magic
tech gf180mcuD
magscale 1 10
timestamp 1757859342
<< nwell >>
rect 6878 4466 7074 4984
rect 8323 4983 8917 4984
rect 9497 4983 9930 4984
rect 8323 4959 9930 4983
rect 8271 4839 9930 4959
rect 8323 4718 9930 4839
rect 8364 4566 8445 4718
rect 8364 4495 8519 4566
rect 8364 4467 8445 4495
rect 8368 4466 8445 4467
rect 8805 4353 9930 4718
rect 8413 4223 9930 4353
rect 9497 4221 9930 4223
rect 9750 4220 9930 4221
rect 6880 2597 7058 3613
rect 8885 3607 9074 3796
rect 9429 3607 9611 3789
rect 7576 3150 7711 3170
rect 7576 3146 7712 3150
rect 7134 3078 8282 3146
rect 8361 3125 9613 3607
rect 8361 3108 9614 3125
rect 7576 3071 7712 3078
rect 8500 2890 9614 3108
rect 8829 2889 9614 2890
rect 9433 2885 9614 2889
rect 24 2470 6860 2532
rect 6878 1232 7061 1741
rect 7438 1232 8182 1248
rect 6878 1168 8182 1232
rect 6878 704 7061 1168
rect 7438 700 8182 1168
<< pwell >>
rect 7667 4081 7847 4096
rect 7135 4017 8281 4081
rect 7667 4002 7847 4017
rect 8172 2345 8853 2400
rect 8172 1936 9491 2345
rect 8172 1743 9489 1936
rect 8748 1639 9489 1743
rect 8488 1352 9490 1639
rect 8487 1348 9718 1352
rect 8486 913 9718 1348
rect 8487 693 9718 913
<< psubdiff >>
rect 7667 4002 7847 4096
rect 8654 2220 9342 2246
rect 8654 2124 8744 2220
rect 9289 2124 9342 2220
rect 8654 2094 9342 2124
rect 8496 818 9649 854
rect 8496 752 8617 818
rect 9514 752 9649 818
rect 8496 733 9649 752
<< nsubdiff >>
rect 8502 4925 8725 4942
rect 8502 4872 8526 4925
rect 8701 4872 8725 4925
rect 8502 4854 8725 4872
rect 9349 4917 9562 4930
rect 9349 4867 9369 4917
rect 9537 4867 9562 4917
rect 9349 4852 9562 4867
rect 9770 4795 9850 4850
rect 9770 4429 9790 4795
rect 9836 4429 9850 4795
rect 9770 4360 9850 4429
rect 7576 3150 7711 3170
rect 8738 3163 9254 3191
rect 7576 3071 7712 3150
rect 8738 3065 8812 3163
rect 9213 3065 9254 3163
rect 8738 3046 9254 3065
rect 24 2470 6860 2532
rect 7948 1182 8099 1250
rect 7948 768 7976 1182
rect 8060 768 8099 1182
rect 7948 724 8099 768
<< psubdiffcont >>
rect 8744 2124 9289 2220
rect 8617 752 9514 818
<< nsubdiffcont >>
rect 8526 4872 8701 4925
rect 9369 4867 9537 4917
rect 9790 4429 9836 4795
rect 8812 3065 9213 3163
rect 7976 768 8060 1182
<< polysilicon >>
rect 2290 2750 2360 4750
rect 4530 2750 4600 4750
rect 9186 4628 9322 4709
rect 2290 250 2360 2250
rect 4520 250 4590 2250
rect 7660 1062 7790 1143
<< metal1 >>
rect 8889 4960 9591 4961
rect 8889 4959 10095 4960
rect 6845 4838 7155 4959
rect 8271 4925 10095 4959
rect 8271 4872 8526 4925
rect 8701 4917 10095 4925
rect 8701 4872 9369 4917
rect 8271 4867 9369 4872
rect 9537 4867 10095 4917
rect 8271 4839 10095 4867
rect 8420 4566 8469 4839
rect 8420 4565 8519 4566
rect 8138 4524 8201 4541
rect 7208 4500 7302 4524
rect 7208 4407 7226 4500
rect 7287 4407 7302 4500
rect 8189 4455 8201 4524
rect 8420 4495 8541 4565
rect 8138 4430 8201 4455
rect 7208 4384 7302 4407
rect 8709 4402 8828 4567
rect 9082 4565 9133 4839
rect 9770 4795 9851 4839
rect 9186 4693 9322 4709
rect 9186 4641 9220 4693
rect 9302 4641 9322 4693
rect 9186 4628 9322 4641
rect 9082 4564 9174 4565
rect 9081 4530 9174 4564
rect 9081 4518 9173 4530
rect 8975 4463 9082 4470
rect 8975 4411 8992 4463
rect 9044 4411 9082 4463
rect 8975 4403 9082 4411
rect 9350 4401 9468 4566
rect 9603 4488 9685 4507
rect 9603 4416 9619 4488
rect 9674 4416 9685 4488
rect 9603 4401 9685 4416
rect 9770 4429 9790 4795
rect 9836 4429 9851 4795
rect 9770 4360 9851 4429
rect 8982 4329 9502 4337
rect 8982 4275 9592 4329
rect 8982 4268 9502 4275
rect 8960 4258 9502 4268
rect 7667 4081 7847 4096
rect 8223 4081 9991 4120
rect 7135 4017 9991 4081
rect 7667 4002 7847 4017
rect 8223 3941 9991 4017
rect 9227 3940 9991 3941
rect 7215 3672 7269 3692
rect 7215 3572 7238 3672
rect 8577 3653 8638 3668
rect 8577 3583 8584 3653
rect 8636 3583 8638 3653
rect 9106 3667 9181 3681
rect 9106 3600 9116 3667
rect 9174 3600 9181 3667
rect 7215 3552 7269 3572
rect 8577 3569 8638 3583
rect 8762 3569 8821 3596
rect 9106 3582 9181 3600
rect 8753 3561 8821 3569
rect 9294 3579 9379 3598
rect 8752 3560 8828 3561
rect 8752 3506 8762 3560
rect 8816 3506 8828 3560
rect 8752 3498 8828 3506
rect 9294 3511 9314 3579
rect 9368 3511 9379 3579
rect 9294 3498 9379 3511
rect 8755 3422 9220 3432
rect 8755 3365 9196 3422
rect 8755 3363 9220 3365
rect 8737 3353 9220 3363
rect 6846 3155 7146 3241
rect 6827 3146 7147 3155
rect 7576 3150 7711 3170
rect 8189 3163 9350 3244
rect 7576 3146 7712 3150
rect 8189 3146 8812 3163
rect 6827 3078 8812 3146
rect 6827 2968 7147 3078
rect 7576 3071 7712 3078
rect 8189 3065 8812 3078
rect 9213 3065 9350 3163
rect 8189 2969 9350 3065
rect 8182 2968 9350 2969
rect 6941 2912 7012 2913
rect 6939 2910 7074 2912
rect 6939 2895 7146 2910
rect 6939 2818 7090 2895
rect 7144 2818 7146 2895
rect 6939 2801 7146 2818
rect 37 2456 6847 2542
rect 6941 1774 7012 2801
rect 7195 2638 7318 2664
rect 7195 2552 7222 2638
rect 7295 2552 7318 2638
rect 7195 2530 7318 2552
rect 8174 2617 8275 2637
rect 8174 2538 8193 2617
rect 8268 2538 8275 2617
rect 8174 2523 8275 2538
rect 9871 2305 9991 3940
rect 9466 2303 9991 2305
rect 8414 2226 9991 2303
rect 8095 2220 9991 2226
rect 8095 2124 8744 2220
rect 9289 2124 9991 2220
rect 8095 2033 9991 2124
rect 8521 2032 9472 2033
rect 7231 1788 7331 1812
rect 7231 1774 7254 1788
rect 6941 1697 7254 1774
rect 7231 1689 7254 1697
rect 7313 1689 7331 1788
rect 8513 1782 8583 1794
rect 8513 1713 8524 1782
rect 8576 1713 8583 1782
rect 8696 1777 8780 1796
rect 8696 1724 8714 1777
rect 8766 1724 8780 1777
rect 8696 1715 8780 1724
rect 9100 1791 9171 1806
rect 9100 1733 9112 1791
rect 9164 1733 9171 1791
rect 9100 1727 9171 1733
rect 9283 1795 9362 1809
rect 9283 1735 9297 1795
rect 9350 1735 9362 1795
rect 9100 1718 9126 1727
rect 9283 1723 9362 1735
rect 8513 1699 8583 1713
rect 7231 1670 7331 1689
rect 9322 1685 9362 1723
rect 9322 1631 9490 1685
rect 7951 1517 8639 1583
rect 8678 1513 9231 1584
rect 9437 1499 9490 1631
rect 9437 1442 9715 1499
rect 6846 1249 7159 1371
rect 8590 1323 9560 1341
rect 7081 1000 7127 1249
rect 7081 936 7181 1000
rect 7554 999 7601 1285
rect 8590 1282 8609 1323
rect 8663 1282 9560 1323
rect 8663 1280 9484 1282
rect 7948 1182 8099 1250
rect 7660 1130 7790 1143
rect 7660 1077 7684 1130
rect 7779 1077 7790 1130
rect 7660 1062 7790 1077
rect 7328 951 7411 968
rect 7328 880 7344 951
rect 7396 880 7411 951
rect 7554 929 7638 999
rect 7798 946 7884 964
rect 7328 859 7411 880
rect 7798 878 7811 946
rect 7869 878 7884 946
rect 7798 866 7884 878
rect 7948 768 7976 1182
rect 8060 768 8099 1182
rect 8501 1143 8558 1167
rect 8501 1087 8517 1143
rect 8501 1072 8558 1087
rect 8711 1048 8839 1212
rect 9024 1050 9123 1215
rect 9657 1214 9714 1442
rect 9609 1213 9714 1214
rect 9315 1050 9421 1213
rect 9567 1156 9714 1213
rect 9032 1049 9096 1050
rect 9040 854 9096 1049
rect 9871 854 9991 2033
rect 7948 724 8099 768
rect 8496 818 9991 854
rect 8496 752 8617 818
rect 9514 752 9991 818
rect 8496 734 9991 752
rect 8496 733 9649 734
<< via1 >>
rect 8565 4646 8662 4698
rect 7226 4407 7287 4500
rect 7467 4414 7531 4466
rect 7943 4431 8027 4483
rect 8136 4455 8189 4524
rect 9220 4641 9302 4693
rect 8992 4411 9044 4463
rect 9619 4416 9674 4488
rect 8877 4269 8971 4324
rect 7392 3750 7449 3842
rect 7238 3572 7301 3672
rect 7948 3602 8032 3656
rect 8584 3583 8636 3653
rect 9116 3600 9174 3667
rect 8762 3506 8816 3560
rect 9314 3511 9368 3579
rect 8092 3315 8152 3389
rect 8652 3362 8735 3420
rect 9196 3365 9278 3422
rect 2269 2999 2387 3115
rect 4491 2987 4622 3114
rect 7090 2818 7144 2895
rect 2259 1933 2397 2028
rect 4494 1937 4632 2032
rect 7222 2552 7295 2638
rect 8193 2538 8268 2617
rect 7254 1689 7313 1788
rect 8524 1713 8576 1782
rect 8714 1724 8766 1777
rect 9112 1733 9164 1791
rect 9297 1735 9350 1795
rect 7211 1076 7302 1132
rect 8609 1271 8663 1323
rect 7684 1077 7779 1130
rect 7344 880 7396 951
rect 7811 878 7869 946
rect 8517 1087 8570 1143
rect 8896 944 8964 996
rect 9183 948 9250 1000
<< metal2 >>
rect 6941 4496 7010 5370
rect 7455 5267 7549 5371
rect 7208 4500 7302 4524
rect 7208 4496 7226 4500
rect 6941 4407 7226 4496
rect 7287 4407 7302 4500
rect 6941 4397 7302 4407
rect 7455 4466 7550 5267
rect 7455 4414 7467 4466
rect 7531 4414 7550 4466
rect 7455 4402 7550 4414
rect 7455 4401 7545 4402
rect 6941 3655 7010 4397
rect 7208 4384 7302 4397
rect 7626 4250 7701 5370
rect 7947 4751 8680 4755
rect 7943 4729 8680 4751
rect 7943 4698 8566 4729
rect 7943 4668 8565 4698
rect 7943 4494 8028 4668
rect 8544 4646 8565 4668
rect 8671 4648 8680 4729
rect 8792 4710 8869 4720
rect 8662 4646 8680 4648
rect 8544 4629 8680 4646
rect 8791 4709 9212 4710
rect 8791 4703 9322 4709
rect 8791 4637 9197 4703
rect 9314 4637 9322 4703
rect 8791 4629 9322 4637
rect 8116 4524 8200 4541
rect 7928 4483 8040 4494
rect 7928 4431 7943 4483
rect 8027 4431 8040 4483
rect 7928 4415 8040 4431
rect 8116 4455 8136 4524
rect 8189 4518 8200 4524
rect 8792 4518 8869 4629
rect 9186 4628 9322 4629
rect 8189 4455 8869 4518
rect 9603 4488 9685 4507
rect 8116 4444 8869 4455
rect 8116 4430 8200 4444
rect 8792 4443 8869 4444
rect 8975 4463 9136 4470
rect 8975 4411 8992 4463
rect 9044 4411 9136 4463
rect 9603 4425 9619 4488
rect 8975 4403 9136 4411
rect 7935 4339 8022 4345
rect 8855 4339 8984 4341
rect 7935 4324 8984 4339
rect 7935 4269 8877 4324
rect 8971 4269 8984 4324
rect 7935 4260 8984 4269
rect 7382 4179 7721 4250
rect 7383 3854 7454 4179
rect 7383 3842 7456 3854
rect 7383 3750 7392 3842
rect 7449 3750 7456 3842
rect 7383 3736 7456 3750
rect 7215 3672 7319 3691
rect 7215 3655 7238 3672
rect 6941 3572 7238 3655
rect 7301 3572 7319 3672
rect 7935 3665 8022 4260
rect 8855 4259 8984 4260
rect 8660 4200 8850 4201
rect 9056 4200 9136 4403
rect 9602 4416 9619 4425
rect 9674 4416 9685 4488
rect 9602 4401 9685 4416
rect 8577 4120 9136 4200
rect 9200 4340 9280 4341
rect 9602 4340 9680 4401
rect 9200 4260 9680 4340
rect 9200 4127 9280 4260
rect 9602 4259 9680 4260
rect 7929 3656 8041 3665
rect 8578 3661 8643 4120
rect 7929 3602 7948 3656
rect 8032 3602 8041 3656
rect 7929 3584 8041 3602
rect 8576 3653 8643 3661
rect 6941 3556 7319 3572
rect 8576 3583 8584 3653
rect 8636 3583 8643 3653
rect 8576 3570 8643 3583
rect 8753 3562 8820 3649
rect 8753 3561 8884 3562
rect 2244 3138 2411 3141
rect 4786 3138 6269 3141
rect 2217 3115 6269 3138
rect 2217 2999 2269 3115
rect 2387 3114 6269 3115
rect 2387 2999 4491 3114
rect 2217 2987 4491 2999
rect 4622 3106 6269 3114
rect 4622 2987 6084 3106
rect 6241 2987 6269 3106
rect 2217 2971 6269 2987
rect 2217 2969 4849 2971
rect 6941 2616 7010 3556
rect 7215 3552 7319 3556
rect 8752 3560 8884 3561
rect 8752 3506 8762 3560
rect 8816 3506 8884 3560
rect 8752 3498 8884 3506
rect 8633 3427 8766 3435
rect 8567 3420 8766 3427
rect 7223 3393 7307 3395
rect 8088 3393 8191 3404
rect 7223 3390 8191 3393
rect 7223 3389 8099 3390
rect 7223 3315 8092 3389
rect 7223 3314 8099 3315
rect 8177 3314 8191 3390
rect 7223 3311 8191 3314
rect 7223 3262 7307 3311
rect 8088 3297 8191 3311
rect 8567 3362 8652 3420
rect 8735 3362 8766 3420
rect 8567 3351 8766 3362
rect 8828 3407 8884 3498
rect 8948 3462 9009 4120
rect 9199 3952 9281 4127
rect 9199 3945 9596 3952
rect 9105 3862 9596 3945
rect 9105 3667 9180 3862
rect 9265 3860 9596 3862
rect 9105 3600 9116 3667
rect 9174 3600 9180 3667
rect 9105 3582 9180 3600
rect 9523 3858 9596 3860
rect 9294 3579 9379 3598
rect 9294 3511 9314 3579
rect 9368 3578 9379 3579
rect 9368 3511 9422 3578
rect 9294 3498 9422 3511
rect 8948 3442 9010 3462
rect 7222 2907 7307 3262
rect 7108 2906 7307 2907
rect 7080 2895 7307 2906
rect 7080 2818 7090 2895
rect 7144 2818 7307 2895
rect 7080 2811 7307 2818
rect 7080 2810 7279 2811
rect 7222 2664 7307 2667
rect 7195 2638 7318 2664
rect 7195 2616 7222 2638
rect 6941 2552 7222 2616
rect 7295 2552 7318 2638
rect 6941 2542 7318 2552
rect 6944 2541 7318 2542
rect 7195 2530 7318 2541
rect 8174 2617 8275 2637
rect 8174 2538 8193 2617
rect 8268 2538 8275 2617
rect 8174 2523 8275 2538
rect 8567 2481 8654 3351
rect 8828 3295 8885 3407
rect 8719 3239 8885 3295
rect 8720 3152 8776 3239
rect 8949 3166 9010 3442
rect 9173 3422 9309 3435
rect 9173 3365 9196 3422
rect 9278 3365 9309 3422
rect 9173 3353 9309 3365
rect 9365 3422 9422 3498
rect 9365 3350 9424 3422
rect 9367 3256 9424 3350
rect 8720 3037 8777 3152
rect 8389 2379 8654 2481
rect 8567 2378 8654 2379
rect 8719 2109 8777 3037
rect 8837 3095 9010 3166
rect 9100 3196 9424 3256
rect 9100 3121 9281 3196
rect 9367 3194 9424 3196
rect 8837 2810 8919 3095
rect 8719 2056 8776 2109
rect 5583 2047 5736 2048
rect 2136 2032 5736 2047
rect 2136 2028 4494 2032
rect 2136 1933 2259 2028
rect 2397 1937 4494 2028
rect 4632 2017 5736 2032
rect 4632 1937 5607 2017
rect 2397 1936 5607 1937
rect 5725 1936 5736 2017
rect 2397 1933 5736 1936
rect 2136 1915 5736 1933
rect 5583 1914 5736 1915
rect 8424 2046 8556 2047
rect 8719 2046 8775 2056
rect 8424 2025 8775 2046
rect 8424 1935 8449 2025
rect 8534 1990 8775 2025
rect 8534 1935 8583 1990
rect 8719 1989 8775 1990
rect 8424 1913 8583 1935
rect 8838 1942 8919 2810
rect 9100 2995 9130 3121
rect 9265 2995 9281 3121
rect 9100 2971 9281 2995
rect 8838 1933 8920 1942
rect 7231 1788 7331 1812
rect 8513 1807 8583 1913
rect 7231 1787 7254 1788
rect 7228 1689 7254 1787
rect 7313 1689 7331 1788
rect 7228 1679 7331 1689
rect 7231 1670 7331 1679
rect 8143 1782 8583 1807
rect 8714 1867 8920 1933
rect 8714 1796 8812 1867
rect 8143 1713 8524 1782
rect 8576 1713 8583 1782
rect 8696 1777 8812 1796
rect 8696 1724 8714 1777
rect 8766 1724 8812 1777
rect 8696 1715 8812 1724
rect 9100 1805 9171 2971
rect 9523 2907 9597 3858
rect 9741 3127 9824 3140
rect 9741 2989 9761 3127
rect 9817 2989 9824 3127
rect 9741 2970 9824 2989
rect 9282 2833 9597 2907
rect 9100 1791 9176 1805
rect 9100 1733 9112 1791
rect 9164 1733 9176 1791
rect 9100 1718 9176 1733
rect 9283 1795 9364 2833
rect 9283 1735 9297 1795
rect 9350 1767 9364 1795
rect 9350 1735 9362 1767
rect 9283 1723 9362 1735
rect 8143 1699 8583 1713
rect 8143 1698 8547 1699
rect 6919 1144 7245 1145
rect 7312 1144 7683 1145
rect 6919 1143 7683 1144
rect 6919 1134 7790 1143
rect 6919 1075 6932 1134
rect 6993 1132 7790 1134
rect 6993 1076 7211 1132
rect 7302 1130 7790 1132
rect 7302 1077 7684 1130
rect 7779 1077 7790 1130
rect 7302 1076 7790 1077
rect 6993 1075 7790 1076
rect 6919 1066 7790 1075
rect 7183 1065 7790 1066
rect 7183 1062 7315 1065
rect 7660 1062 7790 1065
rect 7328 951 7411 968
rect 7328 880 7344 951
rect 7396 880 7411 951
rect 7328 859 7411 880
rect 7798 946 7884 964
rect 7798 878 7811 946
rect 7869 942 7884 946
rect 7869 941 8022 942
rect 8143 941 8208 1698
rect 8739 1465 8812 1715
rect 8351 1385 8812 1465
rect 8351 1166 8430 1385
rect 8587 1323 8686 1327
rect 8587 1321 8609 1323
rect 8663 1321 8686 1323
rect 8587 1265 8606 1321
rect 8671 1265 8686 1321
rect 8587 1249 8686 1265
rect 8501 1166 8575 1167
rect 8351 1143 8575 1166
rect 8351 1087 8517 1143
rect 8570 1087 8575 1143
rect 8501 1072 8575 1087
rect 7869 878 8208 941
rect 8878 996 8999 1003
rect 8878 944 8896 996
rect 8964 987 8999 996
rect 8878 929 8901 944
rect 8968 929 8999 987
rect 8878 918 8999 929
rect 9166 1000 9270 1008
rect 9166 990 9183 1000
rect 9250 990 9270 1000
rect 9166 932 9182 990
rect 9251 932 9270 990
rect 9166 914 9270 932
rect 7798 866 7884 878
rect 7339 687 7401 859
rect 7339 685 8444 687
rect 9765 685 9824 2970
rect 7339 626 9825 685
rect 7340 625 9825 626
rect 9765 623 9824 625
<< via2 >>
rect 8566 4698 8671 4729
rect 8566 4648 8662 4698
rect 8662 4648 8671 4698
rect 9197 4693 9314 4703
rect 9197 4641 9220 4693
rect 9220 4641 9302 4693
rect 9302 4641 9314 4693
rect 9197 4637 9314 4641
rect 6084 2987 6241 3106
rect 8099 3389 8177 3390
rect 8099 3315 8152 3389
rect 8152 3315 8177 3389
rect 8099 3314 8177 3315
rect 8193 2538 8268 2617
rect 5607 1936 5725 2017
rect 8449 1935 8534 2025
rect 9130 2995 9265 3121
rect 9761 2989 9817 3127
rect 6932 1075 6993 1134
rect 8606 1271 8609 1321
rect 8609 1271 8663 1321
rect 8663 1271 8671 1321
rect 8606 1265 8671 1271
rect 8901 944 8964 987
rect 8964 944 8968 987
rect 8901 929 8968 944
rect 9182 948 9183 990
rect 9183 948 9250 990
rect 9250 948 9251 990
rect 9182 932 9251 948
<< metal3 >>
rect 8546 4729 8680 4741
rect 8546 4648 8566 4729
rect 8671 4648 8680 4729
rect 8546 4631 8680 4648
rect 9185 4703 9323 4739
rect 9185 4637 9197 4703
rect 9314 4637 9323 4703
rect 9185 4629 9323 4637
rect 8088 3390 8191 3404
rect 8088 3314 8099 3390
rect 8177 3314 8191 3390
rect 8088 3297 8191 3314
rect 6063 3139 9067 3141
rect 9198 3139 10208 3140
rect 6063 3127 10208 3139
rect 6063 3121 9761 3127
rect 6063 3106 9130 3121
rect 6063 2987 6084 3106
rect 6241 2995 9130 3106
rect 9265 2995 9761 3121
rect 6241 2989 9761 2995
rect 9817 2989 10208 3127
rect 6241 2987 10208 2989
rect 6063 2969 10208 2987
rect 9058 2968 9280 2969
rect 7507 2683 7672 2684
rect 7507 2681 8282 2683
rect 7507 2677 8283 2681
rect 7507 2609 7522 2677
rect 7613 2617 8283 2677
rect 7613 2609 8193 2617
rect 7507 2593 8193 2609
rect 7627 2592 8193 2593
rect 8174 2538 8193 2592
rect 8268 2538 8283 2617
rect 8174 2523 8283 2538
rect 5583 2046 8556 2047
rect 5583 2025 10164 2046
rect 5583 2017 8449 2025
rect 5583 1936 5607 2017
rect 5725 1936 8449 2017
rect 5583 1935 8449 1936
rect 8534 1935 10164 2025
rect 5583 1914 10164 1935
rect 8424 1913 10164 1914
rect 8587 1321 8686 1340
rect 8587 1265 8606 1321
rect 8671 1265 8686 1321
rect 8587 1249 8686 1265
rect 6920 1134 7001 1145
rect 6920 1075 6932 1134
rect 6993 1075 7001 1134
rect 6920 1065 7001 1075
rect 8878 987 8999 1003
rect 8878 929 8901 987
rect 8968 929 8999 987
rect 8878 918 8999 929
rect 9166 990 9270 1008
rect 9166 932 9182 990
rect 9251 932 9270 990
rect 9166 914 9270 932
<< via3 >>
rect 8566 4648 8671 4729
rect 9197 4637 9314 4703
rect 8099 3314 8177 3390
rect 7522 2609 7613 2677
rect 8606 1265 8671 1321
rect 6932 1075 6993 1134
rect 8901 929 8968 987
rect 9182 932 9251 990
<< metal4 >>
rect 8545 4729 8681 4751
rect 8545 4648 8566 4729
rect 8671 4648 8681 4729
rect 8545 4629 8681 4648
rect 9166 4737 9263 4739
rect 9166 4703 9324 4737
rect 9166 4637 9197 4703
rect 9314 4637 9324 4703
rect 8547 3869 8680 4629
rect 9166 4628 9324 4637
rect 8088 3390 8191 3404
rect 8088 3314 8099 3390
rect 8177 3314 8191 3390
rect 8088 3297 8191 3314
rect 7009 2677 7627 2682
rect 7009 2676 7522 2677
rect 6920 2609 7522 2676
rect 7613 2676 7627 2677
rect 7613 2609 7750 2676
rect 6920 2598 7750 2609
rect 6920 2595 7627 2598
rect 6920 1134 7002 2595
rect 8089 1341 8176 3297
rect 8548 1933 8679 3869
rect 8548 1813 9000 1933
rect 8089 1321 8687 1341
rect 8089 1265 8606 1321
rect 8671 1265 8687 1321
rect 8089 1251 8687 1265
rect 6920 1075 6932 1134
rect 6993 1075 7002 1134
rect 6920 -144 7002 1075
rect 8878 987 8999 1813
rect 8878 929 8901 987
rect 8968 929 8999 987
rect 8878 918 8999 929
rect 9166 1008 9263 4628
rect 9166 990 9270 1008
rect 9166 932 9182 990
rect 9251 932 9270 990
rect 9166 914 9270 932
use inv_nand3_1  inv_nand3_1_0
timestamp 1757859342
transform 1 0 7134 0 1 2245
box -86 -1022 1377 870
use nand_inv  nand_inv_0
timestamp 1757859342
transform 1 0 7138 0 1 4118
box -90 -90 1230 866
use nand_inv  nand_inv_1
timestamp 1757859342
transform 1 0 7139 0 -1 3961
box -90 -90 1230 866
use nfet_03v3_084  nfet_03v3_084_0
timestamp 1757514670
transform -1 0 8780 0 -1 1865
box 0 0 280 370
use nfet_03v3_084  nfet_03v3_084_1
timestamp 1757514670
transform -1 0 9367 0 -1 1866
box 0 0 280 370
use nfet_03v3_084  nfet_03v3_084_2
timestamp 1757514670
transform 1 0 8492 0 1 978
box 0 0 280 370
use nfet_03v3_084  nfet_03v3_084_3
timestamp 1757514670
transform -1 0 9071 0 -1 1283
box 0 0 280 370
use nfet_03v3_084  nfet_03v3_084_4
timestamp 1757514670
transform -1 0 9360 0 -1 1285
box 0 0 280 370
use nfet_03v3_084  nfet_03v3_084_5
timestamp 1757514670
transform 1 0 9370 0 1 980
box 0 0 280 370
use pfet_03v3_10  pfet_03v3_10_0
timestamp 1757514455
transform 0 -1 6764 1 0 120
box -120 -120 2380 6764
use pfet_03v3_10  pfet_03v3_10_1
timestamp 1757514455
transform 0 -1 6764 1 0 2620
box -120 -120 2380 6764
use pfet_03v3_084  pfet_03v3_084_0
timestamp 1757513722
transform 1 0 8492 0 1 4342
box -79 -72 325 403
use pfet_03v3_084  pfet_03v3_084_1
timestamp 1757513722
transform -1 0 9040 0 -1 4627
box -79 -72 325 403
use pfet_03v3_084  pfet_03v3_084_2
timestamp 1757513722
transform 1 0 9133 0 1 4341
box -79 -72 325 403
use pfet_03v3_084  pfet_03v3_084_3
timestamp 1757513722
transform -1 0 9668 0 -1 4626
box -79 -72 325 403
use pfet_03v3_084  pfet_03v3_084_4
timestamp 1757513722
transform -1 0 8818 0 -1 3722
box -79 -72 325 403
use pfet_03v3_084  pfet_03v3_084_5
timestamp 1757513722
transform -1 0 9360 0 -1 3721
box -79 -72 325 403
use pfet_03v3_084  pfet_03v3_084_6
timestamp 1757513722
transform 1 0 7130 0 1 776
box -79 -72 325 403
use pfet_03v3_084  pfet_03v3_084_7
timestamp 1757513722
transform 1 0 7606 0 1 775
box -79 -72 325 403
<< labels >>
flabel metal2 7455 5231 7548 5371 0 FreeSans 160 0 0 0 CAL_RESULT
port 7 nsew
flabel metal2 6941 5276 7010 5370 0 FreeSans 160 0 0 0 CAL_CYCLE
port 8 nsew
flabel metal2 7628 5237 7700 5368 0 FreeSans 160 0 0 0 EN_COMP
port 1 nsew
flabel metal3 10010 2980 10201 3130 0 FreeSans 320 0 0 0 CAL_P
port 3 nsew
flabel metal3 9968 1922 10148 2030 0 FreeSans 320 0 0 0 CAL_N
port 2 nsew
flabel metal2 8200 4676 8370 4747 0 FreeSans 160 0 0 0 CAL_RESULT_Z
flabel metal2 7941 3673 8015 3820 0 FreeSans 160 0 0 0 EN_COMP_Z
flabel metal1 8209 1521 8471 1579 0 FreeSans 160 0 0 0 LOAD_CALi
flabel metal2 7858 3313 8064 3388 0 FreeSans 160 0 0 0 EN_COMPi
flabel metal2 8204 4445 8387 4517 0 FreeSans 160 0 0 0 CAL_RESULTi
flabel metal1 9826 4839 10095 4960 0 FreeSans 320 0 0 0 VDD
port 4 nsew
flabel metal1 9492 2085 9736 2261 0 FreeSans 320 0 0 0 VSS
port 5 nsew
flabel metal4 6920 -144 7001 -60 0 FreeSans 320 0 0 0 EN
port 6 nsew
flabel metal2 7953 2213 8379 2274 0 FreeSans 160 0 0 0 LOAD_CAL_Z
<< end >>
