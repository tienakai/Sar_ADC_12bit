magic
tech gf180mcuD
magscale 1 10
timestamp 1757750971
<< error_p >>
rect -2100 833 -2089 879
rect -1758 833 -1747 879
rect -1416 833 -1405 879
rect -1074 833 -1063 879
rect -732 833 -721 879
rect -390 833 -379 879
rect -48 833 -37 879
rect 294 833 305 879
rect 636 833 647 879
rect 978 833 989 879
rect 1320 833 1331 879
rect 1662 833 1673 879
rect 2004 833 2015 879
rect -2100 -879 -2089 -833
rect -1758 -879 -1747 -833
rect -1416 -879 -1405 -833
rect -1074 -879 -1063 -833
rect -732 -879 -721 -833
rect -390 -879 -379 -833
rect -48 -879 -37 -833
rect 294 -879 305 -833
rect 636 -879 647 -833
rect 978 -879 989 -833
rect 1320 -879 1331 -833
rect 1662 -879 1673 -833
rect 2004 -879 2015 -833
<< nwell >>
rect -2276 -978 2276 978
<< pmos >>
rect -2102 -800 -2002 800
rect -1760 -800 -1660 800
rect -1418 -800 -1318 800
rect -1076 -800 -976 800
rect -734 -800 -634 800
rect -392 -800 -292 800
rect -50 -800 50 800
rect 292 -800 392 800
rect 634 -800 734 800
rect 976 -800 1076 800
rect 1318 -800 1418 800
rect 1660 -800 1760 800
rect 2002 -800 2102 800
<< pdiff >>
rect -2190 787 -2102 800
rect -2190 -787 -2177 787
rect -2131 -787 -2102 787
rect -2190 -800 -2102 -787
rect -2002 787 -1914 800
rect -2002 -787 -1973 787
rect -1927 -787 -1914 787
rect -2002 -800 -1914 -787
rect -1848 787 -1760 800
rect -1848 -787 -1835 787
rect -1789 -787 -1760 787
rect -1848 -800 -1760 -787
rect -1660 787 -1572 800
rect -1660 -787 -1631 787
rect -1585 -787 -1572 787
rect -1660 -800 -1572 -787
rect -1506 787 -1418 800
rect -1506 -787 -1493 787
rect -1447 -787 -1418 787
rect -1506 -800 -1418 -787
rect -1318 787 -1230 800
rect -1318 -787 -1289 787
rect -1243 -787 -1230 787
rect -1318 -800 -1230 -787
rect -1164 787 -1076 800
rect -1164 -787 -1151 787
rect -1105 -787 -1076 787
rect -1164 -800 -1076 -787
rect -976 787 -888 800
rect -976 -787 -947 787
rect -901 -787 -888 787
rect -976 -800 -888 -787
rect -822 787 -734 800
rect -822 -787 -809 787
rect -763 -787 -734 787
rect -822 -800 -734 -787
rect -634 787 -546 800
rect -634 -787 -605 787
rect -559 -787 -546 787
rect -634 -800 -546 -787
rect -480 787 -392 800
rect -480 -787 -467 787
rect -421 -787 -392 787
rect -480 -800 -392 -787
rect -292 787 -204 800
rect -292 -787 -263 787
rect -217 -787 -204 787
rect -292 -800 -204 -787
rect -138 787 -50 800
rect -138 -787 -125 787
rect -79 -787 -50 787
rect -138 -800 -50 -787
rect 50 787 138 800
rect 50 -787 79 787
rect 125 -787 138 787
rect 50 -800 138 -787
rect 204 787 292 800
rect 204 -787 217 787
rect 263 -787 292 787
rect 204 -800 292 -787
rect 392 787 480 800
rect 392 -787 421 787
rect 467 -787 480 787
rect 392 -800 480 -787
rect 546 787 634 800
rect 546 -787 559 787
rect 605 -787 634 787
rect 546 -800 634 -787
rect 734 787 822 800
rect 734 -787 763 787
rect 809 -787 822 787
rect 734 -800 822 -787
rect 888 787 976 800
rect 888 -787 901 787
rect 947 -787 976 787
rect 888 -800 976 -787
rect 1076 787 1164 800
rect 1076 -787 1105 787
rect 1151 -787 1164 787
rect 1076 -800 1164 -787
rect 1230 787 1318 800
rect 1230 -787 1243 787
rect 1289 -787 1318 787
rect 1230 -800 1318 -787
rect 1418 787 1506 800
rect 1418 -787 1447 787
rect 1493 -787 1506 787
rect 1418 -800 1506 -787
rect 1572 787 1660 800
rect 1572 -787 1585 787
rect 1631 -787 1660 787
rect 1572 -800 1660 -787
rect 1760 787 1848 800
rect 1760 -787 1789 787
rect 1835 -787 1848 787
rect 1760 -800 1848 -787
rect 1914 787 2002 800
rect 1914 -787 1927 787
rect 1973 -787 2002 787
rect 1914 -800 2002 -787
rect 2102 787 2190 800
rect 2102 -787 2131 787
rect 2177 -787 2190 787
rect 2102 -800 2190 -787
<< pdiffc >>
rect -2177 -787 -2131 787
rect -1973 -787 -1927 787
rect -1835 -787 -1789 787
rect -1631 -787 -1585 787
rect -1493 -787 -1447 787
rect -1289 -787 -1243 787
rect -1151 -787 -1105 787
rect -947 -787 -901 787
rect -809 -787 -763 787
rect -605 -787 -559 787
rect -467 -787 -421 787
rect -263 -787 -217 787
rect -125 -787 -79 787
rect 79 -787 125 787
rect 217 -787 263 787
rect 421 -787 467 787
rect 559 -787 605 787
rect 763 -787 809 787
rect 901 -787 947 787
rect 1105 -787 1151 787
rect 1243 -787 1289 787
rect 1447 -787 1493 787
rect 1585 -787 1631 787
rect 1789 -787 1835 787
rect 1927 -787 1973 787
rect 2131 -787 2177 787
<< polysilicon >>
rect -2102 879 -2002 892
rect -2102 833 -2089 879
rect -2015 833 -2002 879
rect -2102 800 -2002 833
rect -1760 879 -1660 892
rect -1760 833 -1747 879
rect -1673 833 -1660 879
rect -1760 800 -1660 833
rect -1418 879 -1318 892
rect -1418 833 -1405 879
rect -1331 833 -1318 879
rect -1418 800 -1318 833
rect -1076 879 -976 892
rect -1076 833 -1063 879
rect -989 833 -976 879
rect -1076 800 -976 833
rect -734 879 -634 892
rect -734 833 -721 879
rect -647 833 -634 879
rect -734 800 -634 833
rect -392 879 -292 892
rect -392 833 -379 879
rect -305 833 -292 879
rect -392 800 -292 833
rect -50 879 50 892
rect -50 833 -37 879
rect 37 833 50 879
rect -50 800 50 833
rect 292 879 392 892
rect 292 833 305 879
rect 379 833 392 879
rect 292 800 392 833
rect 634 879 734 892
rect 634 833 647 879
rect 721 833 734 879
rect 634 800 734 833
rect 976 879 1076 892
rect 976 833 989 879
rect 1063 833 1076 879
rect 976 800 1076 833
rect 1318 879 1418 892
rect 1318 833 1331 879
rect 1405 833 1418 879
rect 1318 800 1418 833
rect 1660 879 1760 892
rect 1660 833 1673 879
rect 1747 833 1760 879
rect 1660 800 1760 833
rect 2002 879 2102 892
rect 2002 833 2015 879
rect 2089 833 2102 879
rect 2002 800 2102 833
rect -2102 -833 -2002 -800
rect -2102 -879 -2089 -833
rect -2015 -879 -2002 -833
rect -2102 -892 -2002 -879
rect -1760 -833 -1660 -800
rect -1760 -879 -1747 -833
rect -1673 -879 -1660 -833
rect -1760 -892 -1660 -879
rect -1418 -833 -1318 -800
rect -1418 -879 -1405 -833
rect -1331 -879 -1318 -833
rect -1418 -892 -1318 -879
rect -1076 -833 -976 -800
rect -1076 -879 -1063 -833
rect -989 -879 -976 -833
rect -1076 -892 -976 -879
rect -734 -833 -634 -800
rect -734 -879 -721 -833
rect -647 -879 -634 -833
rect -734 -892 -634 -879
rect -392 -833 -292 -800
rect -392 -879 -379 -833
rect -305 -879 -292 -833
rect -392 -892 -292 -879
rect -50 -833 50 -800
rect -50 -879 -37 -833
rect 37 -879 50 -833
rect -50 -892 50 -879
rect 292 -833 392 -800
rect 292 -879 305 -833
rect 379 -879 392 -833
rect 292 -892 392 -879
rect 634 -833 734 -800
rect 634 -879 647 -833
rect 721 -879 734 -833
rect 634 -892 734 -879
rect 976 -833 1076 -800
rect 976 -879 989 -833
rect 1063 -879 1076 -833
rect 976 -892 1076 -879
rect 1318 -833 1418 -800
rect 1318 -879 1331 -833
rect 1405 -879 1418 -833
rect 1318 -892 1418 -879
rect 1660 -833 1760 -800
rect 1660 -879 1673 -833
rect 1747 -879 1760 -833
rect 1660 -892 1760 -879
rect 2002 -833 2102 -800
rect 2002 -879 2015 -833
rect 2089 -879 2102 -833
rect 2002 -892 2102 -879
<< polycontact >>
rect -2089 833 -2015 879
rect -1747 833 -1673 879
rect -1405 833 -1331 879
rect -1063 833 -989 879
rect -721 833 -647 879
rect -379 833 -305 879
rect -37 833 37 879
rect 305 833 379 879
rect 647 833 721 879
rect 989 833 1063 879
rect 1331 833 1405 879
rect 1673 833 1747 879
rect 2015 833 2089 879
rect -2089 -879 -2015 -833
rect -1747 -879 -1673 -833
rect -1405 -879 -1331 -833
rect -1063 -879 -989 -833
rect -721 -879 -647 -833
rect -379 -879 -305 -833
rect -37 -879 37 -833
rect 305 -879 379 -833
rect 647 -879 721 -833
rect 989 -879 1063 -833
rect 1331 -879 1405 -833
rect 1673 -879 1747 -833
rect 2015 -879 2089 -833
<< metal1 >>
rect -2100 833 -2089 879
rect -2015 833 -2004 879
rect -1758 833 -1747 879
rect -1673 833 -1662 879
rect -1416 833 -1405 879
rect -1331 833 -1320 879
rect -1074 833 -1063 879
rect -989 833 -978 879
rect -732 833 -721 879
rect -647 833 -636 879
rect -390 833 -379 879
rect -305 833 -294 879
rect -48 833 -37 879
rect 37 833 48 879
rect 294 833 305 879
rect 379 833 390 879
rect 636 833 647 879
rect 721 833 732 879
rect 978 833 989 879
rect 1063 833 1074 879
rect 1320 833 1331 879
rect 1405 833 1416 879
rect 1662 833 1673 879
rect 1747 833 1758 879
rect 2004 833 2015 879
rect 2089 833 2100 879
rect -2177 787 -2131 798
rect -2177 -798 -2131 -787
rect -1973 787 -1927 798
rect -1973 -798 -1927 -787
rect -1835 787 -1789 798
rect -1835 -798 -1789 -787
rect -1631 787 -1585 798
rect -1631 -798 -1585 -787
rect -1493 787 -1447 798
rect -1493 -798 -1447 -787
rect -1289 787 -1243 798
rect -1289 -798 -1243 -787
rect -1151 787 -1105 798
rect -1151 -798 -1105 -787
rect -947 787 -901 798
rect -947 -798 -901 -787
rect -809 787 -763 798
rect -809 -798 -763 -787
rect -605 787 -559 798
rect -605 -798 -559 -787
rect -467 787 -421 798
rect -467 -798 -421 -787
rect -263 787 -217 798
rect -263 -798 -217 -787
rect -125 787 -79 798
rect -125 -798 -79 -787
rect 79 787 125 798
rect 79 -798 125 -787
rect 217 787 263 798
rect 217 -798 263 -787
rect 421 787 467 798
rect 421 -798 467 -787
rect 559 787 605 798
rect 559 -798 605 -787
rect 763 787 809 798
rect 763 -798 809 -787
rect 901 787 947 798
rect 901 -798 947 -787
rect 1105 787 1151 798
rect 1105 -798 1151 -787
rect 1243 787 1289 798
rect 1243 -798 1289 -787
rect 1447 787 1493 798
rect 1447 -798 1493 -787
rect 1585 787 1631 798
rect 1585 -798 1631 -787
rect 1789 787 1835 798
rect 1789 -798 1835 -787
rect 1927 787 1973 798
rect 1927 -798 1973 -787
rect 2131 787 2177 798
rect 2131 -798 2177 -787
rect -2100 -879 -2089 -833
rect -2015 -879 -2004 -833
rect -1758 -879 -1747 -833
rect -1673 -879 -1662 -833
rect -1416 -879 -1405 -833
rect -1331 -879 -1320 -833
rect -1074 -879 -1063 -833
rect -989 -879 -978 -833
rect -732 -879 -721 -833
rect -647 -879 -636 -833
rect -390 -879 -379 -833
rect -305 -879 -294 -833
rect -48 -879 -37 -833
rect 37 -879 48 -833
rect 294 -879 305 -833
rect 379 -879 390 -833
rect 636 -879 647 -833
rect 721 -879 732 -833
rect 978 -879 989 -833
rect 1063 -879 1074 -833
rect 1320 -879 1331 -833
rect 1405 -879 1416 -833
rect 1662 -879 1673 -833
rect 1747 -879 1758 -833
rect 2004 -879 2015 -833
rect 2089 -879 2100 -833
<< properties >>
string gencell pfet_03v3
string library gf180mcu
string parameters w 8 l 0.5 m 1 nf 13 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {pfet_03v3 pfet_06v0}
<< end >>
