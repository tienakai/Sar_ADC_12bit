magic
tech gf180mcuD
magscale 1 10
timestamp 1757721953
<< error_p >>
rect -1272 833 -1261 879
rect -1068 833 -1057 879
rect -864 833 -853 879
rect -660 833 -649 879
rect -456 833 -445 879
rect -252 833 -241 879
rect -48 833 -37 879
rect 156 833 167 879
rect 360 833 371 879
rect 564 833 575 879
rect 768 833 779 879
rect 972 833 983 879
rect 1176 833 1187 879
rect -1272 -879 -1261 -833
rect -1068 -879 -1057 -833
rect -864 -879 -853 -833
rect -660 -879 -649 -833
rect -456 -879 -445 -833
rect -252 -879 -241 -833
rect -48 -879 -37 -833
rect 156 -879 167 -833
rect 360 -879 371 -833
rect 564 -879 575 -833
rect 768 -879 779 -833
rect 972 -879 983 -833
rect 1176 -879 1187 -833
<< nwell >>
rect -1448 -978 1448 978
<< pmos >>
rect -1274 -800 -1174 800
rect -1070 -800 -970 800
rect -866 -800 -766 800
rect -662 -800 -562 800
rect -458 -800 -358 800
rect -254 -800 -154 800
rect -50 -800 50 800
rect 154 -800 254 800
rect 358 -800 458 800
rect 562 -800 662 800
rect 766 -800 866 800
rect 970 -800 1070 800
rect 1174 -800 1274 800
<< pdiff >>
rect -1362 787 -1274 800
rect -1362 -787 -1349 787
rect -1303 -787 -1274 787
rect -1362 -800 -1274 -787
rect -1174 787 -1070 800
rect -1174 -787 -1145 787
rect -1099 -787 -1070 787
rect -1174 -800 -1070 -787
rect -970 787 -866 800
rect -970 -787 -941 787
rect -895 -787 -866 787
rect -970 -800 -866 -787
rect -766 787 -662 800
rect -766 -787 -737 787
rect -691 -787 -662 787
rect -766 -800 -662 -787
rect -562 787 -458 800
rect -562 -787 -533 787
rect -487 -787 -458 787
rect -562 -800 -458 -787
rect -358 787 -254 800
rect -358 -787 -329 787
rect -283 -787 -254 787
rect -358 -800 -254 -787
rect -154 787 -50 800
rect -154 -787 -125 787
rect -79 -787 -50 787
rect -154 -800 -50 -787
rect 50 787 154 800
rect 50 -787 79 787
rect 125 -787 154 787
rect 50 -800 154 -787
rect 254 787 358 800
rect 254 -787 283 787
rect 329 -787 358 787
rect 254 -800 358 -787
rect 458 787 562 800
rect 458 -787 487 787
rect 533 -787 562 787
rect 458 -800 562 -787
rect 662 787 766 800
rect 662 -787 691 787
rect 737 -787 766 787
rect 662 -800 766 -787
rect 866 787 970 800
rect 866 -787 895 787
rect 941 -787 970 787
rect 866 -800 970 -787
rect 1070 787 1174 800
rect 1070 -787 1099 787
rect 1145 -787 1174 787
rect 1070 -800 1174 -787
rect 1274 787 1362 800
rect 1274 -787 1303 787
rect 1349 -787 1362 787
rect 1274 -800 1362 -787
<< pdiffc >>
rect -1349 -787 -1303 787
rect -1145 -787 -1099 787
rect -941 -787 -895 787
rect -737 -787 -691 787
rect -533 -787 -487 787
rect -329 -787 -283 787
rect -125 -787 -79 787
rect 79 -787 125 787
rect 283 -787 329 787
rect 487 -787 533 787
rect 691 -787 737 787
rect 895 -787 941 787
rect 1099 -787 1145 787
rect 1303 -787 1349 787
<< polysilicon >>
rect -1274 879 -1174 892
rect -1274 833 -1261 879
rect -1187 833 -1174 879
rect -1274 800 -1174 833
rect -1070 879 -970 892
rect -1070 833 -1057 879
rect -983 833 -970 879
rect -1070 800 -970 833
rect -866 879 -766 892
rect -866 833 -853 879
rect -779 833 -766 879
rect -866 800 -766 833
rect -662 879 -562 892
rect -662 833 -649 879
rect -575 833 -562 879
rect -662 800 -562 833
rect -458 879 -358 892
rect -458 833 -445 879
rect -371 833 -358 879
rect -458 800 -358 833
rect -254 879 -154 892
rect -254 833 -241 879
rect -167 833 -154 879
rect -254 800 -154 833
rect -50 879 50 892
rect -50 833 -37 879
rect 37 833 50 879
rect -50 800 50 833
rect 154 879 254 892
rect 154 833 167 879
rect 241 833 254 879
rect 154 800 254 833
rect 358 879 458 892
rect 358 833 371 879
rect 445 833 458 879
rect 358 800 458 833
rect 562 879 662 892
rect 562 833 575 879
rect 649 833 662 879
rect 562 800 662 833
rect 766 879 866 892
rect 766 833 779 879
rect 853 833 866 879
rect 766 800 866 833
rect 970 879 1070 892
rect 970 833 983 879
rect 1057 833 1070 879
rect 970 800 1070 833
rect 1174 879 1274 892
rect 1174 833 1187 879
rect 1261 833 1274 879
rect 1174 800 1274 833
rect -1274 -833 -1174 -800
rect -1274 -879 -1261 -833
rect -1187 -879 -1174 -833
rect -1274 -892 -1174 -879
rect -1070 -833 -970 -800
rect -1070 -879 -1057 -833
rect -983 -879 -970 -833
rect -1070 -892 -970 -879
rect -866 -833 -766 -800
rect -866 -879 -853 -833
rect -779 -879 -766 -833
rect -866 -892 -766 -879
rect -662 -833 -562 -800
rect -662 -879 -649 -833
rect -575 -879 -562 -833
rect -662 -892 -562 -879
rect -458 -833 -358 -800
rect -458 -879 -445 -833
rect -371 -879 -358 -833
rect -458 -892 -358 -879
rect -254 -833 -154 -800
rect -254 -879 -241 -833
rect -167 -879 -154 -833
rect -254 -892 -154 -879
rect -50 -833 50 -800
rect -50 -879 -37 -833
rect 37 -879 50 -833
rect -50 -892 50 -879
rect 154 -833 254 -800
rect 154 -879 167 -833
rect 241 -879 254 -833
rect 154 -892 254 -879
rect 358 -833 458 -800
rect 358 -879 371 -833
rect 445 -879 458 -833
rect 358 -892 458 -879
rect 562 -833 662 -800
rect 562 -879 575 -833
rect 649 -879 662 -833
rect 562 -892 662 -879
rect 766 -833 866 -800
rect 766 -879 779 -833
rect 853 -879 866 -833
rect 766 -892 866 -879
rect 970 -833 1070 -800
rect 970 -879 983 -833
rect 1057 -879 1070 -833
rect 970 -892 1070 -879
rect 1174 -833 1274 -800
rect 1174 -879 1187 -833
rect 1261 -879 1274 -833
rect 1174 -892 1274 -879
<< polycontact >>
rect -1261 833 -1187 879
rect -1057 833 -983 879
rect -853 833 -779 879
rect -649 833 -575 879
rect -445 833 -371 879
rect -241 833 -167 879
rect -37 833 37 879
rect 167 833 241 879
rect 371 833 445 879
rect 575 833 649 879
rect 779 833 853 879
rect 983 833 1057 879
rect 1187 833 1261 879
rect -1261 -879 -1187 -833
rect -1057 -879 -983 -833
rect -853 -879 -779 -833
rect -649 -879 -575 -833
rect -445 -879 -371 -833
rect -241 -879 -167 -833
rect -37 -879 37 -833
rect 167 -879 241 -833
rect 371 -879 445 -833
rect 575 -879 649 -833
rect 779 -879 853 -833
rect 983 -879 1057 -833
rect 1187 -879 1261 -833
<< metal1 >>
rect -1272 833 -1261 879
rect -1187 833 -1176 879
rect -1068 833 -1057 879
rect -983 833 -972 879
rect -864 833 -853 879
rect -779 833 -768 879
rect -660 833 -649 879
rect -575 833 -564 879
rect -456 833 -445 879
rect -371 833 -360 879
rect -252 833 -241 879
rect -167 833 -156 879
rect -48 833 -37 879
rect 37 833 48 879
rect 156 833 167 879
rect 241 833 252 879
rect 360 833 371 879
rect 445 833 456 879
rect 564 833 575 879
rect 649 833 660 879
rect 768 833 779 879
rect 853 833 864 879
rect 972 833 983 879
rect 1057 833 1068 879
rect 1176 833 1187 879
rect 1261 833 1272 879
rect -1349 787 -1303 798
rect -1349 -798 -1303 -787
rect -1145 787 -1099 798
rect -1145 -798 -1099 -787
rect -941 787 -895 798
rect -941 -798 -895 -787
rect -737 787 -691 798
rect -737 -798 -691 -787
rect -533 787 -487 798
rect -533 -798 -487 -787
rect -329 787 -283 798
rect -329 -798 -283 -787
rect -125 787 -79 798
rect -125 -798 -79 -787
rect 79 787 125 798
rect 79 -798 125 -787
rect 283 787 329 798
rect 283 -798 329 -787
rect 487 787 533 798
rect 487 -798 533 -787
rect 691 787 737 798
rect 691 -798 737 -787
rect 895 787 941 798
rect 895 -798 941 -787
rect 1099 787 1145 798
rect 1099 -798 1145 -787
rect 1303 787 1349 798
rect 1303 -798 1349 -787
rect -1272 -879 -1261 -833
rect -1187 -879 -1176 -833
rect -1068 -879 -1057 -833
rect -983 -879 -972 -833
rect -864 -879 -853 -833
rect -779 -879 -768 -833
rect -660 -879 -649 -833
rect -575 -879 -564 -833
rect -456 -879 -445 -833
rect -371 -879 -360 -833
rect -252 -879 -241 -833
rect -167 -879 -156 -833
rect -48 -879 -37 -833
rect 37 -879 48 -833
rect 156 -879 167 -833
rect 241 -879 252 -833
rect 360 -879 371 -833
rect 445 -879 456 -833
rect 564 -879 575 -833
rect 649 -879 660 -833
rect 768 -879 779 -833
rect 853 -879 864 -833
rect 972 -879 983 -833
rect 1057 -879 1068 -833
rect 1176 -879 1187 -833
rect 1261 -879 1272 -833
<< properties >>
string gencell pfet_03v3
string library gf180mcu
string parameters w 8 l 0.5 m 1 nf 13 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {pfet_03v3 pfet_06v0}
<< end >>
