magic
tech gf180mcuD
magscale 1 10
timestamp 1757721953
<< error_p >>
rect -48 833 -37 879
rect -48 -879 -37 -833
<< nwell >>
rect -300 -1010 300 1010
<< pmos >>
rect -50 -800 50 800
<< pdiff >>
rect -138 787 -50 800
rect -138 -787 -125 787
rect -79 -787 -50 787
rect -138 -800 -50 -787
rect 50 787 138 800
rect 50 -787 79 787
rect 125 -787 138 787
rect 50 -800 138 -787
<< pdiffc >>
rect -125 -787 -79 787
rect 79 -787 125 787
<< nsubdiff >>
rect -276 914 276 986
rect -276 870 -204 914
rect -276 -870 -263 870
rect -217 -870 -204 870
rect 204 870 276 914
rect -276 -914 -204 -870
rect 204 -870 217 870
rect 263 -870 276 870
rect 204 -914 276 -870
rect -276 -986 276 -914
<< nsubdiffcont >>
rect -263 -870 -217 870
rect 217 -870 263 870
<< polysilicon >>
rect -50 879 50 892
rect -50 833 -37 879
rect 37 833 50 879
rect -50 800 50 833
rect -50 -833 50 -800
rect -50 -879 -37 -833
rect 37 -879 50 -833
rect -50 -892 50 -879
<< polycontact >>
rect -37 833 37 879
rect -37 -879 37 -833
<< metal1 >>
rect -263 927 263 973
rect -263 870 -217 927
rect -48 833 -37 879
rect 37 833 48 879
rect 217 870 263 927
rect -125 787 -79 798
rect -125 -798 -79 -787
rect 79 787 125 798
rect 79 -798 125 -787
rect -263 -927 -217 -870
rect -48 -879 -37 -833
rect 37 -879 48 -833
rect 217 -927 263 -870
rect -263 -973 263 -927
<< properties >>
string FIXED_BBOX -240 -950 240 950
string gencell pfet_03v3
string library gf180mcu
string parameters w 8 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {pfet_03v3 pfet_06v0}
<< end >>
