magic
tech gf180mcuD
magscale 1 10
timestamp 1757325932
<< nwell >>
rect 1290 -346 2174 443
<< pwell >>
rect 308 -346 1290 443
<< nmos >>
rect 420 -176 476 224
rect 580 -176 636 224
rect 740 -176 796 224
rect 900 -176 956 224
rect 1060 -176 1116 224
<< pmos >>
rect 1464 -176 1520 224
rect 1624 -176 1680 224
rect 1784 -176 1840 224
rect 1944 -176 2000 224
<< ndiff >>
rect 332 211 420 224
rect 332 -163 345 211
rect 391 -163 420 211
rect 332 -176 420 -163
rect 476 211 580 224
rect 476 -163 505 211
rect 551 -163 580 211
rect 476 -176 580 -163
rect 636 211 740 224
rect 636 -163 665 211
rect 711 -163 740 211
rect 636 -176 740 -163
rect 796 211 900 224
rect 796 -163 825 211
rect 871 -163 900 211
rect 796 -176 900 -163
rect 956 211 1060 224
rect 956 -163 985 211
rect 1031 -163 1060 211
rect 956 -176 1060 -163
rect 1116 211 1204 224
rect 1116 -163 1145 211
rect 1191 -163 1204 211
rect 1116 -176 1204 -163
<< pdiff >>
rect 1376 211 1464 224
rect 1376 -163 1389 211
rect 1435 -163 1464 211
rect 1376 -176 1464 -163
rect 1520 211 1624 224
rect 1520 -163 1549 211
rect 1595 -163 1624 211
rect 1520 -176 1624 -163
rect 1680 211 1784 224
rect 1680 -163 1709 211
rect 1755 -163 1784 211
rect 1680 -176 1784 -163
rect 1840 211 1944 224
rect 1840 -163 1869 211
rect 1915 -163 1944 211
rect 1840 -176 1944 -163
rect 2000 211 2088 224
rect 2000 -163 2029 211
rect 2075 -163 2088 211
rect 2000 -176 2088 -163
<< ndiffc >>
rect 345 -163 391 211
rect 505 -163 551 211
rect 665 -163 711 211
rect 825 -163 871 211
rect 985 -163 1031 211
rect 1145 -163 1191 211
<< pdiffc >>
rect 1389 -163 1435 211
rect 1549 -163 1595 211
rect 1709 -163 1755 211
rect 1869 -163 1915 211
rect 2029 -163 2075 211
<< psubdiff >>
rect 341 -257 540 -242
rect 341 -303 360 -257
rect 519 -303 540 -257
rect 341 -316 540 -303
<< nsubdiff >>
rect 2009 384 2149 398
rect 2009 338 2023 384
rect 2135 338 2149 384
rect 2009 325 2149 338
<< psubdiffcont >>
rect 360 -303 519 -257
<< nsubdiffcont >>
rect 2023 338 2135 384
<< polysilicon >>
rect 420 268 636 304
rect 420 224 476 268
rect 580 224 636 268
rect 740 268 956 304
rect 740 224 796 268
rect 900 224 956 268
rect 1060 224 1116 302
rect 1464 268 2000 304
rect 1464 224 1520 268
rect 1624 224 1680 268
rect 1784 224 1840 268
rect 1944 224 2000 268
rect 420 -220 476 -176
rect 580 -220 636 -176
rect 740 -220 796 -176
rect 900 -220 956 -176
rect 1060 -220 1116 -176
rect 1464 -220 1520 -176
rect 1624 -220 1680 -176
rect 1784 -220 1840 -176
rect 1944 -220 2000 -176
<< metal1 >>
rect 346 384 2172 404
rect 346 338 2023 384
rect 2135 338 2172 384
rect 346 322 2172 338
rect 345 211 391 222
rect 330 -110 345 -106
rect 505 211 551 222
rect 391 -110 406 -106
rect 330 -162 342 -110
rect 394 -162 406 -110
rect 330 -163 345 -162
rect 391 -163 406 -162
rect 330 -174 406 -163
rect 665 211 711 222
rect 505 -174 551 -163
rect 650 -110 665 -106
rect 825 211 871 222
rect 711 -110 726 -106
rect 650 -162 662 -110
rect 714 -162 726 -110
rect 650 -163 665 -162
rect 711 -163 726 -162
rect 650 -174 726 -163
rect 985 211 1031 222
rect 825 -174 871 -163
rect 970 -110 985 -106
rect 1145 211 1191 222
rect 1031 -110 1046 -106
rect 970 -162 982 -110
rect 1034 -162 1046 -110
rect 970 -163 985 -162
rect 1031 -163 1046 -162
rect 970 -174 1046 -163
rect 1374 211 1450 222
rect 1374 210 1389 211
rect 1435 210 1450 211
rect 1374 158 1386 210
rect 1438 158 1450 210
rect 1374 154 1389 158
rect 1145 -174 1191 -163
rect 1435 154 1450 158
rect 1549 211 1595 222
rect 1389 -174 1435 -163
rect 1534 -110 1549 -106
rect 1694 211 1770 222
rect 1694 210 1709 211
rect 1755 210 1770 211
rect 1694 158 1706 210
rect 1758 158 1770 210
rect 1694 154 1709 158
rect 1595 -110 1610 -106
rect 1534 -162 1546 -110
rect 1598 -162 1610 -110
rect 1534 -163 1549 -162
rect 1595 -163 1610 -162
rect 1534 -174 1610 -163
rect 1755 154 1770 158
rect 1869 211 1915 222
rect 1709 -174 1755 -163
rect 1854 -110 1869 -106
rect 2014 211 2090 222
rect 2014 210 2029 211
rect 2075 210 2090 211
rect 2014 158 2026 210
rect 2078 158 2090 210
rect 2014 154 2029 158
rect 1915 -110 1930 -106
rect 1854 -162 1866 -110
rect 1918 -162 1930 -110
rect 1854 -163 1869 -162
rect 1915 -163 1930 -162
rect 1854 -174 1930 -163
rect 2075 154 2090 158
rect 2029 -174 2075 -163
rect 332 -257 2091 -234
rect 332 -303 360 -257
rect 519 -303 2091 -257
rect 332 -316 2091 -303
<< via1 >>
rect 342 -162 345 -110
rect 345 -162 391 -110
rect 391 -162 394 -110
rect 662 -162 665 -110
rect 665 -162 711 -110
rect 711 -162 714 -110
rect 982 -162 985 -110
rect 985 -162 1031 -110
rect 1031 -162 1034 -110
rect 1386 158 1389 210
rect 1389 158 1435 210
rect 1435 158 1438 210
rect 1706 158 1709 210
rect 1709 158 1755 210
rect 1755 158 1758 210
rect 1546 -162 1549 -110
rect 1549 -162 1595 -110
rect 1595 -162 1598 -110
rect 2026 158 2029 210
rect 2029 158 2075 210
rect 2075 158 2078 210
rect 1866 -162 1869 -110
rect 1869 -162 1915 -110
rect 1915 -162 1918 -110
<< metal2 >>
rect 1374 210 2090 222
rect 1374 158 1386 210
rect 1438 158 1706 210
rect 1758 158 2026 210
rect 2078 158 2090 210
rect 1374 154 2090 158
rect 330 -110 1930 -106
rect 330 -162 342 -110
rect 394 -162 662 -110
rect 714 -162 982 -110
rect 1034 -162 1546 -110
rect 1598 -162 1866 -110
rect 1918 -162 1930 -110
rect 330 -174 1930 -162
<< labels >>
flabel polysilicon 1060 242 1116 302 1 FreeSans 320 0 0 0 EN_VIN
port 10 n
flabel polysilicon 1464 268 2000 304 1 FreeSans 320 0 0 0 EN_VREF_Z
port 6 n
flabel metal2 1034 -174 1546 -106 1 FreeSans 400 0 0 0 Cbtm
port 7 n
flabel metal2 1374 154 2090 222 1 FreeSans 400 0 0 0 VREF
port 4 n
flabel polysilicon 740 268 956 304 1 FreeSans 320 0 0 0 EN_VSS
port 9 n
flabel polysilicon 420 268 636 304 1 FreeSans 320 0 0 0 EN_VCM
port 5 n
flabel metal1 505 -174 551 222 1 FreeSans 320 0 0 0 VCM
port 1 n
flabel metal1 825 -174 871 222 1 FreeSans 320 0 0 0 VREF_GND
port 2 n
flabel metal1 1145 -174 1191 222 1 FreeSans 320 0 0 0 VIN
port 3 n
flabel metal1 1376 322 2088 404 1 FreeSans 400 0 0 0 VDD
port 8 n
flabel metal1 332 -316 1204 -234 1 FreeSans 400 0 0 0 VSS
port 11 n
<< end >>
