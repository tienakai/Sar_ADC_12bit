magic
tech gf180mcuD
magscale 1 10
timestamp 1757514455
<< nwell >>
rect -1250 -3370 1250 3370
<< pmos >>
rect -1000 1160 1000 3160
rect -1000 -1024 1000 976
rect -1000 -3208 1000 -1208
<< pdiff >>
rect -1088 3147 -1000 3160
rect -1088 1173 -1075 3147
rect -1029 1173 -1000 3147
rect -1088 1160 -1000 1173
rect 1000 3147 1088 3160
rect 1000 1173 1029 3147
rect 1075 1173 1088 3147
rect 1000 1160 1088 1173
rect -1088 963 -1000 976
rect -1088 -1011 -1075 963
rect -1029 -1011 -1000 963
rect -1088 -1024 -1000 -1011
rect 1000 963 1088 976
rect 1000 -1011 1029 963
rect 1075 -1011 1088 963
rect 1000 -1024 1088 -1011
rect -1088 -1221 -1000 -1208
rect -1088 -3195 -1075 -1221
rect -1029 -3195 -1000 -1221
rect -1088 -3208 -1000 -3195
rect 1000 -1221 1088 -1208
rect 1000 -3195 1029 -1221
rect 1075 -3195 1088 -1221
rect 1000 -3208 1088 -3195
<< pdiffc >>
rect -1075 1173 -1029 3147
rect 1029 1173 1075 3147
rect -1075 -1011 -1029 963
rect 1029 -1011 1075 963
rect -1075 -3195 -1029 -1221
rect 1029 -3195 1075 -1221
<< nsubdiff >>
rect -1226 3274 1226 3346
rect -1226 3230 -1154 3274
rect -1226 -3230 -1213 3230
rect -1167 -3230 -1154 3230
rect 1154 3230 1226 3274
rect -1226 -3274 -1154 -3230
rect 1154 -3230 1167 3230
rect 1213 -3230 1226 3230
rect 1154 -3274 1226 -3230
rect -1226 -3287 1226 -3274
rect -1226 -3333 -1110 -3287
rect 1110 -3333 1226 -3287
rect -1226 -3346 1226 -3333
<< nsubdiffcont >>
rect -1213 -3230 -1167 3230
rect 1167 -3230 1213 3230
rect -1110 -3333 1110 -3287
<< polysilicon >>
rect -1000 3239 1000 3252
rect -1000 3193 -987 3239
rect 987 3193 1000 3239
rect -1000 3160 1000 3193
rect -1000 1116 1000 1160
rect -1000 1055 1000 1068
rect -1000 1009 -987 1055
rect 987 1009 1000 1055
rect -1000 976 1000 1009
rect -1000 -1068 1000 -1024
rect -1000 -1129 1000 -1116
rect -1000 -1175 -987 -1129
rect 987 -1175 1000 -1129
rect -1000 -1208 1000 -1175
rect -1000 -3252 1000 -3208
<< polycontact >>
rect -987 3193 987 3239
rect -987 1009 987 1055
rect -987 -1175 987 -1129
<< metal1 >>
rect -1213 3287 1213 3333
rect -1213 3230 -1167 3287
rect -998 3193 -987 3239
rect 987 3193 998 3239
rect 1167 3230 1213 3287
rect -1075 3147 -1029 3158
rect -1075 1162 -1029 1173
rect 1029 3147 1075 3158
rect 1029 1162 1075 1173
rect -998 1009 -987 1055
rect 987 1009 998 1055
rect -1075 963 -1029 974
rect -1075 -1022 -1029 -1011
rect 1029 963 1075 974
rect 1029 -1022 1075 -1011
rect -998 -1175 -987 -1129
rect 987 -1175 998 -1129
rect -1075 -1221 -1029 -1210
rect -1075 -3206 -1029 -3195
rect 1029 -1221 1075 -1210
rect 1029 -3206 1075 -3195
rect -1213 -3287 -1167 -3230
rect 1167 -3287 1213 -3230
rect -1213 -3333 -1110 -3287
rect 1110 -3333 1213 -3287
<< properties >>
string FIXED_BBOX -1190 -3310 1190 3310
string gencell pfet_03v3
string library gf180mcu
string parameters w 10 l 10 m 3 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {pfet_03v3 pfet_06v0}
<< end >>
