magic
tech gf180mcuD
magscale 1 10
timestamp 1757217098
<< nwell >>
rect -10911 2167 1726 2169
rect -10941 -311 1726 2167
<< pwell >>
rect 1760 -311 21619 2158
<< nmos >>
rect 2147 0 2203 1600
rect 2315 0 2371 1600
rect 2486 0 2542 1600
rect 2654 0 2710 1600
rect 2825 0 2881 1600
rect 2993 0 3049 1600
rect 3164 0 3220 1600
rect 3332 0 3388 1600
rect 3504 0 3560 1600
rect 3672 0 3728 1600
rect 3843 0 3899 1600
rect 4011 0 4067 1600
rect 4182 0 4238 1600
rect 4350 0 4406 1600
rect 4521 0 4577 1600
rect 4689 0 4745 1600
rect 5061 0 5117 1600
rect 5229 0 5285 1600
rect 5400 0 5456 1600
rect 5568 0 5624 1600
rect 5739 0 5795 1600
rect 5907 0 5963 1600
rect 6078 0 6134 1600
rect 6246 0 6302 1600
rect 6418 0 6474 1600
rect 6586 0 6642 1600
rect 6757 0 6813 1600
rect 6925 0 6981 1600
rect 7096 0 7152 1600
rect 7264 0 7320 1600
rect 7435 0 7491 1600
rect 7603 0 7659 1600
rect 7774 0 7830 1600
rect 7942 0 7998 1600
rect 8113 0 8169 1600
rect 8281 0 8337 1600
rect 8452 0 8508 1600
rect 8620 0 8676 1600
rect 8791 0 8847 1600
rect 8959 0 9015 1600
rect 9131 0 9187 1600
rect 9299 0 9355 1600
rect 9470 0 9526 1600
rect 9638 0 9694 1600
rect 9809 0 9865 1600
rect 9977 0 10033 1600
rect 10148 0 10204 1600
rect 10316 0 10372 1600
rect 10675 0 10731 1600
rect 10843 0 10899 1600
rect 11014 0 11070 1600
rect 11182 0 11238 1600
rect 11353 0 11409 1600
rect 11521 0 11577 1600
rect 11692 0 11748 1600
rect 11860 0 11916 1600
rect 12032 0 12088 1600
rect 12200 0 12256 1600
rect 12371 0 12427 1600
rect 12539 0 12595 1600
rect 12710 0 12766 1600
rect 12878 0 12934 1600
rect 13049 0 13105 1600
rect 13217 0 13273 1600
rect 13575 0 13631 1600
rect 13743 0 13799 1600
rect 13914 0 13970 1600
rect 14082 0 14138 1600
rect 14253 0 14309 1600
rect 14421 0 14477 1600
rect 14592 0 14648 1600
rect 14760 0 14816 1600
rect 15115 0 15171 1600
rect 15283 0 15339 1600
rect 15454 0 15510 1600
rect 15622 0 15678 1600
rect 15985 0 16041 1600
rect 16153 0 16209 1600
rect 16525 0 16581 1600
rect 16693 0 16749 1600
rect 16864 0 16920 1600
rect 17032 0 17088 1600
rect 17203 0 17259 1600
rect 17371 0 17427 1600
rect 17542 0 17598 1600
rect 17904 800 17960 1600
rect 18286 1200 18342 1600
rect 18457 1200 18513 1600
rect 18834 1200 18890 1600
rect 19005 1200 19061 1600
rect 19395 1200 19451 1600
rect 19566 1200 19622 1600
rect 19944 1200 20000 1600
rect 20115 1200 20171 1600
rect 20790 1130 20846 1730
rect 18373 -11 18429 789
rect 18544 -11 18600 789
rect 18885 -11 18941 789
rect 19056 -11 19112 789
rect 19404 -11 19460 789
rect 19575 -11 19631 789
rect 19924 -11 19980 789
rect 20095 -11 20151 789
rect 20456 -11 20512 789
rect 20627 -11 20683 789
rect 20974 -11 21030 789
rect 21145 -11 21201 789
<< pmos >>
rect -10481 0 -10425 1600
rect -10315 0 -10259 1600
rect -10150 0 -10094 1600
rect -9984 0 -9928 1600
rect -9819 0 -9763 1600
rect -9653 0 -9597 1600
rect -9488 0 -9432 1600
rect -9322 0 -9266 1600
rect -9155 0 -9099 1600
rect -8989 0 -8933 1600
rect -8824 0 -8768 1600
rect -8658 0 -8602 1600
rect -8493 0 -8437 1600
rect -8327 0 -8271 1600
rect -8162 0 -8106 1600
rect -7996 0 -7940 1600
rect -7830 0 -7774 1600
rect -7664 0 -7608 1600
rect -7499 0 -7443 1600
rect -7333 0 -7277 1600
rect -7168 0 -7112 1600
rect -7002 0 -6946 1600
rect -6837 0 -6781 1600
rect -6671 0 -6615 1600
rect -6504 0 -6448 1600
rect -6338 0 -6282 1600
rect -6173 0 -6117 1600
rect -6007 0 -5951 1600
rect -5842 0 -5786 1600
rect -5676 0 -5620 1600
rect -5511 0 -5455 1600
rect -5345 0 -5289 1600
rect -5178 0 -5122 1600
rect -5012 0 -4956 1600
rect -4847 0 -4791 1600
rect -4681 0 -4625 1600
rect -4516 0 -4460 1600
rect -4350 0 -4294 1600
rect -4185 0 -4129 1600
rect -4019 0 -3963 1600
rect -3852 0 -3796 1600
rect -3686 0 -3630 1600
rect -3521 0 -3465 1600
rect -3355 0 -3299 1600
rect -3190 0 -3134 1600
rect -3024 0 -2968 1600
rect -2859 0 -2803 1600
rect -2693 0 -2637 1600
rect -2529 0 -2473 1600
rect -2363 0 -2307 1600
rect -2198 0 -2142 1600
rect -2032 0 -1976 1600
rect -1867 0 -1811 1600
rect -1701 0 -1645 1600
rect -1536 0 -1480 1600
rect -1370 0 -1314 1600
rect -1204 0 -1148 1600
rect -1038 0 -982 1600
rect -873 0 -817 1600
rect -707 0 -651 1600
rect -542 0 -486 1600
rect -376 0 -320 1600
rect 0 0 56 1600
rect 166 0 222 1600
rect 553 0 609 1600
rect 719 0 775 1600
rect 1122 0 1178 1600
rect 1288 0 1344 1600
<< ndiff >>
rect 20693 1699 20790 1730
rect 2036 1559 2147 1600
rect 2036 40 2068 1559
rect 2114 40 2147 1559
rect 2036 0 2147 40
rect 2203 1559 2315 1600
rect 2203 40 2240 1559
rect 2286 40 2315 1559
rect 2203 0 2315 40
rect 2371 1559 2486 1600
rect 2371 40 2408 1559
rect 2454 40 2486 1559
rect 2371 0 2486 40
rect 2542 1559 2654 1600
rect 2542 40 2579 1559
rect 2625 40 2654 1559
rect 2542 0 2654 40
rect 2710 1559 2825 1600
rect 2710 40 2747 1559
rect 2793 40 2825 1559
rect 2710 0 2825 40
rect 2881 1559 2993 1600
rect 2881 40 2918 1559
rect 2964 40 2993 1559
rect 2881 0 2993 40
rect 3049 1559 3164 1600
rect 3049 40 3086 1559
rect 3132 40 3164 1559
rect 3049 0 3164 40
rect 3220 1559 3332 1600
rect 3220 40 3257 1559
rect 3303 40 3332 1559
rect 3220 0 3332 40
rect 3388 1559 3504 1600
rect 3388 40 3425 1559
rect 3471 40 3504 1559
rect 3388 0 3504 40
rect 3560 1559 3672 1600
rect 3560 40 3597 1559
rect 3643 40 3672 1559
rect 3560 0 3672 40
rect 3728 1559 3843 1600
rect 3728 40 3765 1559
rect 3811 40 3843 1559
rect 3728 0 3843 40
rect 3899 1559 4011 1600
rect 3899 40 3936 1559
rect 3982 40 4011 1559
rect 3899 0 4011 40
rect 4067 1559 4182 1600
rect 4067 40 4104 1559
rect 4150 40 4182 1559
rect 4067 0 4182 40
rect 4238 1559 4350 1600
rect 4238 40 4275 1559
rect 4321 40 4350 1559
rect 4238 0 4350 40
rect 4406 1559 4521 1600
rect 4406 40 4443 1559
rect 4489 40 4521 1559
rect 4406 0 4521 40
rect 4577 1559 4689 1600
rect 4577 40 4614 1559
rect 4660 40 4689 1559
rect 4577 0 4689 40
rect 4745 1559 4860 1600
rect 4745 40 4782 1559
rect 4828 40 4860 1559
rect 4745 0 4860 40
rect 4950 1559 5061 1600
rect 4950 40 4982 1559
rect 5028 40 5061 1559
rect 4950 0 5061 40
rect 5117 1559 5229 1600
rect 5117 40 5154 1559
rect 5200 40 5229 1559
rect 5117 0 5229 40
rect 5285 1559 5400 1600
rect 5285 40 5322 1559
rect 5368 40 5400 1559
rect 5285 0 5400 40
rect 5456 1559 5568 1600
rect 5456 40 5493 1559
rect 5539 40 5568 1559
rect 5456 0 5568 40
rect 5624 1559 5739 1600
rect 5624 40 5661 1559
rect 5707 40 5739 1559
rect 5624 0 5739 40
rect 5795 1559 5907 1600
rect 5795 40 5832 1559
rect 5878 40 5907 1559
rect 5795 0 5907 40
rect 5963 1559 6078 1600
rect 5963 40 6000 1559
rect 6046 40 6078 1559
rect 5963 0 6078 40
rect 6134 1559 6246 1600
rect 6134 40 6171 1559
rect 6217 40 6246 1559
rect 6134 0 6246 40
rect 6302 1559 6418 1600
rect 6302 40 6339 1559
rect 6385 40 6418 1559
rect 6302 0 6418 40
rect 6474 1559 6586 1600
rect 6474 40 6511 1559
rect 6557 40 6586 1559
rect 6474 0 6586 40
rect 6642 1559 6757 1600
rect 6642 40 6679 1559
rect 6725 40 6757 1559
rect 6642 0 6757 40
rect 6813 1559 6925 1600
rect 6813 40 6850 1559
rect 6896 40 6925 1559
rect 6813 0 6925 40
rect 6981 1559 7096 1600
rect 6981 40 7018 1559
rect 7064 40 7096 1559
rect 6981 0 7096 40
rect 7152 1559 7264 1600
rect 7152 40 7189 1559
rect 7235 40 7264 1559
rect 7152 0 7264 40
rect 7320 1559 7435 1600
rect 7320 40 7357 1559
rect 7403 40 7435 1559
rect 7320 0 7435 40
rect 7491 1559 7603 1600
rect 7491 40 7528 1559
rect 7574 40 7603 1559
rect 7491 0 7603 40
rect 7659 1559 7774 1600
rect 7659 40 7696 1559
rect 7742 40 7774 1559
rect 7659 0 7774 40
rect 7830 1559 7942 1600
rect 7830 40 7867 1559
rect 7913 40 7942 1559
rect 7830 0 7942 40
rect 7998 1559 8113 1600
rect 7998 40 8035 1559
rect 8081 40 8113 1559
rect 7998 0 8113 40
rect 8169 1559 8281 1600
rect 8169 40 8206 1559
rect 8252 40 8281 1559
rect 8169 0 8281 40
rect 8337 1559 8452 1600
rect 8337 40 8374 1559
rect 8420 40 8452 1559
rect 8337 0 8452 40
rect 8508 1559 8620 1600
rect 8508 40 8545 1559
rect 8591 40 8620 1559
rect 8508 0 8620 40
rect 8676 1559 8791 1600
rect 8676 40 8713 1559
rect 8759 40 8791 1559
rect 8676 0 8791 40
rect 8847 1559 8959 1600
rect 8847 40 8884 1559
rect 8930 40 8959 1559
rect 8847 0 8959 40
rect 9015 1559 9131 1600
rect 9015 40 9052 1559
rect 9098 40 9131 1559
rect 9015 0 9131 40
rect 9187 1559 9299 1600
rect 9187 40 9224 1559
rect 9270 40 9299 1559
rect 9187 0 9299 40
rect 9355 1559 9470 1600
rect 9355 40 9392 1559
rect 9438 40 9470 1559
rect 9355 0 9470 40
rect 9526 1559 9638 1600
rect 9526 40 9563 1559
rect 9609 40 9638 1559
rect 9526 0 9638 40
rect 9694 1559 9809 1600
rect 9694 40 9731 1559
rect 9777 40 9809 1559
rect 9694 0 9809 40
rect 9865 1559 9977 1600
rect 9865 40 9902 1559
rect 9948 40 9977 1559
rect 9865 0 9977 40
rect 10033 1559 10148 1600
rect 10033 40 10070 1559
rect 10116 40 10148 1559
rect 10033 0 10148 40
rect 10204 1559 10316 1600
rect 10204 40 10241 1559
rect 10287 40 10316 1559
rect 10204 0 10316 40
rect 10372 1559 10487 1600
rect 10372 40 10409 1559
rect 10455 40 10487 1559
rect 10372 0 10487 40
rect 10560 1559 10675 1600
rect 10560 40 10597 1559
rect 10643 40 10675 1559
rect 10560 0 10675 40
rect 10731 1559 10843 1600
rect 10731 40 10768 1559
rect 10814 40 10843 1559
rect 10731 0 10843 40
rect 10899 1559 11014 1600
rect 10899 40 10936 1559
rect 10982 40 11014 1559
rect 10899 0 11014 40
rect 11070 1559 11182 1600
rect 11070 40 11107 1559
rect 11153 40 11182 1559
rect 11070 0 11182 40
rect 11238 1559 11353 1600
rect 11238 40 11275 1559
rect 11321 40 11353 1559
rect 11238 0 11353 40
rect 11409 1559 11521 1600
rect 11409 40 11446 1559
rect 11492 40 11521 1559
rect 11409 0 11521 40
rect 11577 1559 11692 1600
rect 11577 40 11614 1559
rect 11660 40 11692 1559
rect 11577 0 11692 40
rect 11748 1559 11860 1600
rect 11748 40 11785 1559
rect 11831 40 11860 1559
rect 11748 0 11860 40
rect 11916 1559 12032 1600
rect 11916 40 11953 1559
rect 11999 40 12032 1559
rect 11916 0 12032 40
rect 12088 1559 12200 1600
rect 12088 40 12125 1559
rect 12171 40 12200 1559
rect 12088 0 12200 40
rect 12256 1559 12371 1600
rect 12256 40 12293 1559
rect 12339 40 12371 1559
rect 12256 0 12371 40
rect 12427 1559 12539 1600
rect 12427 40 12464 1559
rect 12510 40 12539 1559
rect 12427 0 12539 40
rect 12595 1559 12710 1600
rect 12595 40 12632 1559
rect 12678 40 12710 1559
rect 12595 0 12710 40
rect 12766 1559 12878 1600
rect 12766 40 12803 1559
rect 12849 40 12878 1559
rect 12766 0 12878 40
rect 12934 1559 13049 1600
rect 12934 40 12971 1559
rect 13017 40 13049 1559
rect 12934 0 13049 40
rect 13105 1559 13217 1600
rect 13105 40 13142 1559
rect 13188 40 13217 1559
rect 13105 0 13217 40
rect 13273 1559 13388 1600
rect 13273 40 13310 1559
rect 13356 40 13388 1559
rect 13273 0 13388 40
rect 13460 1559 13575 1600
rect 13460 40 13496 1559
rect 13542 40 13575 1559
rect 13460 0 13575 40
rect 13631 1559 13743 1600
rect 13631 40 13668 1559
rect 13714 40 13743 1559
rect 13631 0 13743 40
rect 13799 1559 13914 1600
rect 13799 40 13836 1559
rect 13882 40 13914 1559
rect 13799 0 13914 40
rect 13970 1559 14082 1600
rect 13970 40 14007 1559
rect 14053 40 14082 1559
rect 13970 0 14082 40
rect 14138 1559 14253 1600
rect 14138 40 14175 1559
rect 14221 40 14253 1559
rect 14138 0 14253 40
rect 14309 1559 14421 1600
rect 14309 40 14346 1559
rect 14392 40 14421 1559
rect 14309 0 14421 40
rect 14477 1559 14592 1600
rect 14477 40 14514 1559
rect 14560 40 14592 1559
rect 14477 0 14592 40
rect 14648 1559 14760 1600
rect 14648 40 14685 1559
rect 14731 40 14760 1559
rect 14648 0 14760 40
rect 14816 1559 14931 1600
rect 14816 40 14853 1559
rect 14899 40 14931 1559
rect 14816 0 14931 40
rect 15000 1559 15115 1600
rect 15000 40 15037 1559
rect 15083 40 15115 1559
rect 15000 0 15115 40
rect 15171 1559 15283 1600
rect 15171 40 15208 1559
rect 15254 40 15283 1559
rect 15171 0 15283 40
rect 15339 1559 15454 1600
rect 15339 40 15376 1559
rect 15422 40 15454 1559
rect 15339 0 15454 40
rect 15510 1559 15622 1600
rect 15510 40 15547 1559
rect 15593 40 15622 1559
rect 15510 0 15622 40
rect 15678 1559 15793 1600
rect 15678 40 15715 1559
rect 15761 40 15793 1559
rect 15678 0 15793 40
rect 15870 1559 15985 1600
rect 15870 40 15907 1559
rect 15953 40 15985 1559
rect 15870 0 15985 40
rect 16041 1559 16153 1600
rect 16041 40 16078 1559
rect 16124 40 16153 1559
rect 16041 0 16153 40
rect 16209 1559 16324 1600
rect 16209 40 16246 1559
rect 16292 40 16324 1559
rect 16209 0 16324 40
rect 16410 1559 16525 1600
rect 16410 40 16447 1559
rect 16493 40 16525 1559
rect 16410 0 16525 40
rect 16581 1559 16693 1600
rect 16581 40 16618 1559
rect 16664 40 16693 1559
rect 16581 0 16693 40
rect 16749 1559 16864 1600
rect 16749 40 16786 1559
rect 16832 40 16864 1559
rect 16749 0 16864 40
rect 16920 1559 17032 1600
rect 16920 40 16957 1559
rect 17003 40 17032 1559
rect 16920 0 17032 40
rect 17088 1559 17203 1600
rect 17088 40 17125 1559
rect 17171 40 17203 1559
rect 17088 0 17203 40
rect 17259 1559 17371 1600
rect 17259 40 17296 1559
rect 17342 40 17371 1559
rect 17259 0 17371 40
rect 17427 1559 17542 1600
rect 17427 40 17464 1559
rect 17510 40 17542 1559
rect 17427 0 17542 40
rect 17598 1559 17713 1600
rect 17598 40 17635 1559
rect 17681 40 17713 1559
rect 17789 1559 17904 1600
rect 17789 830 17826 1559
rect 17872 830 17904 1559
rect 17789 800 17904 830
rect 17960 1559 18075 1600
rect 17960 830 17997 1559
rect 18043 830 18075 1559
rect 18171 1559 18286 1600
rect 18171 1241 18208 1559
rect 18254 1241 18286 1559
rect 18171 1200 18286 1241
rect 18342 1559 18457 1600
rect 18342 1240 18379 1559
rect 18425 1240 18457 1559
rect 18342 1200 18457 1240
rect 18513 1559 18627 1600
rect 18513 1240 18550 1559
rect 18596 1240 18627 1559
rect 18513 1200 18627 1240
rect 18721 1559 18834 1600
rect 18721 1240 18758 1559
rect 18804 1240 18834 1559
rect 18721 1200 18834 1240
rect 18890 1559 19005 1600
rect 18890 1240 18927 1559
rect 18973 1240 19005 1559
rect 18890 1200 19005 1240
rect 19061 1559 19176 1600
rect 19061 1240 19098 1559
rect 19144 1240 19176 1559
rect 19061 1200 19176 1240
rect 19282 1559 19395 1600
rect 19282 1240 19319 1559
rect 19365 1240 19395 1559
rect 19282 1200 19395 1240
rect 19451 1559 19566 1600
rect 19451 1240 19488 1559
rect 19534 1240 19566 1559
rect 19451 1200 19566 1240
rect 19622 1559 19737 1600
rect 19622 1240 19659 1559
rect 19705 1240 19737 1559
rect 19622 1200 19737 1240
rect 19831 1559 19944 1600
rect 19831 1240 19868 1559
rect 19914 1240 19944 1559
rect 19831 1200 19944 1240
rect 20000 1559 20115 1600
rect 20000 1240 20037 1559
rect 20083 1240 20115 1559
rect 20000 1200 20115 1240
rect 20171 1559 20286 1600
rect 20171 1240 20208 1559
rect 20254 1240 20286 1559
rect 20171 1200 20286 1240
rect 20693 1160 20708 1699
rect 20759 1160 20790 1699
rect 20693 1130 20790 1160
rect 20846 1699 20942 1730
rect 20846 1160 20875 1699
rect 20926 1160 20942 1699
rect 20846 1130 20942 1160
rect 17960 800 18075 830
rect 17598 0 17713 40
rect 18258 748 18373 789
rect 18258 19 18295 748
rect 18341 19 18373 748
rect 18258 -11 18373 19
rect 18429 748 18544 789
rect 18429 19 18466 748
rect 18512 19 18544 748
rect 18429 -11 18544 19
rect 18600 748 18713 789
rect 18600 19 18637 748
rect 18683 19 18713 748
rect 18600 -11 18713 19
rect 18772 748 18885 789
rect 18772 19 18809 748
rect 18855 19 18885 748
rect 18772 -11 18885 19
rect 18941 748 19056 789
rect 18941 19 18978 748
rect 19024 19 19056 748
rect 18941 -11 19056 19
rect 19112 748 19227 789
rect 19112 19 19149 748
rect 19195 19 19227 748
rect 19112 -11 19227 19
rect 19291 748 19404 789
rect 19291 718 19328 748
rect 19291 624 19327 718
rect 19291 19 19328 624
rect 19374 19 19404 748
rect 19291 -11 19404 19
rect 19460 748 19575 789
rect 19460 19 19497 748
rect 19543 19 19575 748
rect 19460 -11 19575 19
rect 19631 748 19746 789
rect 19631 530 19668 748
rect 19631 430 19666 530
rect 19631 19 19668 430
rect 19714 19 19746 748
rect 19631 -11 19746 19
rect 19811 748 19924 789
rect 19811 717 19848 748
rect 19811 623 19847 717
rect 19811 19 19848 623
rect 19894 19 19924 748
rect 19811 -11 19924 19
rect 19980 748 20095 789
rect 19980 19 20017 748
rect 20063 19 20095 748
rect 19980 -11 20095 19
rect 20151 748 20266 789
rect 20151 530 20188 748
rect 20151 430 20185 530
rect 20151 19 20188 430
rect 20234 19 20266 748
rect 20151 -11 20266 19
rect 20343 748 20456 789
rect 20343 729 20380 748
rect 20343 635 20375 729
rect 20343 19 20380 635
rect 20426 19 20456 748
rect 20343 -11 20456 19
rect 20512 748 20627 789
rect 20512 19 20549 748
rect 20595 19 20627 748
rect 20512 -11 20627 19
rect 20683 748 20798 789
rect 20683 530 20720 748
rect 20683 430 20716 530
rect 20683 19 20720 430
rect 20766 19 20798 748
rect 20683 -11 20798 19
rect 20861 748 20974 789
rect 20861 724 20898 748
rect 20944 724 20974 748
rect 20861 630 20894 724
rect 20945 630 20974 724
rect 20861 19 20898 630
rect 20944 19 20974 630
rect 20861 -11 20974 19
rect 21030 748 21145 789
rect 21030 19 21067 748
rect 21113 19 21145 748
rect 21030 -11 21145 19
rect 21201 748 21316 789
rect 21201 530 21238 748
rect 21201 430 21233 530
rect 21201 19 21238 430
rect 21284 19 21316 748
rect 21201 -11 21316 19
<< pdiff >>
rect -10592 1560 -10481 1600
rect -10592 40 -10560 1560
rect -10514 40 -10481 1560
rect -10592 0 -10481 40
rect -10425 1560 -10315 1600
rect -10425 40 -10394 1560
rect -10348 40 -10315 1560
rect -10425 0 -10315 40
rect -10259 1560 -10150 1600
rect -10259 40 -10229 1560
rect -10183 40 -10150 1560
rect -10259 0 -10150 40
rect -10094 1560 -9984 1600
rect -10094 40 -10063 1560
rect -10017 236 -9984 1560
rect -10015 125 -9984 236
rect -10017 40 -9984 125
rect -10094 0 -9984 40
rect -9928 1560 -9819 1600
rect -9928 40 -9898 1560
rect -9852 40 -9819 1560
rect -9928 0 -9819 40
rect -9763 1560 -9653 1600
rect -9763 235 -9732 1560
rect -9763 124 -9734 235
rect -9763 40 -9732 124
rect -9686 40 -9653 1560
rect -9763 0 -9653 40
rect -9597 1560 -9488 1600
rect -9597 40 -9567 1560
rect -9521 40 -9488 1560
rect -9597 0 -9488 40
rect -9432 1560 -9322 1600
rect -9432 234 -9401 1560
rect -9432 123 -9403 234
rect -9432 40 -9401 123
rect -9355 40 -9322 1560
rect -9432 0 -9322 40
rect -9266 1560 -9155 1600
rect -9266 40 -9234 1560
rect -9188 40 -9155 1560
rect -9266 0 -9155 40
rect -9099 1560 -8989 1600
rect -9099 237 -9068 1560
rect -9099 126 -9070 237
rect -9099 40 -9068 126
rect -9022 40 -8989 1560
rect -9099 0 -8989 40
rect -8933 1560 -8824 1600
rect -8933 40 -8903 1560
rect -8857 40 -8824 1560
rect -8933 0 -8824 40
rect -8768 1560 -8658 1600
rect -8768 237 -8737 1560
rect -8768 126 -8739 237
rect -8768 40 -8737 126
rect -8691 40 -8658 1560
rect -8768 0 -8658 40
rect -8602 1560 -8493 1600
rect -8602 40 -8572 1560
rect -8526 40 -8493 1560
rect -8602 0 -8493 40
rect -8437 1560 -8327 1600
rect -8437 239 -8406 1560
rect -8437 128 -8408 239
rect -8437 40 -8406 128
rect -8360 40 -8327 1560
rect -8437 0 -8327 40
rect -8271 1560 -8162 1600
rect -8271 40 -8241 1560
rect -8195 40 -8162 1560
rect -8271 0 -8162 40
rect -8106 1560 -7996 1600
rect -8106 241 -8075 1560
rect -8029 241 -7996 1560
rect -8106 130 -8076 241
rect -8028 130 -7996 241
rect -8106 40 -8075 130
rect -8029 40 -7996 130
rect -8106 0 -7996 40
rect -7940 1560 -7830 1600
rect -7940 40 -7909 1560
rect -7863 40 -7830 1560
rect -7940 0 -7830 40
rect -7774 1560 -7664 1600
rect -7774 241 -7743 1560
rect -7774 130 -7745 241
rect -7774 40 -7743 130
rect -7697 40 -7664 1560
rect -7774 0 -7664 40
rect -7608 1560 -7499 1600
rect -7608 40 -7578 1560
rect -7532 40 -7499 1560
rect -7608 0 -7499 40
rect -7443 1560 -7333 1600
rect -7443 241 -7412 1560
rect -7366 241 -7333 1560
rect -7443 130 -7413 241
rect -7365 130 -7333 241
rect -7443 40 -7412 130
rect -7366 40 -7333 130
rect -7443 0 -7333 40
rect -7277 1560 -7168 1600
rect -7277 40 -7247 1560
rect -7201 40 -7168 1560
rect -7277 0 -7168 40
rect -7112 1560 -7002 1600
rect -7112 241 -7081 1560
rect -7035 241 -7002 1560
rect -7112 130 -7082 241
rect -7034 130 -7002 241
rect -7112 40 -7081 130
rect -7035 40 -7002 130
rect -7112 0 -7002 40
rect -6946 1560 -6837 1600
rect -6946 40 -6916 1560
rect -6870 40 -6837 1560
rect -6946 0 -6837 40
rect -6781 1560 -6671 1600
rect -6781 241 -6750 1560
rect -6781 130 -6752 241
rect -6781 40 -6750 130
rect -6704 40 -6671 1560
rect -6781 0 -6671 40
rect -6615 1560 -6504 1600
rect -6615 40 -6583 1560
rect -6537 40 -6504 1560
rect -6615 0 -6504 40
rect -6448 1560 -6338 1600
rect -6448 241 -6417 1560
rect -6448 130 -6419 241
rect -6448 40 -6417 130
rect -6371 40 -6338 1560
rect -6448 0 -6338 40
rect -6282 1560 -6173 1600
rect -6282 40 -6252 1560
rect -6206 40 -6173 1560
rect -6282 0 -6173 40
rect -6117 1560 -6007 1600
rect -6117 241 -6086 1560
rect -6117 130 -6088 241
rect -6117 40 -6086 130
rect -6040 40 -6007 1560
rect -6117 0 -6007 40
rect -5951 1560 -5842 1600
rect -5951 40 -5921 1560
rect -5875 40 -5842 1560
rect -5951 0 -5842 40
rect -5786 1560 -5676 1600
rect -5786 40 -5755 1560
rect -5709 251 -5676 1560
rect -5707 140 -5676 251
rect -5709 40 -5676 140
rect -5786 0 -5676 40
rect -5620 1560 -5511 1600
rect -5620 40 -5590 1560
rect -5544 40 -5511 1560
rect -5620 0 -5511 40
rect -5455 1560 -5345 1600
rect -5455 251 -5424 1560
rect -5455 140 -5426 251
rect -5455 40 -5424 140
rect -5378 40 -5345 1560
rect -5455 0 -5345 40
rect -5289 1560 -5178 1600
rect -5289 40 -5257 1560
rect -5211 40 -5178 1560
rect -5289 0 -5178 40
rect -5122 1560 -5012 1600
rect -5122 40 -5091 1560
rect -5045 40 -5012 1560
rect -5122 0 -5012 40
rect -4956 1560 -4847 1600
rect -4956 40 -4926 1560
rect -4880 40 -4847 1560
rect -4956 0 -4847 40
rect -4791 1560 -4681 1600
rect -4791 40 -4760 1560
rect -4714 252 -4681 1560
rect -4712 150 -4681 252
rect -4714 40 -4681 150
rect -4791 0 -4681 40
rect -4625 1560 -4516 1600
rect -4625 40 -4595 1560
rect -4549 40 -4516 1560
rect -4625 0 -4516 40
rect -4460 1560 -4350 1600
rect -4460 252 -4429 1560
rect -4383 252 -4350 1560
rect -4460 150 -4430 252
rect -4382 150 -4350 252
rect -4460 40 -4429 150
rect -4383 40 -4350 150
rect -4460 0 -4350 40
rect -4294 1560 -4185 1600
rect -4294 40 -4264 1560
rect -4218 40 -4185 1560
rect -4294 0 -4185 40
rect -4129 1560 -4019 1600
rect -4129 252 -4098 1560
rect -4129 150 -4100 252
rect -4129 40 -4098 150
rect -4052 40 -4019 1560
rect -4129 0 -4019 40
rect -3963 1560 -3852 1600
rect -3963 40 -3931 1560
rect -3885 40 -3852 1560
rect -3963 0 -3852 40
rect -3796 1560 -3686 1600
rect -3796 252 -3765 1560
rect -3719 252 -3686 1560
rect -3796 150 -3766 252
rect -3718 150 -3686 252
rect -3796 40 -3765 150
rect -3719 40 -3686 150
rect -3796 0 -3686 40
rect -3630 1560 -3521 1600
rect -3630 40 -3600 1560
rect -3554 40 -3521 1560
rect -3630 0 -3521 40
rect -3465 1560 -3355 1600
rect -3465 252 -3434 1560
rect -3388 252 -3355 1560
rect -3465 150 -3435 252
rect -3387 150 -3355 252
rect -3465 40 -3434 150
rect -3388 40 -3355 150
rect -3465 0 -3355 40
rect -3299 1560 -3190 1600
rect -3299 40 -3269 1560
rect -3223 40 -3190 1560
rect -3299 0 -3190 40
rect -3134 1560 -3024 1600
rect -3134 251 -3103 1560
rect -3134 149 -3105 251
rect -3134 40 -3103 149
rect -3057 40 -3024 1560
rect -3134 0 -3024 40
rect -2968 1560 -2859 1600
rect -2968 40 -2938 1560
rect -2892 40 -2859 1560
rect -2968 0 -2859 40
rect -2803 1560 -2693 1600
rect -2803 252 -2772 1560
rect -2803 150 -2774 252
rect -2803 40 -2772 150
rect -2726 40 -2693 1560
rect -2803 0 -2693 40
rect -2637 1560 -2529 1600
rect -2637 40 -2608 1560
rect -2562 40 -2529 1560
rect -2637 0 -2529 40
rect -2473 1560 -2363 1600
rect -2473 252 -2442 1560
rect -2396 252 -2363 1560
rect -2473 150 -2443 252
rect -2395 150 -2363 252
rect -2473 40 -2442 150
rect -2396 40 -2363 150
rect -2473 0 -2363 40
rect -2307 1560 -2198 1600
rect -2307 40 -2277 1560
rect -2231 40 -2198 1560
rect -2307 0 -2198 40
rect -2142 1560 -2032 1600
rect -2142 252 -2111 1560
rect -2065 252 -2032 1560
rect -2142 150 -2112 252
rect -2064 150 -2032 252
rect -2142 40 -2111 150
rect -2065 40 -2032 150
rect -2142 0 -2032 40
rect -1976 1560 -1867 1600
rect -1976 40 -1946 1560
rect -1900 40 -1867 1560
rect -1976 0 -1867 40
rect -1811 1560 -1701 1600
rect -1811 252 -1780 1560
rect -1811 150 -1782 252
rect -1811 40 -1780 150
rect -1734 40 -1701 1560
rect -1811 0 -1701 40
rect -1645 1560 -1536 1600
rect -1645 40 -1615 1560
rect -1569 40 -1536 1560
rect -1645 0 -1536 40
rect -1480 1560 -1370 1600
rect -1480 252 -1449 1560
rect -1403 252 -1370 1560
rect -1480 150 -1450 252
rect -1402 150 -1370 252
rect -1480 40 -1449 150
rect -1403 40 -1370 150
rect -1480 0 -1370 40
rect -1314 1560 -1204 1600
rect -1314 40 -1283 1560
rect -1237 40 -1204 1560
rect -1314 0 -1204 40
rect -1148 1560 -1038 1600
rect -1148 252 -1117 1560
rect -1148 150 -1119 252
rect -1148 40 -1117 150
rect -1071 40 -1038 1560
rect -1148 0 -1038 40
rect -982 1560 -873 1600
rect -982 40 -952 1560
rect -906 40 -873 1560
rect -982 0 -873 40
rect -817 1560 -707 1600
rect -817 252 -786 1560
rect -740 252 -707 1560
rect -817 150 -787 252
rect -739 150 -707 252
rect -817 40 -786 150
rect -740 40 -707 150
rect -817 0 -707 40
rect -651 1560 -542 1600
rect -651 40 -621 1560
rect -575 40 -542 1560
rect -651 0 -542 40
rect -486 1560 -376 1600
rect -486 252 -455 1560
rect -409 252 -376 1560
rect -486 150 -456 252
rect -408 150 -376 252
rect -486 40 -455 150
rect -409 40 -376 150
rect -486 0 -376 40
rect -320 1560 -209 1600
rect -320 40 -289 1560
rect -243 40 -209 1560
rect -320 0 -209 40
rect -111 1560 0 1600
rect -111 252 -79 1560
rect -111 150 -85 252
rect -111 40 -79 150
rect -33 40 0 1560
rect -111 0 0 40
rect 56 1560 166 1600
rect 56 40 87 1560
rect 133 40 166 1560
rect 56 0 166 40
rect 222 1560 333 1600
rect 222 252 253 1560
rect 299 252 333 1560
rect 222 150 251 252
rect 303 150 333 252
rect 222 40 253 150
rect 299 40 333 150
rect 222 0 333 40
rect 442 1560 553 1600
rect 442 252 474 1560
rect 442 150 467 252
rect 442 40 474 150
rect 520 40 553 1560
rect 442 0 553 40
rect 609 1560 719 1600
rect 609 40 640 1560
rect 686 40 719 1560
rect 609 0 719 40
rect 775 1560 886 1600
rect 775 40 806 1560
rect 852 40 886 1560
rect 775 0 886 40
rect 1011 1560 1122 1600
rect 1011 255 1043 1560
rect 1011 150 1041 255
rect 1011 40 1043 150
rect 1089 40 1122 1560
rect 1011 0 1122 40
rect 1178 1560 1288 1600
rect 1178 40 1209 1560
rect 1255 40 1288 1560
rect 1178 0 1288 40
rect 1344 1560 1455 1600
rect 1344 40 1375 1560
rect 1421 255 1455 1560
rect 1423 150 1455 255
rect 1421 40 1455 150
rect 1344 0 1455 40
<< ndiffc >>
rect 2068 40 2114 1559
rect 2240 40 2286 1559
rect 2408 40 2454 1559
rect 2579 40 2625 1559
rect 2747 40 2793 1559
rect 2918 40 2964 1559
rect 3086 40 3132 1559
rect 3257 40 3303 1559
rect 3425 40 3471 1559
rect 3597 40 3643 1559
rect 3765 40 3811 1559
rect 3936 40 3982 1559
rect 4104 40 4150 1559
rect 4275 40 4321 1559
rect 4443 40 4489 1559
rect 4614 40 4660 1559
rect 4782 40 4828 1559
rect 4982 40 5028 1559
rect 5154 40 5200 1559
rect 5322 40 5368 1559
rect 5493 40 5539 1559
rect 5661 40 5707 1559
rect 5832 40 5878 1559
rect 6000 40 6046 1559
rect 6171 40 6217 1559
rect 6339 40 6385 1559
rect 6511 40 6557 1559
rect 6679 40 6725 1559
rect 6850 40 6896 1559
rect 7018 40 7064 1559
rect 7189 40 7235 1559
rect 7357 40 7403 1559
rect 7528 40 7574 1559
rect 7696 40 7742 1559
rect 7867 40 7913 1559
rect 8035 40 8081 1559
rect 8206 40 8252 1559
rect 8374 40 8420 1559
rect 8545 40 8591 1559
rect 8713 40 8759 1559
rect 8884 40 8930 1559
rect 9052 40 9098 1559
rect 9224 40 9270 1559
rect 9392 40 9438 1559
rect 9563 40 9609 1559
rect 9731 40 9777 1559
rect 9902 40 9948 1559
rect 10070 40 10116 1559
rect 10241 40 10287 1559
rect 10409 40 10455 1559
rect 10597 40 10643 1559
rect 10768 40 10814 1559
rect 10936 40 10982 1559
rect 11107 40 11153 1559
rect 11275 40 11321 1559
rect 11446 40 11492 1559
rect 11614 40 11660 1559
rect 11785 40 11831 1559
rect 11953 40 11999 1559
rect 12125 40 12171 1559
rect 12293 40 12339 1559
rect 12464 40 12510 1559
rect 12632 40 12678 1559
rect 12803 40 12849 1559
rect 12971 40 13017 1559
rect 13142 40 13188 1559
rect 13310 40 13356 1559
rect 13496 40 13542 1559
rect 13668 40 13714 1559
rect 13836 40 13882 1559
rect 14007 40 14053 1559
rect 14175 40 14221 1559
rect 14346 40 14392 1559
rect 14514 40 14560 1559
rect 14685 40 14731 1559
rect 14853 40 14899 1559
rect 15037 40 15083 1559
rect 15208 40 15254 1559
rect 15376 40 15422 1559
rect 15547 40 15593 1559
rect 15715 40 15761 1559
rect 15907 40 15953 1559
rect 16078 40 16124 1559
rect 16246 40 16292 1559
rect 16447 40 16493 1559
rect 16618 40 16664 1559
rect 16786 40 16832 1559
rect 16957 40 17003 1559
rect 17125 40 17171 1559
rect 17296 40 17342 1559
rect 17464 40 17510 1559
rect 17635 40 17681 1559
rect 17826 830 17872 1559
rect 17997 830 18043 1559
rect 18208 1241 18254 1559
rect 18379 1240 18425 1559
rect 18550 1240 18596 1559
rect 18758 1240 18804 1559
rect 18927 1240 18973 1559
rect 19098 1240 19144 1559
rect 19319 1240 19365 1559
rect 19488 1240 19534 1559
rect 19659 1240 19705 1559
rect 19868 1240 19914 1559
rect 20037 1240 20083 1559
rect 20208 1240 20254 1559
rect 20708 1160 20759 1699
rect 20875 1160 20926 1699
rect 18295 19 18341 748
rect 18466 19 18512 748
rect 18637 19 18683 748
rect 18809 19 18855 748
rect 18978 19 19024 748
rect 19149 19 19195 748
rect 19328 718 19374 748
rect 19327 624 19374 718
rect 19328 19 19374 624
rect 19497 19 19543 748
rect 19668 530 19714 748
rect 19666 430 19714 530
rect 19668 19 19714 430
rect 19848 717 19894 748
rect 19847 623 19894 717
rect 19848 19 19894 623
rect 20017 19 20063 748
rect 20188 530 20234 748
rect 20185 430 20234 530
rect 20188 19 20234 430
rect 20380 729 20426 748
rect 20375 635 20426 729
rect 20380 19 20426 635
rect 20549 19 20595 748
rect 20720 530 20766 748
rect 20716 430 20766 530
rect 20720 19 20766 430
rect 20898 724 20944 748
rect 20894 630 20945 724
rect 20898 19 20944 630
rect 21067 19 21113 748
rect 21238 530 21284 748
rect 21233 430 21284 530
rect 21238 19 21284 430
<< pdiffc >>
rect -10560 40 -10514 1560
rect -10394 40 -10348 1560
rect -10229 40 -10183 1560
rect -10063 236 -10017 1560
rect -10063 125 -10015 236
rect -10063 40 -10017 125
rect -9898 40 -9852 1560
rect -9732 235 -9686 1560
rect -9734 124 -9686 235
rect -9732 40 -9686 124
rect -9567 40 -9521 1560
rect -9401 234 -9355 1560
rect -9403 123 -9355 234
rect -9401 40 -9355 123
rect -9234 40 -9188 1560
rect -9068 237 -9022 1560
rect -9070 126 -9022 237
rect -9068 40 -9022 126
rect -8903 40 -8857 1560
rect -8737 237 -8691 1560
rect -8739 126 -8691 237
rect -8737 40 -8691 126
rect -8572 40 -8526 1560
rect -8406 239 -8360 1560
rect -8408 128 -8360 239
rect -8406 40 -8360 128
rect -8241 40 -8195 1560
rect -8075 241 -8029 1560
rect -8076 130 -8028 241
rect -8075 40 -8029 130
rect -7909 40 -7863 1560
rect -7743 241 -7697 1560
rect -7745 130 -7697 241
rect -7743 40 -7697 130
rect -7578 40 -7532 1560
rect -7412 241 -7366 1560
rect -7413 130 -7365 241
rect -7412 40 -7366 130
rect -7247 40 -7201 1560
rect -7081 241 -7035 1560
rect -7082 130 -7034 241
rect -7081 40 -7035 130
rect -6916 40 -6870 1560
rect -6750 241 -6704 1560
rect -6752 130 -6704 241
rect -6750 40 -6704 130
rect -6583 40 -6537 1560
rect -6417 241 -6371 1560
rect -6419 130 -6371 241
rect -6417 40 -6371 130
rect -6252 40 -6206 1560
rect -6086 241 -6040 1560
rect -6088 130 -6040 241
rect -6086 40 -6040 130
rect -5921 40 -5875 1560
rect -5755 251 -5709 1560
rect -5755 140 -5707 251
rect -5755 40 -5709 140
rect -5590 40 -5544 1560
rect -5424 251 -5378 1560
rect -5426 140 -5378 251
rect -5424 40 -5378 140
rect -5257 40 -5211 1560
rect -5091 40 -5045 1560
rect -4926 40 -4880 1560
rect -4760 252 -4714 1560
rect -4760 150 -4712 252
rect -4760 40 -4714 150
rect -4595 40 -4549 1560
rect -4429 252 -4383 1560
rect -4430 150 -4382 252
rect -4429 40 -4383 150
rect -4264 40 -4218 1560
rect -4098 252 -4052 1560
rect -4100 150 -4052 252
rect -4098 40 -4052 150
rect -3931 40 -3885 1560
rect -3765 252 -3719 1560
rect -3766 150 -3718 252
rect -3765 40 -3719 150
rect -3600 40 -3554 1560
rect -3434 252 -3388 1560
rect -3435 150 -3387 252
rect -3434 40 -3388 150
rect -3269 40 -3223 1560
rect -3103 251 -3057 1560
rect -3105 149 -3057 251
rect -3103 40 -3057 149
rect -2938 40 -2892 1560
rect -2772 252 -2726 1560
rect -2774 150 -2726 252
rect -2772 40 -2726 150
rect -2608 40 -2562 1560
rect -2442 252 -2396 1560
rect -2443 150 -2395 252
rect -2442 40 -2396 150
rect -2277 40 -2231 1560
rect -2111 252 -2065 1560
rect -2112 150 -2064 252
rect -2111 40 -2065 150
rect -1946 40 -1900 1560
rect -1780 252 -1734 1560
rect -1782 150 -1734 252
rect -1780 40 -1734 150
rect -1615 40 -1569 1560
rect -1449 252 -1403 1560
rect -1450 150 -1402 252
rect -1449 40 -1403 150
rect -1283 40 -1237 1560
rect -1117 252 -1071 1560
rect -1119 150 -1071 252
rect -1117 40 -1071 150
rect -952 40 -906 1560
rect -786 252 -740 1560
rect -787 150 -739 252
rect -786 40 -740 150
rect -621 40 -575 1560
rect -455 252 -409 1560
rect -456 150 -408 252
rect -455 40 -409 150
rect -289 40 -243 1560
rect -79 252 -33 1560
rect -85 150 -33 252
rect -79 40 -33 150
rect 87 40 133 1560
rect 253 252 299 1560
rect 251 150 303 252
rect 253 40 299 150
rect 474 252 520 1560
rect 467 150 520 252
rect 474 40 520 150
rect 640 40 686 1560
rect 806 40 852 1560
rect 1043 255 1089 1560
rect 1041 150 1089 255
rect 1043 40 1089 150
rect 1209 40 1255 1560
rect 1375 255 1421 1560
rect 1375 150 1423 255
rect 1375 40 1421 150
<< psubdiff >>
rect 11175 2122 11357 2124
rect 16255 2123 16359 2124
rect 17219 2123 18810 2124
rect 13872 2122 20553 2123
rect 10518 2121 20553 2122
rect 21359 2121 21584 2122
rect 1799 2120 4831 2121
rect 6395 2120 6574 2121
rect 7655 2120 21584 2121
rect 1799 2110 21584 2120
rect 1799 2107 17623 2110
rect 1799 2106 6883 2107
rect 1799 2101 3780 2106
rect 1799 2007 2184 2101
rect 2745 2012 3780 2101
rect 4341 2099 6883 2106
rect 4341 2012 5230 2099
rect 2745 2007 5230 2012
rect 1799 2005 5230 2007
rect 5791 2013 6883 2099
rect 7444 2104 9727 2107
rect 7444 2013 8198 2104
rect 5791 2010 8198 2013
rect 8759 2013 9727 2104
rect 10288 2106 17623 2107
rect 10288 2102 16308 2106
rect 10288 2013 11480 2102
rect 8759 2010 11480 2013
rect 5791 2008 11480 2010
rect 12041 2100 16308 2102
rect 12041 2098 14532 2100
rect 12041 2008 12864 2098
rect 5791 2005 12864 2008
rect 1799 2004 12864 2005
rect 13425 2006 14532 2098
rect 15093 2012 16308 2100
rect 16869 2016 17623 2106
rect 18184 2107 21584 2110
rect 18184 2016 19309 2107
rect 16869 2013 19309 2016
rect 19870 2100 21584 2107
rect 19870 2013 20507 2100
rect 16869 2012 20507 2013
rect 15093 2006 20507 2012
rect 21068 2006 21584 2100
rect 13425 2004 21584 2006
rect 1799 1991 21584 2004
rect 1799 1990 14000 1991
rect 1799 1716 1919 1990
rect 4800 1989 7665 1990
rect 8848 1989 9027 1990
rect 12591 1989 12773 1990
rect 13819 1989 14000 1990
rect 14507 1989 14688 1991
rect 12591 1988 12769 1989
rect 13820 1988 14000 1989
rect 14508 1988 14688 1989
rect 15140 1988 15319 1991
rect 15478 1988 15657 1991
rect 18757 1990 20553 1991
rect 21359 1990 21584 1991
rect 13820 1987 13998 1988
rect 14508 1987 14686 1988
rect 15140 1987 15317 1988
rect 15478 1987 15655 1988
rect 1799 1361 1827 1716
rect 1899 1361 1919 1716
rect 1799 920 1919 1361
rect 1799 565 1824 920
rect 1896 565 1919 920
rect 1799 352 1919 565
rect 1799 -3 1820 352
rect 1892 -3 1919 352
rect 21427 1717 21584 1990
rect 21427 1156 21469 1717
rect 21563 1156 21584 1717
rect 1799 -148 1919 -3
rect 21427 538 21584 1156
rect 21427 -23 21462 538
rect 21556 -23 21584 538
rect 1799 -149 17252 -148
rect 18821 -149 20526 -147
rect 21427 -149 21584 -23
rect 1799 -161 21584 -149
rect 1799 -165 7595 -161
rect 1799 -168 3667 -165
rect 1799 -262 2224 -168
rect 2785 -259 3667 -168
rect 4228 -172 6375 -165
rect 4228 -259 5075 -172
rect 2785 -262 5075 -259
rect 1799 -266 5075 -262
rect 5636 -259 6375 -172
rect 6936 -255 7595 -165
rect 8156 -162 21584 -161
rect 8156 -165 18628 -162
rect 8156 -168 13452 -165
rect 8156 -255 9024 -168
rect 6936 -259 9024 -255
rect 5636 -262 9024 -259
rect 9585 -262 10334 -168
rect 10895 -262 11982 -168
rect 12543 -259 13452 -168
rect 14013 -259 15071 -165
rect 15632 -169 18628 -165
rect 15632 -259 16873 -169
rect 12543 -262 16873 -259
rect 5636 -263 16873 -262
rect 17434 -256 18628 -169
rect 19189 -165 21584 -162
rect 19189 -256 20208 -165
rect 17434 -259 20208 -256
rect 20769 -259 21584 -165
rect 17434 -263 21584 -259
rect 5636 -266 21584 -263
rect 1799 -279 21584 -266
rect 1799 -280 1919 -279
rect 4844 -281 21584 -279
rect 17245 -282 21435 -281
<< nsubdiff >>
rect -10891 2120 1583 2121
rect -10891 2094 1689 2120
rect -10891 2089 -4309 2094
rect -10891 2087 -6214 2089
rect -10891 2024 -10645 2087
rect -10260 2084 -6214 2087
rect -10260 2024 -9736 2084
rect -10891 2021 -9736 2024
rect -9351 2083 -6214 2084
rect -9351 2082 -7244 2083
rect -9351 2021 -8322 2082
rect -10891 2019 -8322 2021
rect -7937 2020 -7244 2082
rect -6859 2026 -6214 2083
rect -5829 2079 -4309 2089
rect -5829 2026 -5186 2079
rect -6859 2020 -5186 2026
rect -7937 2019 -5186 2020
rect -10891 2016 -5186 2019
rect -4801 2031 -4309 2079
rect -3924 2092 1689 2094
rect -3924 2031 -3355 2092
rect -4801 2029 -3355 2031
rect -2970 2091 1689 2092
rect -2970 2029 -2495 2091
rect -4801 2028 -2495 2029
rect -2110 2089 1689 2091
rect -2110 2087 -162 2089
rect -2110 2028 -1528 2087
rect -4801 2024 -1528 2028
rect -1143 2026 -162 2087
rect 223 2026 876 2089
rect 1261 2026 1689 2089
rect -1143 2024 1689 2026
rect -4801 2016 1689 2024
rect -10891 2015 1689 2016
rect -10892 2000 1689 2015
rect -10892 1990 1690 2000
rect -10892 1846 -10768 1990
rect -9281 1988 -7136 1990
rect -6513 1988 -4368 1990
rect -10892 1461 -10868 1846
rect -10805 1461 -10768 1846
rect 1570 1740 1690 1990
rect -10892 1249 -10768 1461
rect -10892 864 -10860 1249
rect -10797 864 -10768 1249
rect -10892 451 -10768 864
rect -10892 66 -10855 451
rect -10792 66 -10768 451
rect -10892 -148 -10768 66
rect 1570 1355 1600 1740
rect 1663 1355 1690 1740
rect 1570 971 1690 1355
rect 1570 586 1599 971
rect 1662 586 1690 971
rect 1570 379 1690 586
rect 1570 -6 1598 379
rect 1661 -6 1690 379
rect 1570 -110 1690 -6
rect 1569 -148 1690 -110
rect -10893 -175 1690 -148
rect -10893 -182 -8567 -175
rect -10893 -245 -10444 -182
rect -10059 -183 -8567 -182
rect -10059 -245 -9441 -183
rect -10893 -246 -9441 -245
rect -9056 -238 -8567 -183
rect -8182 -179 626 -175
rect -8182 -181 -4325 -179
rect -8182 -238 -7658 -181
rect -9056 -244 -7658 -238
rect -7273 -184 -4325 -181
rect -7273 -186 -5464 -184
rect -7273 -244 -6670 -186
rect -9056 -246 -6670 -244
rect -10893 -249 -6670 -246
rect -6285 -247 -5464 -186
rect -5079 -242 -4325 -184
rect -3940 -185 626 -179
rect -3940 -242 -3208 -185
rect -5079 -247 -3208 -242
rect -6285 -248 -3208 -247
rect -2823 -191 -1140 -185
rect -2823 -248 -2261 -191
rect -6285 -249 -2261 -248
rect -10893 -254 -2261 -249
rect -1876 -248 -1140 -191
rect -755 -248 -270 -185
rect 115 -238 626 -185
rect 1011 -238 1690 -175
rect 115 -248 1690 -238
rect -1876 -254 1690 -248
rect -10893 -280 1690 -254
rect -10893 -281 1687 -280
<< psubdiffcont >>
rect 2184 2007 2745 2101
rect 3780 2012 4341 2106
rect 5230 2005 5791 2099
rect 6883 2013 7444 2107
rect 8198 2010 8759 2104
rect 9727 2013 10288 2107
rect 11480 2008 12041 2102
rect 12864 2004 13425 2098
rect 14532 2006 15093 2100
rect 16308 2012 16869 2106
rect 17623 2016 18184 2110
rect 19309 2013 19870 2107
rect 20507 2006 21068 2100
rect 1827 1361 1899 1716
rect 1824 565 1896 920
rect 1820 -3 1892 352
rect 21469 1156 21563 1717
rect 21462 -23 21556 538
rect 2224 -262 2785 -168
rect 3667 -259 4228 -165
rect 5075 -266 5636 -172
rect 6375 -259 6936 -165
rect 7595 -255 8156 -161
rect 9024 -262 9585 -168
rect 10334 -262 10895 -168
rect 11982 -262 12543 -168
rect 13452 -259 14013 -165
rect 15071 -259 15632 -165
rect 16873 -263 17434 -169
rect 18628 -256 19189 -162
rect 20208 -259 20769 -165
<< nsubdiffcont >>
rect -10645 2024 -10260 2087
rect -9736 2021 -9351 2084
rect -8322 2019 -7937 2082
rect -7244 2020 -6859 2083
rect -6214 2026 -5829 2089
rect -5186 2016 -4801 2079
rect -4309 2031 -3924 2094
rect -3355 2029 -2970 2092
rect -2495 2028 -2110 2091
rect -1528 2024 -1143 2087
rect -162 2026 223 2089
rect 876 2026 1261 2089
rect -10868 1461 -10805 1846
rect -10860 864 -10797 1249
rect -10855 66 -10792 451
rect 1600 1355 1663 1740
rect 1599 586 1662 971
rect 1598 -6 1661 379
rect -10444 -245 -10059 -182
rect -9441 -246 -9056 -183
rect -8567 -238 -8182 -175
rect -7658 -244 -7273 -181
rect -6670 -249 -6285 -186
rect -5464 -247 -5079 -184
rect -4325 -242 -3940 -179
rect -3208 -248 -2823 -185
rect -2261 -254 -1876 -191
rect -1140 -248 -755 -185
rect -270 -248 115 -185
rect 626 -238 1011 -175
<< polysilicon >>
rect -7642 1767 -7538 1791
rect -7642 1720 -7618 1767
rect -7645 1703 -7618 1720
rect -7557 1703 -7538 1767
rect -3653 1770 -3549 1794
rect -3653 1723 -3629 1770
rect -3656 1706 -3629 1723
rect -3568 1706 -3549 1770
rect -1925 1768 -1821 1792
rect -1925 1721 -1901 1768
rect -1928 1710 -1901 1721
rect -3656 1704 -3549 1706
rect -2529 1704 -1901 1710
rect -1840 1710 -1821 1768
rect -969 1764 -865 1788
rect -969 1717 -945 1764
rect -972 1710 -945 1717
rect -1840 1704 -1314 1710
rect -7645 1702 -7538 1703
rect -10481 1645 -5289 1702
rect -10481 1600 -10425 1645
rect -10315 1600 -10259 1645
rect -10150 1600 -10094 1645
rect -9984 1600 -9928 1645
rect -9819 1600 -9763 1645
rect -9653 1600 -9597 1645
rect -9488 1600 -9432 1645
rect -9322 1600 -9266 1645
rect -9155 1600 -9099 1645
rect -8989 1600 -8933 1645
rect -8824 1600 -8768 1645
rect -8658 1600 -8602 1645
rect -8493 1600 -8437 1645
rect -8327 1600 -8271 1645
rect -8162 1600 -8106 1645
rect -7996 1600 -7940 1645
rect -7830 1600 -7774 1645
rect -7664 1600 -7608 1645
rect -7499 1600 -7443 1645
rect -7333 1600 -7277 1645
rect -7168 1600 -7112 1645
rect -7002 1600 -6946 1645
rect -6837 1600 -6781 1645
rect -6671 1600 -6615 1645
rect -6504 1600 -6448 1645
rect -6338 1600 -6282 1645
rect -6173 1600 -6117 1645
rect -6007 1600 -5951 1645
rect -5842 1600 -5786 1645
rect -5676 1600 -5620 1645
rect -5511 1600 -5455 1645
rect -5345 1600 -5289 1645
rect -5178 1645 -2637 1704
rect -5178 1600 -5122 1645
rect -5012 1600 -4956 1645
rect -4847 1600 -4791 1645
rect -4681 1600 -4625 1645
rect -4516 1600 -4460 1645
rect -4350 1600 -4294 1645
rect -4185 1600 -4129 1645
rect -4019 1600 -3963 1645
rect -3852 1600 -3796 1645
rect -3686 1600 -3630 1645
rect -3521 1600 -3465 1645
rect -3355 1600 -3299 1645
rect -3190 1600 -3134 1645
rect -3024 1600 -2968 1645
rect -2859 1600 -2803 1645
rect -2693 1600 -2637 1645
rect -2529 1646 -1314 1704
rect -2529 1600 -2473 1646
rect -2363 1600 -2307 1646
rect -2198 1600 -2142 1646
rect -2032 1600 -1976 1646
rect -1867 1600 -1811 1646
rect -1701 1600 -1645 1646
rect -1536 1600 -1480 1646
rect -1370 1600 -1314 1646
rect -1204 1700 -945 1710
rect -884 1710 -865 1764
rect -475 1757 -370 1781
rect -475 1710 -451 1757
rect -884 1700 -651 1710
rect -1204 1648 -651 1700
rect -1204 1600 -1148 1648
rect -1038 1600 -982 1648
rect -873 1600 -817 1648
rect -707 1600 -651 1648
rect -542 1693 -451 1710
rect -390 1710 -370 1757
rect -46 1742 59 1766
rect -390 1693 -320 1710
rect -542 1648 -320 1693
rect -46 1678 -22 1742
rect 39 1678 59 1742
rect -46 1650 59 1678
rect 167 1742 272 1766
rect 167 1678 191 1742
rect 252 1678 272 1742
rect 167 1650 272 1678
rect 505 1743 610 1767
rect 505 1679 529 1743
rect 590 1679 610 1743
rect 505 1651 610 1679
rect 720 1742 825 1766
rect 720 1678 744 1742
rect 805 1678 825 1742
rect -542 1600 -486 1648
rect -376 1600 -320 1648
rect 0 1600 56 1650
rect 166 1600 222 1650
rect 553 1600 609 1651
rect 720 1650 825 1678
rect 1075 1740 1180 1764
rect 1075 1676 1099 1740
rect 1160 1676 1180 1740
rect 719 1600 775 1650
rect 1075 1648 1180 1676
rect 1288 1742 1393 1766
rect 1288 1678 1312 1742
rect 1373 1678 1393 1742
rect 1288 1650 1393 1678
rect 1122 1600 1178 1648
rect 1288 1600 1344 1650
rect -10481 -50 -10425 0
rect -10315 -50 -10259 0
rect -10150 -50 -10094 0
rect -9984 -50 -9928 0
rect -9819 -50 -9763 0
rect -9653 -50 -9597 0
rect -9488 -50 -9432 0
rect -9322 -50 -9266 0
rect -9155 -50 -9099 0
rect -8989 -50 -8933 0
rect -8824 -50 -8768 0
rect -8658 -50 -8602 0
rect -8493 -50 -8437 0
rect -8327 -50 -8271 0
rect -8162 -50 -8106 0
rect -7996 -50 -7940 0
rect -7830 -50 -7774 0
rect -7664 -50 -7608 0
rect -7499 -50 -7443 0
rect -7333 -50 -7277 0
rect -7168 -50 -7112 0
rect -7002 -50 -6946 0
rect -6837 -50 -6781 0
rect -6671 -50 -6615 0
rect -6504 -50 -6448 0
rect -6338 -50 -6282 0
rect -6173 -50 -6117 0
rect -6007 -50 -5951 0
rect -5842 -50 -5786 0
rect -5676 -50 -5620 0
rect -5511 -50 -5455 0
rect -5345 -50 -5289 0
rect -5178 -50 -5122 0
rect -5012 -50 -4956 0
rect -4847 -50 -4791 0
rect -4681 -50 -4625 0
rect -4516 -50 -4460 0
rect -4350 -50 -4294 0
rect -4185 -50 -4129 0
rect -4019 -50 -3963 0
rect -3852 -50 -3796 0
rect -3686 -50 -3630 0
rect -3521 -50 -3465 0
rect -3355 -50 -3299 0
rect -3190 -50 -3134 0
rect -3024 -50 -2968 0
rect -2859 -50 -2803 0
rect -2693 -50 -2637 0
rect -2529 -50 -2473 0
rect -2363 -50 -2307 0
rect -2198 -50 -2142 0
rect -2032 -50 -1976 0
rect -1867 -50 -1811 0
rect -1701 -50 -1645 0
rect -1536 -50 -1480 0
rect -1370 -50 -1314 0
rect -1204 -50 -1148 0
rect -1038 -50 -982 0
rect -873 -50 -817 0
rect -707 -50 -651 0
rect -542 -50 -486 0
rect -376 -50 -320 0
rect 0 -50 56 0
rect 166 -50 222 0
rect 553 -50 609 0
rect 719 -50 775 0
rect 1122 -50 1178 0
rect 1288 -50 1344 0
rect 20768 1857 20880 1870
rect 3221 1782 3399 1801
rect 3221 1712 3258 1782
rect 3370 1712 3399 1782
rect 3221 1700 3399 1712
rect 6396 1782 6574 1801
rect 6396 1712 6433 1782
rect 6545 1712 6574 1782
rect 6396 1700 6574 1712
rect 8849 1781 9027 1800
rect 8849 1711 8886 1781
rect 8998 1711 9027 1781
rect 8849 1700 9027 1711
rect 11175 1784 11353 1803
rect 11175 1714 11212 1784
rect 11324 1714 11353 1784
rect 11175 1703 11353 1714
rect 12591 1780 12769 1799
rect 20768 1798 20781 1857
rect 20865 1798 20880 1857
rect 12591 1710 12628 1780
rect 12740 1710 12769 1780
rect 11175 1700 11357 1703
rect 12591 1700 12769 1710
rect 13820 1779 13998 1798
rect 13820 1709 13857 1779
rect 13969 1709 13998 1779
rect 13820 1701 13998 1709
rect 14508 1779 14686 1798
rect 14508 1709 14545 1779
rect 14657 1709 14686 1779
rect 14508 1701 14686 1709
rect 15140 1779 15317 1798
rect 15140 1709 15176 1779
rect 15288 1709 15317 1779
rect 15140 1701 15317 1709
rect 15478 1779 15655 1798
rect 20768 1781 20880 1798
rect 15478 1709 15514 1779
rect 15626 1709 15655 1779
rect 15478 1701 15655 1709
rect 15930 1748 16042 1761
rect 2147 1650 4745 1700
rect 2147 1600 2203 1650
rect 2315 1600 2371 1650
rect 2486 1600 2542 1650
rect 2654 1600 2710 1650
rect 2825 1600 2881 1650
rect 2993 1600 3049 1650
rect 3164 1600 3220 1650
rect 3332 1600 3388 1650
rect 3504 1600 3560 1650
rect 3672 1600 3728 1650
rect 3843 1600 3899 1650
rect 4011 1600 4067 1650
rect 4182 1600 4238 1650
rect 4350 1600 4406 1650
rect 4521 1600 4577 1650
rect 4689 1600 4745 1650
rect 5061 1650 7659 1700
rect 5061 1600 5117 1650
rect 5229 1600 5285 1650
rect 5400 1600 5456 1650
rect 5568 1600 5624 1650
rect 5739 1600 5795 1650
rect 5907 1600 5963 1650
rect 6078 1600 6134 1650
rect 6246 1600 6302 1650
rect 6418 1600 6474 1650
rect 6586 1600 6642 1650
rect 6757 1600 6813 1650
rect 6925 1600 6981 1650
rect 7096 1600 7152 1650
rect 7264 1600 7320 1650
rect 7435 1600 7491 1650
rect 7603 1600 7659 1650
rect 7774 1650 10372 1700
rect 7774 1600 7830 1650
rect 7942 1600 7998 1650
rect 8113 1600 8169 1650
rect 8281 1600 8337 1650
rect 8452 1600 8508 1650
rect 8620 1600 8676 1650
rect 8791 1600 8847 1650
rect 8959 1600 9015 1650
rect 9131 1600 9187 1650
rect 9299 1600 9355 1650
rect 9470 1600 9526 1650
rect 9638 1600 9694 1650
rect 9809 1600 9865 1650
rect 9977 1600 10033 1650
rect 10148 1600 10204 1650
rect 10316 1600 10372 1650
rect 10675 1649 11916 1700
rect 10675 1600 10731 1649
rect 10843 1600 10899 1649
rect 11014 1600 11070 1649
rect 11182 1600 11238 1649
rect 11353 1600 11409 1649
rect 11521 1600 11577 1649
rect 11692 1600 11748 1649
rect 11860 1600 11916 1649
rect 12032 1649 13273 1700
rect 12032 1600 12088 1649
rect 12200 1600 12256 1649
rect 12371 1600 12427 1649
rect 12539 1600 12595 1649
rect 12710 1600 12766 1649
rect 12878 1600 12934 1649
rect 13049 1600 13105 1649
rect 13217 1600 13273 1649
rect 13575 1649 14138 1701
rect 13575 1600 13631 1649
rect 13743 1600 13799 1649
rect 13914 1600 13970 1649
rect 14082 1600 14138 1649
rect 14253 1649 14816 1701
rect 15140 1700 15320 1701
rect 15478 1700 15658 1701
rect 14253 1600 14309 1649
rect 14421 1600 14477 1649
rect 14592 1600 14648 1649
rect 14760 1600 14816 1649
rect 15115 1649 15339 1700
rect 15115 1600 15171 1649
rect 15283 1600 15339 1649
rect 15454 1649 15678 1700
rect 15930 1689 15943 1748
rect 16027 1689 16042 1748
rect 15930 1670 16042 1689
rect 16153 1748 16265 1761
rect 16153 1689 16166 1748
rect 16250 1689 16265 1748
rect 16725 1750 16887 1766
rect 16725 1696 16752 1750
rect 16870 1696 16887 1750
rect 16725 1691 16887 1696
rect 17235 1746 17397 1762
rect 17235 1692 17262 1746
rect 17380 1692 17397 1746
rect 17235 1691 17397 1692
rect 17527 1741 17616 1771
rect 16153 1670 16265 1689
rect 15454 1600 15510 1649
rect 15622 1600 15678 1649
rect 15985 1600 16041 1670
rect 16153 1600 16209 1670
rect 16525 1649 17088 1691
rect 16525 1600 16581 1649
rect 16693 1600 16749 1649
rect 16864 1600 16920 1649
rect 17032 1600 17088 1649
rect 17203 1649 17427 1691
rect 17203 1600 17259 1649
rect 17371 1600 17427 1649
rect 17527 1673 17542 1741
rect 17599 1673 17616 1741
rect 17527 1648 17616 1673
rect 17889 1741 17978 1771
rect 17889 1673 17904 1741
rect 17961 1673 17978 1741
rect 17889 1648 17978 1673
rect 18259 1741 18348 1771
rect 18259 1673 18274 1741
rect 18331 1673 18348 1741
rect 18259 1648 18348 1673
rect 18431 1741 18520 1771
rect 18431 1673 18446 1741
rect 18503 1673 18520 1741
rect 18431 1648 18520 1673
rect 18803 1741 18892 1771
rect 18803 1673 18818 1741
rect 18875 1673 18892 1741
rect 18803 1648 18892 1673
rect 18976 1741 19065 1771
rect 18976 1673 18991 1741
rect 19048 1673 19065 1741
rect 18976 1648 19065 1673
rect 19364 1741 19453 1771
rect 19364 1673 19379 1741
rect 19436 1673 19453 1741
rect 19364 1648 19453 1673
rect 19537 1741 19626 1770
rect 19537 1673 19552 1741
rect 19609 1673 19626 1741
rect 19537 1648 19626 1673
rect 19913 1741 20002 1770
rect 19913 1673 19928 1741
rect 19985 1673 20002 1741
rect 19913 1648 20002 1673
rect 20086 1741 20175 1770
rect 20086 1673 20101 1741
rect 20158 1673 20175 1741
rect 20790 1730 20846 1781
rect 20086 1648 20175 1673
rect 17542 1600 17598 1648
rect 17904 1600 17960 1648
rect 18286 1600 18342 1648
rect 18457 1600 18513 1648
rect 18834 1600 18890 1648
rect 19005 1600 19061 1648
rect 19395 1600 19451 1648
rect 19566 1600 19622 1648
rect 19944 1600 20000 1648
rect 20115 1600 20171 1648
rect 18286 1150 18342 1200
rect 18457 1150 18513 1200
rect 18834 1150 18890 1200
rect 19005 1150 19061 1200
rect 19395 1150 19451 1200
rect 19566 1150 19622 1200
rect 19944 1150 20000 1200
rect 20115 1150 20171 1200
rect 20790 1080 20846 1130
rect 18344 943 18466 973
rect 18534 955 18640 971
rect 18344 874 18377 943
rect 18440 874 18466 943
rect 18344 835 18466 874
rect 18533 936 18640 955
rect 18533 867 18552 936
rect 18615 867 18640 936
rect 18533 850 18640 867
rect 18534 835 18640 850
rect 18879 935 18970 970
rect 19040 955 19135 970
rect 18879 866 18893 935
rect 18956 866 18970 935
rect 17904 750 17960 800
rect 18373 789 18429 835
rect 18534 834 18629 835
rect 18544 789 18600 834
rect 18879 833 18970 866
rect 19039 936 19135 955
rect 19039 867 19058 936
rect 19121 867 19135 936
rect 19039 850 19135 867
rect 19040 834 19135 850
rect 19398 935 19489 970
rect 19559 955 19654 970
rect 19398 866 19412 935
rect 19475 866 19489 935
rect 19050 833 19112 834
rect 19398 833 19489 866
rect 19558 936 19654 955
rect 19558 867 19577 936
rect 19640 867 19654 936
rect 19558 850 19654 867
rect 19559 834 19654 850
rect 19918 935 20009 970
rect 20079 955 20174 970
rect 19918 866 19932 935
rect 19995 866 20009 935
rect 19569 833 19631 834
rect 19918 833 20009 866
rect 20078 936 20174 955
rect 20078 867 20097 936
rect 20160 867 20174 936
rect 20078 850 20174 867
rect 20079 834 20174 850
rect 20450 935 20541 970
rect 20611 955 20706 970
rect 20450 866 20464 935
rect 20527 866 20541 935
rect 20089 833 20151 834
rect 20450 833 20541 866
rect 20610 936 20706 955
rect 20610 867 20629 936
rect 20692 867 20706 936
rect 20610 850 20706 867
rect 20611 834 20706 850
rect 20968 935 21059 970
rect 21129 955 21224 970
rect 20968 866 20982 935
rect 21045 866 21059 935
rect 20621 833 20683 834
rect 20968 833 21059 866
rect 21128 936 21224 955
rect 21128 867 21147 936
rect 21210 867 21224 936
rect 21128 850 21224 867
rect 21129 834 21224 850
rect 21139 833 21201 834
rect 18885 789 18941 833
rect 19056 789 19112 833
rect 19404 789 19460 833
rect 19575 789 19631 833
rect 19924 789 19980 833
rect 20095 789 20151 833
rect 20456 789 20512 833
rect 20627 789 20683 833
rect 20974 789 21030 833
rect 21145 789 21201 833
rect 2147 -50 2203 0
rect 2315 -50 2371 0
rect 2486 -50 2542 0
rect 2654 -50 2710 0
rect 2825 -50 2881 0
rect 2993 -50 3049 0
rect 3164 -50 3220 0
rect 3332 -50 3388 0
rect 3504 -50 3560 0
rect 3672 -50 3728 0
rect 3843 -50 3899 0
rect 4011 -50 4067 0
rect 4182 -50 4238 0
rect 4350 -50 4406 0
rect 4521 -50 4577 0
rect 4689 -50 4745 0
rect 5061 -50 5117 0
rect 5229 -50 5285 0
rect 5400 -50 5456 0
rect 5568 -50 5624 0
rect 5739 -50 5795 0
rect 5907 -50 5963 0
rect 6078 -50 6134 0
rect 6246 -50 6302 0
rect 6418 -50 6474 0
rect 6586 -50 6642 0
rect 6757 -50 6813 0
rect 6925 -50 6981 0
rect 7096 -50 7152 0
rect 7264 -50 7320 0
rect 7435 -50 7491 0
rect 7603 -50 7659 0
rect 7774 -50 7830 0
rect 7942 -50 7998 0
rect 8113 -50 8169 0
rect 8281 -50 8337 0
rect 8452 -50 8508 0
rect 8620 -50 8676 0
rect 8791 -50 8847 0
rect 8959 -50 9015 0
rect 9131 -50 9187 0
rect 9299 -50 9355 0
rect 9470 -50 9526 0
rect 9638 -50 9694 0
rect 9809 -50 9865 0
rect 9977 -50 10033 0
rect 10148 -50 10204 0
rect 10316 -50 10372 0
rect 10675 -50 10731 0
rect 10843 -50 10899 0
rect 11014 -50 11070 0
rect 11182 -50 11238 0
rect 11353 -50 11409 0
rect 11521 -50 11577 0
rect 11692 -50 11748 0
rect 11860 -50 11916 0
rect 12032 -50 12088 0
rect 12200 -50 12256 0
rect 12371 -50 12427 0
rect 12539 -50 12595 0
rect 12710 -50 12766 0
rect 12878 -50 12934 0
rect 13049 -50 13105 0
rect 13217 -50 13273 0
rect 13575 -50 13631 0
rect 13743 -50 13799 0
rect 13914 -50 13970 0
rect 14082 -50 14138 0
rect 14253 -50 14309 0
rect 14421 -50 14477 0
rect 14592 -50 14648 0
rect 14760 -50 14816 0
rect 15115 -50 15171 0
rect 15283 -50 15339 0
rect 15454 -50 15510 0
rect 15622 -50 15678 0
rect 15985 -50 16041 0
rect 16153 -50 16209 0
rect 16525 -50 16581 0
rect 16693 -50 16749 0
rect 16864 -50 16920 0
rect 17032 -50 17088 0
rect 17203 -50 17259 0
rect 17371 -50 17427 0
rect 17542 -50 17598 0
rect 18373 -60 18429 -11
rect 18544 -60 18600 -11
rect 18885 -60 18941 -11
rect 19056 -60 19112 -11
rect 19404 -60 19460 -11
rect 19575 -60 19631 -11
rect 19924 -60 19980 -11
rect 20095 -60 20151 -11
rect 20456 -60 20512 -11
rect 20627 -60 20683 -11
rect 20974 -60 21030 -11
rect 21145 -60 21201 -11
<< polycontact >>
rect -7618 1703 -7557 1767
rect -3629 1706 -3568 1770
rect -1901 1704 -1840 1768
rect -945 1700 -884 1764
rect -451 1693 -390 1757
rect -22 1678 39 1742
rect 191 1678 252 1742
rect 529 1679 590 1743
rect 744 1678 805 1742
rect 1099 1676 1160 1740
rect 1312 1678 1373 1742
rect 3258 1712 3370 1782
rect 6433 1712 6545 1782
rect 8886 1711 8998 1781
rect 11212 1714 11324 1784
rect 20781 1798 20865 1857
rect 12628 1710 12740 1780
rect 13857 1709 13969 1779
rect 14545 1709 14657 1779
rect 15176 1709 15288 1779
rect 15514 1709 15626 1779
rect 15943 1689 16027 1748
rect 16166 1689 16250 1748
rect 16752 1696 16870 1750
rect 17262 1692 17380 1746
rect 17542 1673 17599 1741
rect 17904 1673 17961 1741
rect 18274 1673 18331 1741
rect 18446 1673 18503 1741
rect 18818 1673 18875 1741
rect 18991 1673 19048 1741
rect 19379 1673 19436 1741
rect 19552 1673 19609 1741
rect 19928 1673 19985 1741
rect 20101 1673 20158 1741
rect 18377 874 18440 943
rect 18552 867 18615 936
rect 18893 866 18956 935
rect 19058 867 19121 936
rect 19412 866 19475 935
rect 19577 867 19640 936
rect 19932 866 19995 935
rect 20097 867 20160 936
rect 20464 866 20527 935
rect 20629 867 20692 936
rect 20982 866 21045 935
rect 21147 867 21210 936
<< metal1 >>
rect 11175 2122 11357 2124
rect 16255 2123 16359 2124
rect 17219 2123 18810 2124
rect 13872 2122 20553 2123
rect 10518 2121 20553 2122
rect 21359 2121 21584 2122
rect -10891 2120 1583 2121
rect 1799 2120 4831 2121
rect 6395 2120 6574 2121
rect 7655 2120 21584 2121
rect -10891 2094 1689 2120
rect -10891 2089 -4309 2094
rect -10891 2087 -6214 2089
rect -10891 2024 -10645 2087
rect -10260 2084 -6214 2087
rect -10260 2024 -9736 2084
rect -10891 2021 -9736 2024
rect -9351 2083 -6214 2084
rect -9351 2082 -7244 2083
rect -9351 2021 -8322 2082
rect -10891 2019 -8322 2021
rect -7937 2020 -7244 2082
rect -6859 2026 -6214 2083
rect -5829 2079 -4309 2089
rect -5829 2026 -5186 2079
rect -6859 2020 -5186 2026
rect -7937 2019 -5186 2020
rect -10891 2016 -5186 2019
rect -4801 2031 -4309 2079
rect -3924 2092 1689 2094
rect -3924 2031 -3355 2092
rect -4801 2029 -3355 2031
rect -2970 2091 1689 2092
rect -2970 2029 -2495 2091
rect -4801 2028 -2495 2029
rect -2110 2089 1689 2091
rect -2110 2087 -162 2089
rect -2110 2028 -1528 2087
rect -4801 2024 -1528 2028
rect -1143 2026 -162 2087
rect 223 2026 876 2089
rect 1261 2026 1689 2089
rect -1143 2024 1689 2026
rect -4801 2016 1689 2024
rect -10891 2015 1689 2016
rect -10892 2000 1689 2015
rect 1799 2110 21584 2120
rect 1799 2107 17623 2110
rect 1799 2106 6883 2107
rect 1799 2101 3780 2106
rect 1799 2007 2184 2101
rect 2745 2012 3780 2101
rect 4341 2099 6883 2106
rect 4341 2012 5230 2099
rect 2745 2007 5230 2012
rect 1799 2005 5230 2007
rect 5791 2013 6883 2099
rect 7444 2104 9727 2107
rect 7444 2013 8198 2104
rect 5791 2010 8198 2013
rect 8759 2013 9727 2104
rect 10288 2106 17623 2107
rect 10288 2102 16308 2106
rect 10288 2013 11480 2102
rect 8759 2010 11480 2013
rect 5791 2008 11480 2010
rect 12041 2100 16308 2102
rect 12041 2098 14532 2100
rect 12041 2008 12864 2098
rect 5791 2005 12864 2008
rect 1799 2004 12864 2005
rect 13425 2006 14532 2098
rect 15093 2012 16308 2100
rect 16869 2016 17623 2106
rect 18184 2107 21584 2110
rect 18184 2016 19309 2107
rect 16869 2013 19309 2016
rect 19870 2100 21584 2107
rect 19870 2013 20507 2100
rect 16869 2012 20507 2013
rect 15093 2006 20507 2012
rect 21068 2006 21584 2100
rect 13425 2004 21584 2006
rect -10892 1990 1690 2000
rect -10892 1846 -10768 1990
rect -9281 1988 -7136 1990
rect -6513 1988 -4368 1990
rect -10892 1461 -10868 1846
rect -10805 1461 -10768 1846
rect -7643 1767 -7538 1792
rect -7643 1703 -7618 1767
rect -7557 1703 -7538 1767
rect -7643 1675 -7538 1703
rect -3654 1770 -3549 1795
rect -3654 1706 -3629 1770
rect -3568 1706 -3549 1770
rect -3654 1678 -3549 1706
rect -1926 1768 -1821 1793
rect -1926 1704 -1901 1768
rect -1840 1704 -1821 1768
rect -1926 1676 -1821 1704
rect -970 1764 -865 1789
rect -970 1700 -945 1764
rect -884 1700 -865 1764
rect -970 1672 -865 1700
rect -476 1757 -371 1782
rect -476 1693 -451 1757
rect -390 1693 -371 1757
rect -476 1665 -371 1693
rect -47 1742 58 1767
rect -47 1678 -22 1742
rect 39 1678 58 1742
rect -47 1650 58 1678
rect 166 1742 271 1767
rect 166 1678 191 1742
rect 252 1678 271 1742
rect 166 1650 271 1678
rect 504 1743 609 1768
rect 504 1679 529 1743
rect 590 1679 609 1743
rect 504 1651 609 1679
rect 719 1742 824 1767
rect 719 1678 744 1742
rect 805 1678 824 1742
rect 719 1650 824 1678
rect 1074 1740 1179 1765
rect 1074 1676 1099 1740
rect 1160 1676 1179 1740
rect 1074 1648 1179 1676
rect 1287 1742 1392 1767
rect 1287 1678 1312 1742
rect 1373 1678 1392 1742
rect 1287 1650 1392 1678
rect 1570 1740 1690 1990
rect -10892 1249 -10768 1461
rect -10892 864 -10860 1249
rect -10797 864 -10768 1249
rect -10892 451 -10768 864
rect -10892 66 -10855 451
rect -10792 66 -10768 451
rect -10892 -148 -10768 66
rect -10570 1560 -10506 1571
rect -10570 1549 -10560 1560
rect -10514 1549 -10506 1560
rect -10570 50 -10561 1549
rect -10509 50 -10506 1549
rect -10570 40 -10560 50
rect -10514 40 -10506 50
rect -10570 30 -10506 40
rect -10401 1560 -10337 1571
rect -10401 40 -10394 1560
rect -10348 1549 -10337 1560
rect -10341 48 -10337 1549
rect -10348 40 -10337 48
rect -10401 30 -10337 40
rect -10239 1560 -10175 1571
rect -10239 1549 -10229 1560
rect -10183 1549 -10175 1560
rect -10239 50 -10230 1549
rect -10178 50 -10175 1549
rect -10239 40 -10229 50
rect -10183 40 -10175 50
rect -10239 30 -10175 40
rect -10070 1560 -10006 1571
rect -10070 40 -10063 1560
rect -10017 1549 -10006 1560
rect -10010 236 -10006 1549
rect -9908 1560 -9844 1571
rect -9908 1549 -9898 1560
rect -9852 1549 -9844 1560
rect -10008 125 -10004 236
rect -10010 48 -10006 125
rect -10017 40 -10006 48
rect -10070 30 -10006 40
rect -9908 50 -9899 1549
rect -9847 50 -9844 1549
rect -9908 40 -9898 50
rect -9852 40 -9844 50
rect -9908 30 -9844 40
rect -9739 1560 -9675 1571
rect -9739 235 -9732 1560
rect -9686 1549 -9675 1560
rect -9739 124 -9734 235
rect -9739 40 -9732 124
rect -9679 48 -9675 1549
rect -9686 40 -9675 48
rect -9739 30 -9675 40
rect -9577 1560 -9513 1571
rect -9577 1549 -9567 1560
rect -9521 1549 -9513 1560
rect -9577 50 -9568 1549
rect -9516 50 -9513 1549
rect -9577 40 -9567 50
rect -9521 40 -9513 50
rect -9577 30 -9513 40
rect -9408 1560 -9344 1571
rect -9408 234 -9401 1560
rect -9355 1549 -9344 1560
rect -9408 123 -9403 234
rect -9408 40 -9401 123
rect -9348 48 -9344 1549
rect -9355 40 -9344 48
rect -9408 30 -9344 40
rect -9244 1560 -9180 1571
rect -9244 1549 -9234 1560
rect -9188 1549 -9180 1560
rect -9244 50 -9235 1549
rect -9183 50 -9180 1549
rect -9244 40 -9234 50
rect -9188 40 -9180 50
rect -9244 30 -9180 40
rect -9075 1560 -9011 1571
rect -9075 237 -9068 1560
rect -9022 1549 -9011 1560
rect -9075 126 -9070 237
rect -9075 40 -9068 126
rect -9015 48 -9011 1549
rect -9022 40 -9011 48
rect -9075 30 -9011 40
rect -8913 1560 -8849 1571
rect -8913 1549 -8903 1560
rect -8857 1549 -8849 1560
rect -8913 50 -8904 1549
rect -8852 50 -8849 1549
rect -8913 40 -8903 50
rect -8857 40 -8849 50
rect -8913 30 -8849 40
rect -8744 1560 -8680 1571
rect -8744 237 -8737 1560
rect -8691 1549 -8680 1560
rect -8744 126 -8739 237
rect -8744 40 -8737 126
rect -8684 48 -8680 1549
rect -8691 40 -8680 48
rect -8744 30 -8680 40
rect -8582 1560 -8518 1571
rect -8582 1549 -8572 1560
rect -8526 1549 -8518 1560
rect -8582 50 -8573 1549
rect -8521 50 -8518 1549
rect -8582 40 -8572 50
rect -8526 40 -8518 50
rect -8582 30 -8518 40
rect -8413 1560 -8349 1571
rect -8413 239 -8406 1560
rect -8360 1549 -8349 1560
rect -8413 128 -8408 239
rect -8413 40 -8406 128
rect -8353 48 -8349 1549
rect -8360 40 -8349 48
rect -8413 30 -8349 40
rect -8251 1560 -8187 1571
rect -8251 1549 -8241 1560
rect -8195 1549 -8187 1560
rect -8251 50 -8242 1549
rect -8190 50 -8187 1549
rect -8251 40 -8241 50
rect -8195 40 -8187 50
rect -8251 30 -8187 40
rect -8082 1560 -8018 1571
rect -8082 241 -8075 1560
rect -8029 1549 -8018 1560
rect -8022 241 -8018 1549
rect -7919 1560 -7855 1571
rect -7919 1549 -7909 1560
rect -7863 1549 -7855 1560
rect -8082 130 -8076 241
rect -8021 130 -8017 241
rect -8082 40 -8075 130
rect -8022 48 -8018 130
rect -8029 40 -8018 48
rect -8082 30 -8018 40
rect -7919 50 -7910 1549
rect -7858 50 -7855 1549
rect -7919 40 -7909 50
rect -7863 40 -7855 50
rect -7919 30 -7855 40
rect -7750 1560 -7686 1571
rect -7750 241 -7743 1560
rect -7697 1549 -7686 1560
rect -7750 130 -7745 241
rect -7750 40 -7743 130
rect -7690 48 -7686 1549
rect -7697 40 -7686 48
rect -7750 30 -7686 40
rect -7588 1560 -7524 1571
rect -7588 1549 -7578 1560
rect -7532 1549 -7524 1560
rect -7588 50 -7579 1549
rect -7527 50 -7524 1549
rect -7588 40 -7578 50
rect -7532 40 -7524 50
rect -7588 30 -7524 40
rect -7419 1560 -7355 1571
rect -7419 241 -7412 1560
rect -7366 1549 -7355 1560
rect -7359 241 -7355 1549
rect -7257 1560 -7193 1571
rect -7257 1549 -7247 1560
rect -7201 1549 -7193 1560
rect -7419 130 -7413 241
rect -7358 130 -7354 241
rect -7419 40 -7412 130
rect -7359 48 -7355 130
rect -7366 40 -7355 48
rect -7419 30 -7355 40
rect -7257 50 -7248 1549
rect -7196 50 -7193 1549
rect -7257 40 -7247 50
rect -7201 40 -7193 50
rect -7257 30 -7193 40
rect -7088 1560 -7024 1571
rect -7088 241 -7081 1560
rect -7035 1549 -7024 1560
rect -7028 241 -7024 1549
rect -6926 1560 -6862 1571
rect -6926 1549 -6916 1560
rect -6870 1549 -6862 1560
rect -7088 130 -7082 241
rect -7027 130 -7023 241
rect -7088 40 -7081 130
rect -7028 48 -7024 130
rect -7035 40 -7024 48
rect -7088 30 -7024 40
rect -6926 50 -6917 1549
rect -6865 50 -6862 1549
rect -6926 40 -6916 50
rect -6870 40 -6862 50
rect -6926 30 -6862 40
rect -6757 1560 -6693 1571
rect -6757 241 -6750 1560
rect -6704 1549 -6693 1560
rect -6757 130 -6752 241
rect -6757 40 -6750 130
rect -6697 48 -6693 1549
rect -6704 40 -6693 48
rect -6757 30 -6693 40
rect -6593 1560 -6529 1571
rect -6593 1549 -6583 1560
rect -6537 1549 -6529 1560
rect -6593 50 -6584 1549
rect -6532 50 -6529 1549
rect -6593 40 -6583 50
rect -6537 40 -6529 50
rect -6593 30 -6529 40
rect -6424 1560 -6360 1571
rect -6424 241 -6417 1560
rect -6371 1549 -6360 1560
rect -6424 130 -6419 241
rect -6424 40 -6417 130
rect -6364 48 -6360 1549
rect -6371 40 -6360 48
rect -6424 30 -6360 40
rect -6262 1560 -6198 1571
rect -6262 1549 -6252 1560
rect -6206 1549 -6198 1560
rect -6262 50 -6253 1549
rect -6201 50 -6198 1549
rect -6262 40 -6252 50
rect -6206 40 -6198 50
rect -6262 30 -6198 40
rect -6093 1560 -6029 1571
rect -6093 241 -6086 1560
rect -6040 1549 -6029 1560
rect -6093 130 -6088 241
rect -6093 40 -6086 130
rect -6033 48 -6029 1549
rect -6040 40 -6029 48
rect -6093 30 -6029 40
rect -5931 1560 -5867 1571
rect -5931 1549 -5921 1560
rect -5875 1549 -5867 1560
rect -5931 50 -5922 1549
rect -5870 50 -5867 1549
rect -5931 40 -5921 50
rect -5875 40 -5867 50
rect -5931 30 -5867 40
rect -5762 1560 -5698 1571
rect -5762 40 -5755 1560
rect -5709 1549 -5698 1560
rect -5702 251 -5698 1549
rect -5600 1560 -5536 1571
rect -5600 1549 -5590 1560
rect -5544 1549 -5536 1560
rect -5700 140 -5696 251
rect -5702 48 -5698 140
rect -5709 40 -5698 48
rect -5762 30 -5698 40
rect -5600 50 -5591 1549
rect -5539 50 -5536 1549
rect -5600 40 -5590 50
rect -5544 40 -5536 50
rect -5600 30 -5536 40
rect -5431 1560 -5367 1571
rect -5431 251 -5424 1560
rect -5378 1549 -5367 1560
rect -5431 140 -5426 251
rect -5431 40 -5424 140
rect -5371 48 -5367 1549
rect -5378 40 -5367 48
rect -5431 30 -5367 40
rect -5267 1560 -5203 1571
rect -5267 1549 -5257 1560
rect -5211 1549 -5203 1560
rect -5267 50 -5258 1549
rect -5206 50 -5203 1549
rect -5267 40 -5257 50
rect -5211 40 -5203 50
rect -5267 30 -5203 40
rect -5098 1560 -5034 1571
rect -5098 40 -5091 1560
rect -5045 1549 -5034 1560
rect -5038 48 -5034 1549
rect -5045 40 -5034 48
rect -5098 30 -5034 40
rect -4936 1560 -4872 1571
rect -4936 1549 -4926 1560
rect -4880 1549 -4872 1560
rect -4936 50 -4927 1549
rect -4875 50 -4872 1549
rect -4936 40 -4926 50
rect -4880 40 -4872 50
rect -4936 30 -4872 40
rect -4767 1560 -4703 1571
rect -4767 40 -4760 1560
rect -4714 1549 -4703 1560
rect -4707 252 -4703 1549
rect -4605 1560 -4541 1571
rect -4605 1549 -4595 1560
rect -4549 1549 -4541 1560
rect -4705 150 -4701 252
rect -4707 48 -4703 150
rect -4714 40 -4703 48
rect -4767 30 -4703 40
rect -4605 50 -4596 1549
rect -4544 50 -4541 1549
rect -4605 40 -4595 50
rect -4549 40 -4541 50
rect -4605 30 -4541 40
rect -4436 1560 -4372 1571
rect -4436 252 -4429 1560
rect -4383 1549 -4372 1560
rect -4376 252 -4372 1549
rect -4274 1560 -4210 1571
rect -4274 1549 -4264 1560
rect -4218 1549 -4210 1560
rect -4436 150 -4430 252
rect -4375 150 -4371 252
rect -4436 40 -4429 150
rect -4376 48 -4372 150
rect -4383 40 -4372 48
rect -4436 30 -4372 40
rect -4274 50 -4265 1549
rect -4213 50 -4210 1549
rect -4274 40 -4264 50
rect -4218 40 -4210 50
rect -4274 30 -4210 40
rect -4105 1560 -4041 1571
rect -4105 252 -4098 1560
rect -4052 1549 -4041 1560
rect -4105 150 -4100 252
rect -4105 40 -4098 150
rect -4045 48 -4041 1549
rect -4052 40 -4041 48
rect -4105 30 -4041 40
rect -3941 1560 -3877 1571
rect -3941 1549 -3931 1560
rect -3885 1549 -3877 1560
rect -3941 50 -3932 1549
rect -3880 50 -3877 1549
rect -3941 40 -3931 50
rect -3885 40 -3877 50
rect -3941 30 -3877 40
rect -3772 1560 -3708 1571
rect -3772 252 -3765 1560
rect -3719 1549 -3708 1560
rect -3712 252 -3708 1549
rect -3610 1560 -3546 1571
rect -3610 1549 -3600 1560
rect -3554 1549 -3546 1560
rect -3772 150 -3766 252
rect -3711 150 -3707 252
rect -3772 40 -3765 150
rect -3712 48 -3708 150
rect -3719 40 -3708 48
rect -3772 30 -3708 40
rect -3610 50 -3601 1549
rect -3549 50 -3546 1549
rect -3610 40 -3600 50
rect -3554 40 -3546 50
rect -3610 30 -3546 40
rect -3441 1560 -3377 1571
rect -3441 252 -3434 1560
rect -3388 1549 -3377 1560
rect -3381 252 -3377 1549
rect -3279 1560 -3215 1571
rect -3279 1549 -3269 1560
rect -3223 1549 -3215 1560
rect -3441 150 -3435 252
rect -3380 150 -3376 252
rect -3441 40 -3434 150
rect -3381 48 -3377 150
rect -3388 40 -3377 48
rect -3441 30 -3377 40
rect -3279 50 -3270 1549
rect -3218 50 -3215 1549
rect -3279 40 -3269 50
rect -3223 40 -3215 50
rect -3279 30 -3215 40
rect -3110 1560 -3046 1571
rect -3110 251 -3103 1560
rect -3057 1549 -3046 1560
rect -3110 149 -3105 251
rect -3110 40 -3103 149
rect -3050 48 -3046 1549
rect -3057 40 -3046 48
rect -3110 30 -3046 40
rect -2948 1560 -2884 1571
rect -2948 1549 -2938 1560
rect -2892 1549 -2884 1560
rect -2948 50 -2939 1549
rect -2887 50 -2884 1549
rect -2948 40 -2938 50
rect -2892 40 -2884 50
rect -2948 30 -2884 40
rect -2779 1560 -2715 1571
rect -2779 252 -2772 1560
rect -2726 1549 -2715 1560
rect -2779 150 -2774 252
rect -2779 40 -2772 150
rect -2719 48 -2715 1549
rect -2726 40 -2715 48
rect -2779 30 -2715 40
rect -2618 1560 -2554 1571
rect -2618 1549 -2608 1560
rect -2562 1549 -2554 1560
rect -2618 50 -2609 1549
rect -2557 50 -2554 1549
rect -2618 40 -2608 50
rect -2562 40 -2554 50
rect -2618 30 -2554 40
rect -2449 1560 -2385 1571
rect -2449 252 -2442 1560
rect -2396 1549 -2385 1560
rect -2389 252 -2385 1549
rect -2287 1560 -2223 1571
rect -2287 1549 -2277 1560
rect -2231 1549 -2223 1560
rect -2449 150 -2443 252
rect -2388 150 -2384 252
rect -2449 40 -2442 150
rect -2389 48 -2385 150
rect -2396 40 -2385 48
rect -2449 30 -2385 40
rect -2287 50 -2278 1549
rect -2226 50 -2223 1549
rect -2287 40 -2277 50
rect -2231 40 -2223 50
rect -2287 30 -2223 40
rect -2118 1560 -2054 1571
rect -2118 252 -2111 1560
rect -2065 1549 -2054 1560
rect -2058 252 -2054 1549
rect -1956 1560 -1892 1571
rect -1956 1549 -1946 1560
rect -1900 1549 -1892 1560
rect -2118 150 -2112 252
rect -2057 150 -2053 252
rect -2118 40 -2111 150
rect -2058 48 -2054 150
rect -2065 40 -2054 48
rect -2118 30 -2054 40
rect -1956 50 -1947 1549
rect -1895 50 -1892 1549
rect -1956 40 -1946 50
rect -1900 40 -1892 50
rect -1956 30 -1892 40
rect -1787 1560 -1723 1571
rect -1787 252 -1780 1560
rect -1734 1549 -1723 1560
rect -1787 150 -1782 252
rect -1787 40 -1780 150
rect -1727 48 -1723 1549
rect -1734 40 -1723 48
rect -1787 30 -1723 40
rect -1625 1560 -1561 1571
rect -1625 1549 -1615 1560
rect -1569 1549 -1561 1560
rect -1625 50 -1616 1549
rect -1564 50 -1561 1549
rect -1625 40 -1615 50
rect -1569 40 -1561 50
rect -1625 30 -1561 40
rect -1456 1560 -1392 1571
rect -1456 252 -1449 1560
rect -1403 1549 -1392 1560
rect -1396 252 -1392 1549
rect -1293 1560 -1229 1571
rect -1293 1549 -1283 1560
rect -1237 1549 -1229 1560
rect -1456 150 -1450 252
rect -1395 150 -1391 252
rect -1456 40 -1449 150
rect -1396 48 -1392 150
rect -1403 40 -1392 48
rect -1456 30 -1392 40
rect -1293 50 -1284 1549
rect -1232 50 -1229 1549
rect -1293 40 -1283 50
rect -1237 40 -1229 50
rect -1293 30 -1229 40
rect -1124 1560 -1060 1571
rect -1124 252 -1117 1560
rect -1071 1549 -1060 1560
rect -1124 150 -1119 252
rect -1124 40 -1117 150
rect -1064 48 -1060 1549
rect -1071 40 -1060 48
rect -1124 30 -1060 40
rect -962 1560 -898 1571
rect -962 1549 -952 1560
rect -906 1549 -898 1560
rect -962 50 -953 1549
rect -901 50 -898 1549
rect -962 40 -952 50
rect -906 40 -898 50
rect -962 30 -898 40
rect -793 1560 -729 1571
rect -793 252 -786 1560
rect -740 1549 -729 1560
rect -733 252 -729 1549
rect -631 1560 -567 1571
rect -631 1549 -621 1560
rect -575 1549 -567 1560
rect -793 150 -787 252
rect -732 150 -728 252
rect -793 40 -786 150
rect -733 48 -729 150
rect -740 40 -729 48
rect -793 30 -729 40
rect -631 50 -622 1549
rect -570 50 -567 1549
rect -631 40 -621 50
rect -575 40 -567 50
rect -631 30 -567 40
rect -462 1560 -398 1571
rect -462 252 -455 1560
rect -409 1549 -398 1560
rect -402 252 -398 1549
rect -296 1560 -232 1571
rect -462 150 -456 252
rect -401 150 -397 252
rect -462 40 -455 150
rect -402 48 -398 150
rect -409 40 -398 48
rect -462 30 -398 40
rect -296 40 -289 1560
rect -243 1549 -232 1560
rect -236 48 -232 1549
rect -89 1560 -25 1571
rect -89 1549 -79 1560
rect -33 1549 -25 1560
rect -89 252 -80 1549
rect -90 150 -85 252
rect -243 40 -232 48
rect -296 30 -232 40
rect -89 50 -80 150
rect -28 50 -25 1549
rect -89 40 -79 50
rect -33 40 -25 50
rect -89 30 -25 40
rect 80 1560 144 1571
rect 80 40 87 1560
rect 133 1549 144 1560
rect 140 48 144 1549
rect 133 40 144 48
rect 80 30 144 40
rect 246 1560 310 1571
rect 246 252 253 1560
rect 299 1549 310 1560
rect 306 252 310 1549
rect 464 1560 528 1571
rect 464 1549 474 1560
rect 520 1549 528 1560
rect 464 252 473 1549
rect 246 150 251 252
rect 308 150 310 252
rect 462 150 467 252
rect 246 40 253 150
rect 306 48 310 150
rect 299 40 310 48
rect 246 30 310 40
rect 464 50 473 150
rect 525 50 528 1549
rect 464 40 474 50
rect 520 40 528 50
rect 464 30 528 40
rect 633 1560 697 1571
rect 633 40 640 1560
rect 686 1549 697 1560
rect 693 48 697 1549
rect 686 40 697 48
rect 633 30 697 40
rect 799 1560 863 1571
rect 799 40 806 1560
rect 852 1549 863 1560
rect 859 48 863 1549
rect 852 40 863 48
rect 799 30 863 40
rect 1033 1560 1097 1571
rect 1033 1549 1043 1560
rect 1089 1549 1097 1560
rect 1033 255 1042 1549
rect 1033 150 1041 255
rect 1033 50 1042 150
rect 1094 255 1097 1549
rect 1202 1560 1266 1571
rect 1094 150 1098 255
rect 1094 50 1097 150
rect 1033 40 1043 50
rect 1089 40 1097 50
rect 1033 30 1097 40
rect 1202 40 1209 1560
rect 1255 1549 1266 1560
rect 1262 48 1266 1549
rect 1255 40 1266 48
rect 1202 30 1266 40
rect 1368 1560 1432 1571
rect 1368 40 1375 1560
rect 1421 1549 1432 1560
rect 1428 48 1432 1549
rect 1421 40 1432 48
rect 1368 30 1432 40
rect 1570 1355 1600 1740
rect 1663 1355 1690 1740
rect 1570 971 1690 1355
rect 1570 586 1599 971
rect 1662 586 1690 971
rect 1570 379 1690 586
rect 1570 -6 1598 379
rect 1661 -6 1690 379
rect 1570 -110 1690 -6
rect 1569 -148 1690 -110
rect -10893 -175 1690 -148
rect -10893 -182 -8567 -175
rect -10893 -245 -10444 -182
rect -10059 -183 -8567 -182
rect -10059 -245 -9441 -183
rect -10893 -246 -9441 -245
rect -9056 -238 -8567 -183
rect -8182 -179 626 -175
rect -8182 -181 -4325 -179
rect -8182 -238 -7658 -181
rect -9056 -244 -7658 -238
rect -7273 -184 -4325 -181
rect -7273 -186 -5464 -184
rect -7273 -244 -6670 -186
rect -9056 -246 -6670 -244
rect -10893 -249 -6670 -246
rect -6285 -247 -5464 -186
rect -5079 -242 -4325 -184
rect -3940 -185 626 -179
rect -3940 -242 -3208 -185
rect -5079 -247 -3208 -242
rect -6285 -248 -3208 -247
rect -2823 -191 -1140 -185
rect -2823 -248 -2261 -191
rect -6285 -249 -2261 -248
rect -10893 -254 -2261 -249
rect -1876 -248 -1140 -191
rect -755 -248 -270 -185
rect 115 -238 626 -185
rect 1011 -238 1690 -175
rect 115 -248 1690 -238
rect -1876 -254 1690 -248
rect -10893 -280 1690 -254
rect 1799 1991 21584 2004
rect 1799 1990 14000 1991
rect 1799 1716 1919 1990
rect 4800 1989 7665 1990
rect 8848 1989 9027 1990
rect 12591 1989 12773 1990
rect 13819 1989 14000 1990
rect 14507 1989 14688 1991
rect 12591 1988 12769 1989
rect 13820 1988 14000 1989
rect 14508 1988 14688 1989
rect 15140 1988 15319 1991
rect 15478 1988 15657 1991
rect 18757 1990 20553 1991
rect 21359 1990 21584 1991
rect 13820 1987 13998 1988
rect 14508 1987 14686 1988
rect 15140 1987 15317 1988
rect 15478 1987 15655 1988
rect 20768 1857 20880 1872
rect 1799 1361 1827 1716
rect 1899 1361 1919 1716
rect 3221 1782 3399 1801
rect 3221 1712 3258 1782
rect 3370 1712 3399 1782
rect 3221 1690 3399 1712
rect 6396 1782 6574 1801
rect 6396 1712 6433 1782
rect 6545 1712 6574 1782
rect 6396 1690 6574 1712
rect 8849 1781 9027 1800
rect 8849 1711 8886 1781
rect 8998 1711 9027 1781
rect 8849 1689 9027 1711
rect 11175 1784 11353 1803
rect 11175 1714 11212 1784
rect 11324 1714 11353 1784
rect 11175 1692 11353 1714
rect 12591 1780 12769 1799
rect 20768 1798 20781 1857
rect 20865 1798 20880 1857
rect 12591 1710 12628 1780
rect 12740 1710 12769 1780
rect 12591 1688 12769 1710
rect 13820 1779 13998 1798
rect 13820 1709 13857 1779
rect 13969 1709 13998 1779
rect 13820 1687 13998 1709
rect 14508 1779 14686 1798
rect 14508 1709 14545 1779
rect 14657 1709 14686 1779
rect 14508 1687 14686 1709
rect 15140 1779 15317 1798
rect 15140 1709 15176 1779
rect 15288 1709 15317 1779
rect 15140 1688 15317 1709
rect 15478 1779 15655 1798
rect 20768 1781 20880 1798
rect 15478 1709 15514 1779
rect 15626 1709 15655 1779
rect 15478 1688 15655 1709
rect 15930 1748 16043 1763
rect 15930 1689 15943 1748
rect 16027 1689 16043 1748
rect 15930 1670 16043 1689
rect 16153 1748 16265 1763
rect 16153 1689 16166 1748
rect 16250 1689 16265 1748
rect 16153 1670 16265 1689
rect 16726 1750 16887 1767
rect 16726 1696 16752 1750
rect 16870 1696 16887 1750
rect 16726 1678 16887 1696
rect 17236 1746 17397 1763
rect 17236 1692 17262 1746
rect 17380 1692 17397 1746
rect 17236 1674 17397 1692
rect 17527 1741 17616 1771
rect 17527 1673 17542 1741
rect 17599 1673 17616 1741
rect 17527 1648 17616 1673
rect 17889 1741 17978 1771
rect 17889 1673 17904 1741
rect 17961 1673 17978 1741
rect 17889 1648 17978 1673
rect 18259 1741 18348 1771
rect 18259 1673 18274 1741
rect 18331 1673 18348 1741
rect 18259 1648 18348 1673
rect 18431 1741 18520 1771
rect 18431 1673 18446 1741
rect 18503 1673 18520 1741
rect 18431 1648 18520 1673
rect 18803 1741 18892 1771
rect 18803 1673 18818 1741
rect 18875 1673 18892 1741
rect 18803 1648 18892 1673
rect 18976 1741 19065 1771
rect 18976 1673 18991 1741
rect 19048 1673 19065 1741
rect 18976 1648 19065 1673
rect 19364 1741 19453 1771
rect 19364 1673 19379 1741
rect 19436 1673 19453 1741
rect 19364 1648 19453 1673
rect 19537 1741 19626 1770
rect 19537 1673 19552 1741
rect 19609 1673 19626 1741
rect 19537 1648 19626 1673
rect 19913 1741 20002 1770
rect 19913 1673 19928 1741
rect 19985 1673 20002 1741
rect 19913 1648 20002 1673
rect 20086 1741 20175 1770
rect 20086 1673 20101 1741
rect 20158 1673 20175 1741
rect 21427 1717 21584 1990
rect 20086 1648 20175 1673
rect 20698 1699 20771 1713
rect 1799 920 1919 1361
rect 1799 565 1824 920
rect 1896 565 1919 920
rect 1799 352 1919 565
rect 1799 -3 1820 352
rect 1892 -3 1919 352
rect 2058 1559 2121 1572
rect 2058 1550 2068 1559
rect 2114 1550 2121 1559
rect 2058 53 2067 1550
rect 2119 53 2121 1550
rect 2058 40 2068 53
rect 2114 40 2121 53
rect 2058 30 2121 40
rect 2230 1559 2293 1572
rect 2230 1550 2240 1559
rect 2286 1550 2293 1559
rect 2230 53 2239 1550
rect 2291 53 2293 1550
rect 2230 40 2240 53
rect 2286 40 2293 53
rect 2230 30 2293 40
rect 2398 1559 2461 1572
rect 2398 1550 2408 1559
rect 2454 1550 2461 1559
rect 2398 53 2407 1550
rect 2459 53 2461 1550
rect 2398 40 2408 53
rect 2454 40 2461 53
rect 2398 30 2461 40
rect 2569 1559 2632 1572
rect 2569 1550 2579 1559
rect 2625 1550 2632 1559
rect 2569 53 2578 1550
rect 2630 53 2632 1550
rect 2569 40 2579 53
rect 2625 40 2632 53
rect 2569 30 2632 40
rect 2737 1559 2800 1572
rect 2737 1550 2747 1559
rect 2793 1550 2800 1559
rect 2737 53 2746 1550
rect 2798 53 2800 1550
rect 2737 40 2747 53
rect 2793 40 2800 53
rect 2737 30 2800 40
rect 2908 1559 2971 1572
rect 2908 1550 2918 1559
rect 2964 1550 2971 1559
rect 2908 53 2917 1550
rect 2969 53 2971 1550
rect 2908 40 2918 53
rect 2964 40 2971 53
rect 2908 30 2971 40
rect 3076 1559 3139 1572
rect 3076 1550 3086 1559
rect 3132 1550 3139 1559
rect 3076 53 3085 1550
rect 3137 53 3139 1550
rect 3076 40 3086 53
rect 3132 40 3139 53
rect 3076 30 3139 40
rect 3247 1559 3310 1572
rect 3247 1550 3257 1559
rect 3303 1550 3310 1559
rect 3247 53 3256 1550
rect 3308 53 3310 1550
rect 3247 40 3257 53
rect 3303 40 3310 53
rect 3247 30 3310 40
rect 3415 1559 3478 1572
rect 3415 1550 3425 1559
rect 3471 1550 3478 1559
rect 3415 53 3424 1550
rect 3476 53 3478 1550
rect 3415 40 3425 53
rect 3471 40 3478 53
rect 3415 30 3478 40
rect 3587 1559 3650 1572
rect 3587 1550 3597 1559
rect 3643 1550 3650 1559
rect 3587 53 3596 1550
rect 3648 53 3650 1550
rect 3587 40 3597 53
rect 3643 40 3650 53
rect 3587 30 3650 40
rect 3755 1559 3818 1572
rect 3755 1550 3765 1559
rect 3811 1550 3818 1559
rect 3755 53 3764 1550
rect 3816 53 3818 1550
rect 3755 40 3765 53
rect 3811 40 3818 53
rect 3755 30 3818 40
rect 3926 1559 3989 1572
rect 3926 1550 3936 1559
rect 3982 1550 3989 1559
rect 3926 53 3935 1550
rect 3987 53 3989 1550
rect 3926 40 3936 53
rect 3982 40 3989 53
rect 3926 30 3989 40
rect 4094 1559 4157 1572
rect 4094 1550 4104 1559
rect 4150 1550 4157 1559
rect 4094 53 4103 1550
rect 4155 53 4157 1550
rect 4094 40 4104 53
rect 4150 40 4157 53
rect 4094 30 4157 40
rect 4265 1559 4328 1572
rect 4265 1550 4275 1559
rect 4321 1550 4328 1559
rect 4265 53 4274 1550
rect 4326 53 4328 1550
rect 4265 40 4275 53
rect 4321 40 4328 53
rect 4265 30 4328 40
rect 4433 1559 4496 1572
rect 4433 1550 4443 1559
rect 4489 1550 4496 1559
rect 4433 53 4442 1550
rect 4494 53 4496 1550
rect 4433 40 4443 53
rect 4489 40 4496 53
rect 4433 30 4496 40
rect 4604 1559 4667 1572
rect 4604 1550 4614 1559
rect 4660 1550 4667 1559
rect 4604 53 4613 1550
rect 4665 53 4667 1550
rect 4604 40 4614 53
rect 4660 40 4667 53
rect 4604 30 4667 40
rect 4772 1559 4835 1572
rect 4772 1550 4782 1559
rect 4828 1550 4835 1559
rect 4772 53 4781 1550
rect 4833 53 4835 1550
rect 4772 40 4782 53
rect 4828 40 4835 53
rect 4772 30 4835 40
rect 4972 1559 5035 1572
rect 4972 1550 4982 1559
rect 5028 1550 5035 1559
rect 4972 53 4981 1550
rect 5033 53 5035 1550
rect 4972 40 4982 53
rect 5028 40 5035 53
rect 4972 30 5035 40
rect 5144 1559 5207 1572
rect 5144 1550 5154 1559
rect 5200 1550 5207 1559
rect 5144 53 5153 1550
rect 5205 53 5207 1550
rect 5144 40 5154 53
rect 5200 40 5207 53
rect 5144 30 5207 40
rect 5312 1559 5375 1572
rect 5312 1550 5322 1559
rect 5368 1550 5375 1559
rect 5312 53 5321 1550
rect 5373 53 5375 1550
rect 5312 40 5322 53
rect 5368 40 5375 53
rect 5312 30 5375 40
rect 5483 1559 5546 1572
rect 5483 1550 5493 1559
rect 5539 1550 5546 1559
rect 5483 53 5492 1550
rect 5544 53 5546 1550
rect 5483 40 5493 53
rect 5539 40 5546 53
rect 5483 30 5546 40
rect 5651 1559 5714 1572
rect 5651 1550 5661 1559
rect 5707 1550 5714 1559
rect 5651 53 5660 1550
rect 5712 53 5714 1550
rect 5651 40 5661 53
rect 5707 40 5714 53
rect 5651 30 5714 40
rect 5822 1559 5885 1572
rect 5822 1550 5832 1559
rect 5878 1550 5885 1559
rect 5822 53 5831 1550
rect 5883 53 5885 1550
rect 5822 40 5832 53
rect 5878 40 5885 53
rect 5822 30 5885 40
rect 5990 1559 6053 1572
rect 5990 1550 6000 1559
rect 6046 1550 6053 1559
rect 5990 53 5999 1550
rect 6051 53 6053 1550
rect 5990 40 6000 53
rect 6046 40 6053 53
rect 5990 30 6053 40
rect 6161 1559 6224 1572
rect 6161 1550 6171 1559
rect 6217 1550 6224 1559
rect 6161 53 6170 1550
rect 6222 53 6224 1550
rect 6161 40 6171 53
rect 6217 40 6224 53
rect 6161 30 6224 40
rect 6329 1559 6392 1572
rect 6329 1550 6339 1559
rect 6385 1550 6392 1559
rect 6329 53 6338 1550
rect 6390 53 6392 1550
rect 6329 40 6339 53
rect 6385 40 6392 53
rect 6329 30 6392 40
rect 6501 1559 6564 1572
rect 6501 1550 6511 1559
rect 6557 1550 6564 1559
rect 6501 53 6510 1550
rect 6562 53 6564 1550
rect 6501 40 6511 53
rect 6557 40 6564 53
rect 6501 30 6564 40
rect 6669 1559 6732 1572
rect 6669 1550 6679 1559
rect 6725 1550 6732 1559
rect 6669 53 6678 1550
rect 6730 53 6732 1550
rect 6669 40 6679 53
rect 6725 40 6732 53
rect 6669 30 6732 40
rect 6840 1559 6903 1572
rect 6840 1550 6850 1559
rect 6896 1550 6903 1559
rect 6840 53 6849 1550
rect 6901 53 6903 1550
rect 6840 40 6850 53
rect 6896 40 6903 53
rect 6840 30 6903 40
rect 7008 1559 7071 1572
rect 7008 1550 7018 1559
rect 7064 1550 7071 1559
rect 7008 53 7017 1550
rect 7069 53 7071 1550
rect 7008 40 7018 53
rect 7064 40 7071 53
rect 7008 30 7071 40
rect 7179 1559 7242 1572
rect 7179 1550 7189 1559
rect 7235 1550 7242 1559
rect 7179 53 7188 1550
rect 7240 53 7242 1550
rect 7179 40 7189 53
rect 7235 40 7242 53
rect 7179 30 7242 40
rect 7347 1559 7410 1572
rect 7347 1550 7357 1559
rect 7403 1550 7410 1559
rect 7347 53 7356 1550
rect 7408 53 7410 1550
rect 7347 40 7357 53
rect 7403 40 7410 53
rect 7347 30 7410 40
rect 7518 1559 7581 1572
rect 7518 1550 7528 1559
rect 7574 1550 7581 1559
rect 7518 53 7527 1550
rect 7579 53 7581 1550
rect 7518 40 7528 53
rect 7574 40 7581 53
rect 7518 30 7581 40
rect 7686 1559 7749 1572
rect 7686 1550 7696 1559
rect 7742 1550 7749 1559
rect 7686 53 7695 1550
rect 7747 53 7749 1550
rect 7686 40 7696 53
rect 7742 40 7749 53
rect 7686 30 7749 40
rect 7857 1559 7920 1572
rect 7857 1550 7867 1559
rect 7913 1550 7920 1559
rect 7857 53 7866 1550
rect 7918 53 7920 1550
rect 7857 40 7867 53
rect 7913 40 7920 53
rect 7857 30 7920 40
rect 8025 1559 8088 1572
rect 8025 1550 8035 1559
rect 8081 1550 8088 1559
rect 8025 53 8034 1550
rect 8086 53 8088 1550
rect 8025 40 8035 53
rect 8081 40 8088 53
rect 8025 30 8088 40
rect 8196 1559 8259 1572
rect 8196 1550 8206 1559
rect 8252 1550 8259 1559
rect 8196 53 8205 1550
rect 8257 53 8259 1550
rect 8196 40 8206 53
rect 8252 40 8259 53
rect 8196 30 8259 40
rect 8364 1559 8427 1572
rect 8364 1550 8374 1559
rect 8420 1550 8427 1559
rect 8364 53 8373 1550
rect 8425 53 8427 1550
rect 8364 40 8374 53
rect 8420 40 8427 53
rect 8364 30 8427 40
rect 8535 1559 8598 1572
rect 8535 1550 8545 1559
rect 8591 1550 8598 1559
rect 8535 53 8544 1550
rect 8596 53 8598 1550
rect 8535 40 8545 53
rect 8591 40 8598 53
rect 8535 30 8598 40
rect 8703 1559 8766 1572
rect 8703 1550 8713 1559
rect 8759 1550 8766 1559
rect 8703 53 8712 1550
rect 8764 53 8766 1550
rect 8703 40 8713 53
rect 8759 40 8766 53
rect 8703 30 8766 40
rect 8874 1559 8937 1572
rect 8874 1550 8884 1559
rect 8930 1550 8937 1559
rect 8874 53 8883 1550
rect 8935 53 8937 1550
rect 8874 40 8884 53
rect 8930 40 8937 53
rect 8874 30 8937 40
rect 9042 1559 9105 1572
rect 9042 1550 9052 1559
rect 9098 1550 9105 1559
rect 9042 53 9051 1550
rect 9103 53 9105 1550
rect 9042 40 9052 53
rect 9098 40 9105 53
rect 9042 30 9105 40
rect 9214 1559 9277 1572
rect 9214 1550 9224 1559
rect 9270 1550 9277 1559
rect 9214 53 9223 1550
rect 9275 53 9277 1550
rect 9214 40 9224 53
rect 9270 40 9277 53
rect 9214 30 9277 40
rect 9382 1559 9445 1572
rect 9382 1550 9392 1559
rect 9438 1550 9445 1559
rect 9382 53 9391 1550
rect 9443 53 9445 1550
rect 9382 40 9392 53
rect 9438 40 9445 53
rect 9382 30 9445 40
rect 9553 1559 9616 1572
rect 9553 1550 9563 1559
rect 9609 1550 9616 1559
rect 9553 53 9562 1550
rect 9614 53 9616 1550
rect 9553 40 9563 53
rect 9609 40 9616 53
rect 9553 30 9616 40
rect 9721 1559 9784 1572
rect 9721 1550 9731 1559
rect 9777 1550 9784 1559
rect 9721 53 9730 1550
rect 9782 53 9784 1550
rect 9721 40 9731 53
rect 9777 40 9784 53
rect 9721 30 9784 40
rect 9892 1559 9955 1572
rect 9892 1550 9902 1559
rect 9948 1550 9955 1559
rect 9892 53 9901 1550
rect 9953 53 9955 1550
rect 9892 40 9902 53
rect 9948 40 9955 53
rect 9892 30 9955 40
rect 10060 1559 10123 1572
rect 10060 1550 10070 1559
rect 10116 1550 10123 1559
rect 10060 53 10069 1550
rect 10121 53 10123 1550
rect 10060 40 10070 53
rect 10116 40 10123 53
rect 10060 30 10123 40
rect 10231 1559 10294 1572
rect 10231 1550 10241 1559
rect 10287 1550 10294 1559
rect 10231 53 10240 1550
rect 10292 53 10294 1550
rect 10231 40 10241 53
rect 10287 40 10294 53
rect 10231 30 10294 40
rect 10399 1559 10462 1572
rect 10399 1550 10409 1559
rect 10455 1550 10462 1559
rect 10399 53 10408 1550
rect 10460 53 10462 1550
rect 10399 40 10409 53
rect 10455 40 10462 53
rect 10399 30 10462 40
rect 10587 1559 10650 1572
rect 10587 1550 10597 1559
rect 10643 1550 10650 1559
rect 10587 53 10596 1550
rect 10648 53 10650 1550
rect 10587 40 10597 53
rect 10643 40 10650 53
rect 10587 30 10650 40
rect 10758 1559 10821 1572
rect 10758 1550 10768 1559
rect 10814 1550 10821 1559
rect 10758 53 10767 1550
rect 10819 53 10821 1550
rect 10758 40 10768 53
rect 10814 40 10821 53
rect 10758 30 10821 40
rect 10926 1559 10989 1572
rect 10926 1550 10936 1559
rect 10982 1550 10989 1559
rect 10926 53 10935 1550
rect 10987 53 10989 1550
rect 10926 40 10936 53
rect 10982 40 10989 53
rect 10926 30 10989 40
rect 11097 1559 11160 1572
rect 11097 1550 11107 1559
rect 11153 1550 11160 1559
rect 11097 53 11106 1550
rect 11158 53 11160 1550
rect 11097 40 11107 53
rect 11153 40 11160 53
rect 11097 30 11160 40
rect 11265 1559 11328 1572
rect 11265 1550 11275 1559
rect 11321 1550 11328 1559
rect 11265 53 11274 1550
rect 11326 53 11328 1550
rect 11265 40 11275 53
rect 11321 40 11328 53
rect 11265 30 11328 40
rect 11436 1559 11499 1572
rect 11436 1550 11446 1559
rect 11492 1550 11499 1559
rect 11436 53 11445 1550
rect 11497 53 11499 1550
rect 11436 40 11446 53
rect 11492 40 11499 53
rect 11436 30 11499 40
rect 11604 1559 11667 1572
rect 11604 1550 11614 1559
rect 11660 1550 11667 1559
rect 11604 53 11613 1550
rect 11665 53 11667 1550
rect 11604 40 11614 53
rect 11660 40 11667 53
rect 11604 30 11667 40
rect 11775 1559 11838 1572
rect 11775 1550 11785 1559
rect 11831 1550 11838 1559
rect 11775 53 11784 1550
rect 11836 53 11838 1550
rect 11775 40 11785 53
rect 11831 40 11838 53
rect 11775 30 11838 40
rect 11943 1559 12006 1572
rect 11943 1550 11953 1559
rect 11999 1550 12006 1559
rect 11943 53 11952 1550
rect 12004 53 12006 1550
rect 11943 40 11953 53
rect 11999 40 12006 53
rect 11943 30 12006 40
rect 12115 1559 12178 1572
rect 12115 1550 12125 1559
rect 12171 1550 12178 1559
rect 12115 53 12124 1550
rect 12176 53 12178 1550
rect 12115 40 12125 53
rect 12171 40 12178 53
rect 12115 30 12178 40
rect 12283 1559 12346 1572
rect 12283 1550 12293 1559
rect 12339 1550 12346 1559
rect 12283 53 12292 1550
rect 12344 53 12346 1550
rect 12283 40 12293 53
rect 12339 40 12346 53
rect 12283 30 12346 40
rect 12454 1559 12517 1572
rect 12454 1550 12464 1559
rect 12510 1550 12517 1559
rect 12454 53 12463 1550
rect 12515 53 12517 1550
rect 12454 40 12464 53
rect 12510 40 12517 53
rect 12454 30 12517 40
rect 12622 1559 12685 1572
rect 12622 1550 12632 1559
rect 12678 1550 12685 1559
rect 12622 53 12631 1550
rect 12683 53 12685 1550
rect 12622 40 12632 53
rect 12678 40 12685 53
rect 12622 30 12685 40
rect 12793 1559 12856 1572
rect 12793 1550 12803 1559
rect 12849 1550 12856 1559
rect 12793 53 12802 1550
rect 12854 53 12856 1550
rect 12793 40 12803 53
rect 12849 40 12856 53
rect 12793 30 12856 40
rect 12961 1559 13024 1572
rect 12961 1550 12971 1559
rect 13017 1550 13024 1559
rect 12961 53 12970 1550
rect 13022 53 13024 1550
rect 12961 40 12971 53
rect 13017 40 13024 53
rect 12961 30 13024 40
rect 13132 1559 13195 1572
rect 13132 1550 13142 1559
rect 13188 1550 13195 1559
rect 13132 53 13141 1550
rect 13193 53 13195 1550
rect 13132 40 13142 53
rect 13188 40 13195 53
rect 13132 30 13195 40
rect 13300 1559 13363 1572
rect 13300 1550 13310 1559
rect 13356 1550 13363 1559
rect 13300 53 13309 1550
rect 13361 53 13363 1550
rect 13300 40 13310 53
rect 13356 40 13363 53
rect 13300 30 13363 40
rect 13486 1559 13549 1572
rect 13486 1550 13496 1559
rect 13542 1550 13549 1559
rect 13486 53 13495 1550
rect 13547 53 13549 1550
rect 13486 40 13496 53
rect 13542 40 13549 53
rect 13486 30 13549 40
rect 13658 1559 13721 1572
rect 13658 1550 13668 1559
rect 13714 1550 13721 1559
rect 13658 53 13667 1550
rect 13719 53 13721 1550
rect 13658 40 13668 53
rect 13714 40 13721 53
rect 13658 30 13721 40
rect 13826 1559 13889 1572
rect 13826 1550 13836 1559
rect 13882 1550 13889 1559
rect 13826 53 13835 1550
rect 13887 53 13889 1550
rect 13826 40 13836 53
rect 13882 40 13889 53
rect 13826 30 13889 40
rect 13997 1559 14060 1572
rect 13997 1550 14007 1559
rect 14053 1550 14060 1559
rect 13997 53 14006 1550
rect 14058 53 14060 1550
rect 13997 40 14007 53
rect 14053 40 14060 53
rect 13997 30 14060 40
rect 14165 1559 14228 1572
rect 14165 1550 14175 1559
rect 14221 1550 14228 1559
rect 14165 53 14174 1550
rect 14226 53 14228 1550
rect 14165 40 14175 53
rect 14221 40 14228 53
rect 14165 30 14228 40
rect 14336 1559 14399 1572
rect 14336 1550 14346 1559
rect 14392 1550 14399 1559
rect 14336 53 14345 1550
rect 14397 53 14399 1550
rect 14336 40 14346 53
rect 14392 40 14399 53
rect 14336 30 14399 40
rect 14504 1559 14567 1572
rect 14504 1550 14514 1559
rect 14560 1550 14567 1559
rect 14504 53 14513 1550
rect 14565 53 14567 1550
rect 14504 40 14514 53
rect 14560 40 14567 53
rect 14504 30 14567 40
rect 14675 1559 14738 1572
rect 14675 1550 14685 1559
rect 14731 1550 14738 1559
rect 14675 53 14684 1550
rect 14736 53 14738 1550
rect 14675 40 14685 53
rect 14731 40 14738 53
rect 14675 30 14738 40
rect 14843 1559 14906 1572
rect 14843 1550 14853 1559
rect 14899 1550 14906 1559
rect 14843 53 14852 1550
rect 14904 53 14906 1550
rect 14843 40 14853 53
rect 14899 40 14906 53
rect 14843 30 14906 40
rect 15027 1559 15090 1572
rect 15027 1550 15037 1559
rect 15083 1550 15090 1559
rect 15027 53 15036 1550
rect 15088 53 15090 1550
rect 15027 40 15037 53
rect 15083 40 15090 53
rect 15027 30 15090 40
rect 15198 1559 15261 1572
rect 15198 1550 15208 1559
rect 15254 1550 15261 1559
rect 15198 53 15207 1550
rect 15259 53 15261 1550
rect 15198 40 15208 53
rect 15254 40 15261 53
rect 15198 30 15261 40
rect 15366 1559 15429 1572
rect 15366 1550 15376 1559
rect 15422 1550 15429 1559
rect 15366 53 15375 1550
rect 15427 53 15429 1550
rect 15366 40 15376 53
rect 15422 40 15429 53
rect 15366 30 15429 40
rect 15537 1559 15600 1572
rect 15537 1550 15547 1559
rect 15593 1550 15600 1559
rect 15537 53 15546 1550
rect 15598 53 15600 1550
rect 15537 40 15547 53
rect 15593 40 15600 53
rect 15537 30 15600 40
rect 15705 1559 15768 1572
rect 15705 1550 15715 1559
rect 15761 1550 15768 1559
rect 15705 53 15714 1550
rect 15766 53 15768 1550
rect 15705 40 15715 53
rect 15761 40 15768 53
rect 15705 30 15768 40
rect 15897 1559 15960 1572
rect 15897 1550 15907 1559
rect 15953 1550 15960 1559
rect 15897 53 15906 1550
rect 15958 53 15960 1550
rect 15897 40 15907 53
rect 15953 40 15960 53
rect 15897 30 15960 40
rect 16068 1559 16131 1572
rect 16068 1550 16078 1559
rect 16124 1550 16131 1559
rect 16068 53 16077 1550
rect 16129 53 16131 1550
rect 16068 40 16078 53
rect 16124 40 16131 53
rect 16068 30 16131 40
rect 16236 1559 16299 1572
rect 16236 1550 16246 1559
rect 16292 1550 16299 1559
rect 16236 53 16245 1550
rect 16297 53 16299 1550
rect 16236 40 16246 53
rect 16292 40 16299 53
rect 16236 30 16299 40
rect 16437 1559 16500 1572
rect 16437 1545 16447 1559
rect 16493 1545 16500 1559
rect 16437 53 16446 1545
rect 16498 53 16500 1545
rect 16437 40 16447 53
rect 16493 40 16500 53
rect 16437 30 16500 40
rect 16608 1559 16671 1572
rect 16608 1545 16618 1559
rect 16664 1545 16671 1559
rect 16608 53 16617 1545
rect 16669 53 16671 1545
rect 16608 40 16618 53
rect 16664 40 16671 53
rect 16608 30 16671 40
rect 16776 1559 16839 1572
rect 16776 1545 16786 1559
rect 16832 1545 16839 1559
rect 16776 53 16785 1545
rect 16837 53 16839 1545
rect 16776 40 16786 53
rect 16832 40 16839 53
rect 16776 30 16839 40
rect 16947 1559 17010 1572
rect 16947 1545 16957 1559
rect 17003 1545 17010 1559
rect 16947 53 16956 1545
rect 17008 53 17010 1545
rect 16947 40 16957 53
rect 17003 40 17010 53
rect 16947 30 17010 40
rect 17115 1559 17178 1572
rect 17115 1545 17125 1559
rect 17171 1545 17178 1559
rect 17115 53 17124 1545
rect 17176 53 17178 1545
rect 17115 40 17125 53
rect 17171 40 17178 53
rect 17115 30 17178 40
rect 17286 1559 17349 1572
rect 17286 1545 17296 1559
rect 17342 1545 17349 1559
rect 17286 53 17295 1545
rect 17347 53 17349 1545
rect 17286 40 17296 53
rect 17342 40 17349 53
rect 17286 30 17349 40
rect 17454 1559 17517 1572
rect 17454 1545 17464 1559
rect 17510 1545 17517 1559
rect 17454 53 17463 1545
rect 17515 53 17517 1545
rect 17454 40 17464 53
rect 17510 40 17517 53
rect 17454 30 17517 40
rect 17625 1559 17688 1572
rect 17625 1545 17635 1559
rect 17681 1545 17688 1559
rect 17625 53 17634 1545
rect 17686 53 17688 1545
rect 17816 1559 17879 1572
rect 17816 1545 17826 1559
rect 17872 1545 17879 1559
rect 17816 830 17825 1545
rect 17877 830 17879 1545
rect 17816 814 17879 830
rect 17987 1559 18050 1572
rect 17987 1545 17997 1559
rect 18043 1545 18050 1559
rect 17987 830 17996 1545
rect 18048 830 18050 1545
rect 18198 1559 18261 1572
rect 18198 1545 18208 1559
rect 18254 1545 18261 1559
rect 18198 1241 18207 1545
rect 18259 1241 18261 1545
rect 18198 1220 18261 1241
rect 18369 1559 18432 1572
rect 18369 1545 18379 1559
rect 18425 1545 18432 1559
rect 18369 1240 18378 1545
rect 18430 1240 18432 1545
rect 18369 1220 18432 1240
rect 18540 1559 18603 1572
rect 18540 1545 18550 1559
rect 18596 1545 18603 1559
rect 18540 1240 18549 1545
rect 18601 1240 18603 1545
rect 18540 1220 18603 1240
rect 18748 1559 18811 1572
rect 18748 1545 18758 1559
rect 18804 1545 18811 1559
rect 18748 1240 18757 1545
rect 18809 1240 18811 1545
rect 18748 1220 18811 1240
rect 18917 1559 18980 1572
rect 18917 1545 18927 1559
rect 18973 1545 18980 1559
rect 18917 1240 18926 1545
rect 18978 1240 18980 1545
rect 18917 1220 18980 1240
rect 19088 1559 19151 1572
rect 19088 1545 19098 1559
rect 19144 1545 19151 1559
rect 19088 1240 19097 1545
rect 19149 1240 19151 1545
rect 19088 1220 19151 1240
rect 19309 1559 19372 1572
rect 19309 1545 19319 1559
rect 19365 1545 19372 1559
rect 19309 1240 19318 1545
rect 19370 1240 19372 1545
rect 19309 1220 19372 1240
rect 19478 1559 19541 1572
rect 19478 1545 19488 1559
rect 19534 1545 19541 1559
rect 19478 1240 19487 1545
rect 19539 1240 19541 1545
rect 19478 1220 19541 1240
rect 19649 1559 19712 1572
rect 19649 1545 19659 1559
rect 19705 1545 19712 1559
rect 19649 1240 19658 1545
rect 19710 1240 19712 1545
rect 19649 1220 19712 1240
rect 19858 1559 19921 1572
rect 19858 1545 19868 1559
rect 19914 1545 19921 1559
rect 19858 1240 19867 1545
rect 19919 1240 19921 1545
rect 19858 1220 19921 1240
rect 20027 1559 20090 1572
rect 20027 1545 20037 1559
rect 20083 1545 20090 1559
rect 20027 1240 20036 1545
rect 20088 1240 20090 1545
rect 20027 1220 20090 1240
rect 20198 1559 20261 1572
rect 20198 1545 20208 1559
rect 20254 1545 20261 1559
rect 20198 1240 20207 1545
rect 20259 1240 20261 1545
rect 20198 1220 20261 1240
rect 20698 1160 20708 1699
rect 20759 1654 20771 1699
rect 20760 1188 20771 1654
rect 20759 1160 20771 1188
rect 20698 1139 20771 1160
rect 20863 1699 20936 1717
rect 20863 1160 20875 1699
rect 20926 1655 20936 1699
rect 20927 1189 20936 1655
rect 20926 1160 20936 1189
rect 20863 1143 20936 1160
rect 21427 1156 21469 1717
rect 21563 1156 21584 1717
rect 18343 943 18466 974
rect 18534 970 18640 971
rect 18343 874 18377 943
rect 18440 874 18466 943
rect 18343 840 18466 874
rect 18533 936 18640 970
rect 18533 867 18552 936
rect 18615 867 18640 936
rect 18533 838 18640 867
rect 18534 835 18640 838
rect 18883 935 18968 969
rect 18883 866 18893 935
rect 18956 866 18968 935
rect 18883 837 18968 866
rect 19039 936 19133 970
rect 19039 867 19058 936
rect 19121 867 19133 936
rect 19039 838 19133 867
rect 19402 935 19487 969
rect 19402 866 19412 935
rect 19475 866 19487 935
rect 19402 837 19487 866
rect 19558 936 19652 970
rect 19558 867 19577 936
rect 19640 867 19652 936
rect 19558 838 19652 867
rect 19922 935 20007 969
rect 19922 866 19932 935
rect 19995 866 20007 935
rect 19922 837 20007 866
rect 20078 936 20172 970
rect 20078 867 20097 936
rect 20160 867 20172 936
rect 20078 838 20172 867
rect 20454 935 20539 969
rect 20454 866 20464 935
rect 20527 866 20539 935
rect 20454 837 20539 866
rect 20610 936 20704 970
rect 20610 867 20629 936
rect 20692 867 20704 936
rect 20610 838 20704 867
rect 20972 935 21057 969
rect 20972 866 20982 935
rect 21045 866 21057 935
rect 20972 837 21057 866
rect 21128 936 21222 970
rect 21128 867 21147 936
rect 21210 867 21222 936
rect 21128 838 21222 867
rect 17987 814 18050 830
rect 17625 40 17635 53
rect 17681 40 17688 53
rect 17625 30 17688 40
rect 18285 748 18348 761
rect 18285 734 18295 748
rect 18341 734 18348 748
rect 18285 19 18294 734
rect 18346 19 18348 734
rect 18285 3 18348 19
rect 18456 748 18519 761
rect 18456 734 18466 748
rect 18512 734 18519 748
rect 18456 19 18465 734
rect 18517 19 18519 734
rect 18456 3 18519 19
rect 18627 748 18690 761
rect 18627 734 18637 748
rect 18683 734 18690 748
rect 18627 19 18636 734
rect 18688 19 18690 734
rect 18627 3 18690 19
rect 18799 748 18862 761
rect 18799 734 18809 748
rect 18855 734 18862 748
rect 18799 19 18808 734
rect 18860 19 18862 734
rect 18799 3 18862 19
rect 18968 748 19031 761
rect 18968 734 18978 748
rect 19024 734 19031 748
rect 18968 19 18977 734
rect 19029 19 19031 734
rect 18968 3 19031 19
rect 19139 748 19202 761
rect 19139 734 19149 748
rect 19195 734 19202 748
rect 19139 19 19148 734
rect 19200 19 19202 734
rect 19318 748 19381 761
rect 19318 734 19328 748
rect 19374 734 19381 748
rect 19318 718 19327 734
rect 19317 624 19326 718
rect 19139 3 19202 19
rect 19318 19 19327 624
rect 19379 19 19381 734
rect 19318 3 19381 19
rect 19487 748 19550 761
rect 19487 734 19497 748
rect 19543 734 19550 748
rect 19487 19 19496 734
rect 19548 19 19550 734
rect 19658 748 19721 761
rect 19658 734 19668 748
rect 19714 734 19721 748
rect 19658 530 19667 734
rect 19656 430 19665 530
rect 19487 3 19550 19
rect 19658 19 19667 430
rect 19719 19 19721 734
rect 19838 748 19901 761
rect 19838 734 19848 748
rect 19894 734 19901 748
rect 19838 717 19847 734
rect 19837 623 19846 717
rect 19658 3 19721 19
rect 19838 19 19847 623
rect 19899 19 19901 734
rect 19838 3 19901 19
rect 20007 748 20070 761
rect 20007 734 20017 748
rect 20063 734 20070 748
rect 20007 19 20016 734
rect 20068 19 20070 734
rect 20178 748 20241 761
rect 20178 734 20188 748
rect 20234 734 20241 748
rect 20178 530 20187 734
rect 20175 430 20184 530
rect 20007 3 20070 19
rect 20178 19 20187 430
rect 20239 19 20241 734
rect 20370 748 20433 761
rect 20370 734 20380 748
rect 20426 734 20433 748
rect 20370 729 20379 734
rect 20365 635 20374 729
rect 20178 3 20241 19
rect 20370 19 20379 635
rect 20431 19 20433 734
rect 20370 3 20433 19
rect 20539 748 20602 761
rect 20539 734 20549 748
rect 20595 734 20602 748
rect 20539 19 20548 734
rect 20600 19 20602 734
rect 20710 748 20773 761
rect 20710 734 20720 748
rect 20766 734 20773 748
rect 20710 530 20719 734
rect 20706 430 20715 530
rect 20539 3 20602 19
rect 20710 19 20719 430
rect 20771 19 20773 734
rect 20888 748 20951 761
rect 20888 734 20898 748
rect 20944 734 20951 748
rect 20888 724 20897 734
rect 20884 630 20893 724
rect 20710 3 20773 19
rect 20888 19 20897 630
rect 20949 19 20951 734
rect 20888 3 20951 19
rect 21057 748 21120 761
rect 21057 734 21067 748
rect 21113 734 21120 748
rect 21057 19 21066 734
rect 21118 19 21120 734
rect 21228 748 21291 761
rect 21228 734 21238 748
rect 21284 734 21291 748
rect 21228 530 21237 734
rect 21223 430 21232 530
rect 21057 3 21120 19
rect 21228 19 21237 430
rect 21289 19 21291 734
rect 21228 3 21291 19
rect 21427 538 21584 1156
rect 1799 -148 1919 -3
rect 21427 -23 21462 538
rect 21556 -23 21584 538
rect 1799 -149 17252 -148
rect 18821 -149 20526 -147
rect 21427 -149 21584 -23
rect 1799 -161 21584 -149
rect 1799 -165 7595 -161
rect 1799 -168 3667 -165
rect 1799 -262 2224 -168
rect 2785 -259 3667 -168
rect 4228 -172 6375 -165
rect 4228 -259 5075 -172
rect 2785 -262 5075 -259
rect 1799 -266 5075 -262
rect 5636 -259 6375 -172
rect 6936 -255 7595 -165
rect 8156 -162 21584 -161
rect 8156 -165 18628 -162
rect 8156 -168 13452 -165
rect 8156 -255 9024 -168
rect 6936 -259 9024 -255
rect 5636 -262 9024 -259
rect 9585 -262 10334 -168
rect 10895 -262 11982 -168
rect 12543 -259 13452 -168
rect 14013 -259 15071 -165
rect 15632 -169 18628 -165
rect 15632 -259 16873 -169
rect 12543 -262 16873 -259
rect 5636 -263 16873 -262
rect 17434 -256 18628 -169
rect 19189 -165 21584 -162
rect 19189 -256 20208 -165
rect 17434 -259 20208 -256
rect 20769 -259 21584 -165
rect 17434 -263 21584 -259
rect 5636 -266 21584 -263
rect 1799 -279 21584 -266
rect 1799 -280 1919 -279
rect -10893 -281 1687 -280
rect 4844 -281 21584 -279
rect 17245 -282 21435 -281
<< via1 >>
rect -10645 2024 -10260 2087
rect -9736 2021 -9351 2084
rect -8322 2019 -7937 2082
rect -7244 2020 -6859 2083
rect -6214 2026 -5829 2089
rect -5186 2016 -4801 2079
rect -4309 2031 -3924 2094
rect -3355 2029 -2970 2092
rect -2495 2028 -2110 2091
rect -1528 2024 -1143 2087
rect -162 2026 223 2089
rect 876 2026 1261 2089
rect 2184 2007 2745 2101
rect 3780 2012 4341 2106
rect 5230 2005 5791 2099
rect 6883 2013 7444 2107
rect 8198 2010 8759 2104
rect 9727 2013 10288 2107
rect 11480 2008 12041 2102
rect 12864 2004 13425 2098
rect 14532 2006 15093 2100
rect 16308 2012 16869 2106
rect 17623 2016 18184 2110
rect 19309 2013 19870 2107
rect 20507 2006 21068 2100
rect -10868 1461 -10805 1846
rect -7618 1703 -7557 1767
rect -3629 1706 -3568 1770
rect -1901 1704 -1840 1768
rect -945 1700 -884 1764
rect -451 1693 -390 1757
rect -22 1678 39 1742
rect 191 1678 252 1742
rect 529 1679 590 1743
rect 744 1678 805 1742
rect 1099 1676 1160 1740
rect 1312 1678 1373 1742
rect -10860 864 -10797 1249
rect -10855 66 -10792 451
rect -10561 50 -10560 1549
rect -10560 50 -10514 1549
rect -10514 50 -10509 1549
rect -10394 48 -10348 1549
rect -10348 48 -10341 1549
rect -10230 50 -10229 1549
rect -10229 50 -10183 1549
rect -10183 50 -10178 1549
rect -10063 236 -10017 1549
rect -10017 236 -10010 1549
rect -10063 125 -10015 236
rect -10015 125 -10008 236
rect -10063 48 -10017 125
rect -10017 48 -10010 125
rect -9899 50 -9898 1549
rect -9898 50 -9852 1549
rect -9852 50 -9847 1549
rect -9732 235 -9686 1549
rect -9734 124 -9686 235
rect -9732 48 -9686 124
rect -9686 48 -9679 1549
rect -9568 50 -9567 1549
rect -9567 50 -9521 1549
rect -9521 50 -9516 1549
rect -9401 234 -9355 1549
rect -9403 123 -9355 234
rect -9401 48 -9355 123
rect -9355 48 -9348 1549
rect -9235 50 -9234 1549
rect -9234 50 -9188 1549
rect -9188 50 -9183 1549
rect -9068 237 -9022 1549
rect -9070 126 -9022 237
rect -9068 48 -9022 126
rect -9022 48 -9015 1549
rect -8904 50 -8903 1549
rect -8903 50 -8857 1549
rect -8857 50 -8852 1549
rect -8737 237 -8691 1549
rect -8739 126 -8691 237
rect -8737 48 -8691 126
rect -8691 48 -8684 1549
rect -8573 50 -8572 1549
rect -8572 50 -8526 1549
rect -8526 50 -8521 1549
rect -8406 239 -8360 1549
rect -8408 128 -8360 239
rect -8406 48 -8360 128
rect -8360 48 -8353 1549
rect -8242 50 -8241 1549
rect -8241 50 -8195 1549
rect -8195 50 -8190 1549
rect -8075 241 -8029 1549
rect -8029 241 -8022 1549
rect -8076 130 -8028 241
rect -8028 130 -8021 241
rect -8075 48 -8029 130
rect -8029 48 -8022 130
rect -7910 50 -7909 1549
rect -7909 50 -7863 1549
rect -7863 50 -7858 1549
rect -7743 241 -7697 1549
rect -7745 130 -7697 241
rect -7743 48 -7697 130
rect -7697 48 -7690 1549
rect -7579 50 -7578 1549
rect -7578 50 -7532 1549
rect -7532 50 -7527 1549
rect -7412 241 -7366 1549
rect -7366 241 -7359 1549
rect -7413 130 -7365 241
rect -7365 130 -7358 241
rect -7412 48 -7366 130
rect -7366 48 -7359 130
rect -7248 50 -7247 1549
rect -7247 50 -7201 1549
rect -7201 50 -7196 1549
rect -7081 241 -7035 1549
rect -7035 241 -7028 1549
rect -7082 130 -7034 241
rect -7034 130 -7027 241
rect -7081 48 -7035 130
rect -7035 48 -7028 130
rect -6917 50 -6916 1549
rect -6916 50 -6870 1549
rect -6870 50 -6865 1549
rect -6750 241 -6704 1549
rect -6752 130 -6704 241
rect -6750 48 -6704 130
rect -6704 48 -6697 1549
rect -6584 50 -6583 1549
rect -6583 50 -6537 1549
rect -6537 50 -6532 1549
rect -6417 241 -6371 1549
rect -6419 130 -6371 241
rect -6417 48 -6371 130
rect -6371 48 -6364 1549
rect -6253 50 -6252 1549
rect -6252 50 -6206 1549
rect -6206 50 -6201 1549
rect -6086 241 -6040 1549
rect -6088 130 -6040 241
rect -6086 48 -6040 130
rect -6040 48 -6033 1549
rect -5922 50 -5921 1549
rect -5921 50 -5875 1549
rect -5875 50 -5870 1549
rect -5755 251 -5709 1549
rect -5709 251 -5702 1549
rect -5755 140 -5707 251
rect -5707 140 -5700 251
rect -5755 48 -5709 140
rect -5709 48 -5702 140
rect -5591 50 -5590 1549
rect -5590 50 -5544 1549
rect -5544 50 -5539 1549
rect -5424 251 -5378 1549
rect -5426 140 -5378 251
rect -5424 48 -5378 140
rect -5378 48 -5371 1549
rect -5258 50 -5257 1549
rect -5257 50 -5211 1549
rect -5211 50 -5206 1549
rect -5091 48 -5045 1549
rect -5045 48 -5038 1549
rect -4927 50 -4926 1549
rect -4926 50 -4880 1549
rect -4880 50 -4875 1549
rect -4760 252 -4714 1549
rect -4714 252 -4707 1549
rect -4760 150 -4712 252
rect -4712 150 -4705 252
rect -4760 48 -4714 150
rect -4714 48 -4707 150
rect -4596 50 -4595 1549
rect -4595 50 -4549 1549
rect -4549 50 -4544 1549
rect -4429 252 -4383 1549
rect -4383 252 -4376 1549
rect -4430 150 -4382 252
rect -4382 150 -4375 252
rect -4429 48 -4383 150
rect -4383 48 -4376 150
rect -4265 50 -4264 1549
rect -4264 50 -4218 1549
rect -4218 50 -4213 1549
rect -4098 252 -4052 1549
rect -4100 150 -4052 252
rect -4098 48 -4052 150
rect -4052 48 -4045 1549
rect -3932 50 -3931 1549
rect -3931 50 -3885 1549
rect -3885 50 -3880 1549
rect -3765 252 -3719 1549
rect -3719 252 -3712 1549
rect -3766 150 -3718 252
rect -3718 150 -3711 252
rect -3765 48 -3719 150
rect -3719 48 -3712 150
rect -3601 50 -3600 1549
rect -3600 50 -3554 1549
rect -3554 50 -3549 1549
rect -3434 252 -3388 1549
rect -3388 252 -3381 1549
rect -3435 150 -3387 252
rect -3387 150 -3380 252
rect -3434 48 -3388 150
rect -3388 48 -3381 150
rect -3270 50 -3269 1549
rect -3269 50 -3223 1549
rect -3223 50 -3218 1549
rect -3103 251 -3057 1549
rect -3105 149 -3057 251
rect -3103 48 -3057 149
rect -3057 48 -3050 1549
rect -2939 50 -2938 1549
rect -2938 50 -2892 1549
rect -2892 50 -2887 1549
rect -2772 252 -2726 1549
rect -2774 150 -2726 252
rect -2772 48 -2726 150
rect -2726 48 -2719 1549
rect -2609 50 -2608 1549
rect -2608 50 -2562 1549
rect -2562 50 -2557 1549
rect -2442 252 -2396 1549
rect -2396 252 -2389 1549
rect -2443 150 -2395 252
rect -2395 150 -2388 252
rect -2442 48 -2396 150
rect -2396 48 -2389 150
rect -2278 50 -2277 1549
rect -2277 50 -2231 1549
rect -2231 50 -2226 1549
rect -2111 252 -2065 1549
rect -2065 252 -2058 1549
rect -2112 150 -2064 252
rect -2064 150 -2057 252
rect -2111 48 -2065 150
rect -2065 48 -2058 150
rect -1947 50 -1946 1549
rect -1946 50 -1900 1549
rect -1900 50 -1895 1549
rect -1780 252 -1734 1549
rect -1782 150 -1734 252
rect -1780 48 -1734 150
rect -1734 48 -1727 1549
rect -1616 50 -1615 1549
rect -1615 50 -1569 1549
rect -1569 50 -1564 1549
rect -1449 252 -1403 1549
rect -1403 252 -1396 1549
rect -1450 150 -1402 252
rect -1402 150 -1395 252
rect -1449 48 -1403 150
rect -1403 48 -1396 150
rect -1284 50 -1283 1549
rect -1283 50 -1237 1549
rect -1237 50 -1232 1549
rect -1117 252 -1071 1549
rect -1119 150 -1071 252
rect -1117 48 -1071 150
rect -1071 48 -1064 1549
rect -953 50 -952 1549
rect -952 50 -906 1549
rect -906 50 -901 1549
rect -786 252 -740 1549
rect -740 252 -733 1549
rect -787 150 -739 252
rect -739 150 -732 252
rect -786 48 -740 150
rect -740 48 -733 150
rect -622 50 -621 1549
rect -621 50 -575 1549
rect -575 50 -570 1549
rect -455 252 -409 1549
rect -409 252 -402 1549
rect -456 150 -408 252
rect -408 150 -401 252
rect -455 48 -409 150
rect -409 48 -402 150
rect -289 48 -243 1549
rect -243 48 -236 1549
rect -80 252 -79 1549
rect -79 252 -33 1549
rect -85 150 -33 252
rect -80 50 -79 150
rect -79 50 -33 150
rect -33 50 -28 1549
rect 87 48 133 1549
rect 133 48 140 1549
rect 253 252 299 1549
rect 299 252 306 1549
rect 473 252 474 1549
rect 474 252 520 1549
rect 251 150 303 252
rect 303 150 308 252
rect 467 150 520 252
rect 253 48 299 150
rect 299 48 306 150
rect 473 50 474 150
rect 474 50 520 150
rect 520 50 525 1549
rect 640 48 686 1549
rect 686 48 693 1549
rect 806 48 852 1549
rect 852 48 859 1549
rect 1042 255 1043 1549
rect 1043 255 1089 1549
rect 1041 150 1089 255
rect 1042 50 1043 150
rect 1043 50 1089 150
rect 1089 50 1094 1549
rect 1209 48 1255 1549
rect 1255 48 1262 1549
rect 1375 255 1421 1549
rect 1421 255 1428 1549
rect 1375 150 1423 255
rect 1423 150 1428 255
rect 1375 48 1421 150
rect 1421 48 1428 150
rect 1600 1355 1663 1740
rect 1599 586 1662 971
rect 1598 -6 1661 379
rect -10444 -245 -10059 -182
rect -9441 -246 -9056 -183
rect -8567 -238 -8182 -175
rect -7658 -244 -7273 -181
rect -6670 -249 -6285 -186
rect -5464 -247 -5079 -184
rect -4325 -242 -3940 -179
rect -3208 -248 -2823 -185
rect -2261 -254 -1876 -191
rect -1140 -248 -755 -185
rect -270 -248 115 -185
rect 626 -238 1011 -175
rect 1827 1361 1899 1716
rect 3258 1712 3370 1782
rect 6433 1712 6545 1782
rect 8886 1711 8998 1781
rect 11212 1714 11324 1784
rect 20781 1798 20865 1857
rect 12628 1710 12740 1780
rect 13857 1709 13969 1779
rect 14545 1709 14657 1779
rect 15176 1709 15288 1779
rect 15514 1709 15626 1779
rect 15943 1689 16027 1748
rect 16166 1689 16250 1748
rect 16752 1696 16870 1750
rect 17262 1692 17380 1746
rect 17542 1673 17599 1741
rect 17904 1673 17961 1741
rect 18274 1673 18331 1741
rect 18446 1673 18503 1741
rect 18818 1673 18875 1741
rect 18991 1673 19048 1741
rect 19379 1673 19436 1741
rect 19552 1673 19609 1741
rect 19928 1673 19985 1741
rect 20101 1673 20158 1741
rect 1824 565 1896 920
rect 1820 -3 1892 352
rect 2067 53 2068 1550
rect 2068 53 2114 1550
rect 2114 53 2119 1550
rect 2239 53 2240 1550
rect 2240 53 2286 1550
rect 2286 53 2291 1550
rect 2407 53 2408 1550
rect 2408 53 2454 1550
rect 2454 53 2459 1550
rect 2578 53 2579 1550
rect 2579 53 2625 1550
rect 2625 53 2630 1550
rect 2746 53 2747 1550
rect 2747 53 2793 1550
rect 2793 53 2798 1550
rect 2917 53 2918 1550
rect 2918 53 2964 1550
rect 2964 53 2969 1550
rect 3085 53 3086 1550
rect 3086 53 3132 1550
rect 3132 53 3137 1550
rect 3256 53 3257 1550
rect 3257 53 3303 1550
rect 3303 53 3308 1550
rect 3424 53 3425 1550
rect 3425 53 3471 1550
rect 3471 53 3476 1550
rect 3596 53 3597 1550
rect 3597 53 3643 1550
rect 3643 53 3648 1550
rect 3764 53 3765 1550
rect 3765 53 3811 1550
rect 3811 53 3816 1550
rect 3935 53 3936 1550
rect 3936 53 3982 1550
rect 3982 53 3987 1550
rect 4103 53 4104 1550
rect 4104 53 4150 1550
rect 4150 53 4155 1550
rect 4274 53 4275 1550
rect 4275 53 4321 1550
rect 4321 53 4326 1550
rect 4442 53 4443 1550
rect 4443 53 4489 1550
rect 4489 53 4494 1550
rect 4613 53 4614 1550
rect 4614 53 4660 1550
rect 4660 53 4665 1550
rect 4781 53 4782 1550
rect 4782 53 4828 1550
rect 4828 53 4833 1550
rect 4981 53 4982 1550
rect 4982 53 5028 1550
rect 5028 53 5033 1550
rect 5153 53 5154 1550
rect 5154 53 5200 1550
rect 5200 53 5205 1550
rect 5321 53 5322 1550
rect 5322 53 5368 1550
rect 5368 53 5373 1550
rect 5492 53 5493 1550
rect 5493 53 5539 1550
rect 5539 53 5544 1550
rect 5660 53 5661 1550
rect 5661 53 5707 1550
rect 5707 53 5712 1550
rect 5831 53 5832 1550
rect 5832 53 5878 1550
rect 5878 53 5883 1550
rect 5999 53 6000 1550
rect 6000 53 6046 1550
rect 6046 53 6051 1550
rect 6170 53 6171 1550
rect 6171 53 6217 1550
rect 6217 53 6222 1550
rect 6338 53 6339 1550
rect 6339 53 6385 1550
rect 6385 53 6390 1550
rect 6510 53 6511 1550
rect 6511 53 6557 1550
rect 6557 53 6562 1550
rect 6678 53 6679 1550
rect 6679 53 6725 1550
rect 6725 53 6730 1550
rect 6849 53 6850 1550
rect 6850 53 6896 1550
rect 6896 53 6901 1550
rect 7017 53 7018 1550
rect 7018 53 7064 1550
rect 7064 53 7069 1550
rect 7188 53 7189 1550
rect 7189 53 7235 1550
rect 7235 53 7240 1550
rect 7356 53 7357 1550
rect 7357 53 7403 1550
rect 7403 53 7408 1550
rect 7527 53 7528 1550
rect 7528 53 7574 1550
rect 7574 53 7579 1550
rect 7695 53 7696 1550
rect 7696 53 7742 1550
rect 7742 53 7747 1550
rect 7866 53 7867 1550
rect 7867 53 7913 1550
rect 7913 53 7918 1550
rect 8034 53 8035 1550
rect 8035 53 8081 1550
rect 8081 53 8086 1550
rect 8205 53 8206 1550
rect 8206 53 8252 1550
rect 8252 53 8257 1550
rect 8373 53 8374 1550
rect 8374 53 8420 1550
rect 8420 53 8425 1550
rect 8544 53 8545 1550
rect 8545 53 8591 1550
rect 8591 53 8596 1550
rect 8712 53 8713 1550
rect 8713 53 8759 1550
rect 8759 53 8764 1550
rect 8883 53 8884 1550
rect 8884 53 8930 1550
rect 8930 53 8935 1550
rect 9051 53 9052 1550
rect 9052 53 9098 1550
rect 9098 53 9103 1550
rect 9223 53 9224 1550
rect 9224 53 9270 1550
rect 9270 53 9275 1550
rect 9391 53 9392 1550
rect 9392 53 9438 1550
rect 9438 53 9443 1550
rect 9562 53 9563 1550
rect 9563 53 9609 1550
rect 9609 53 9614 1550
rect 9730 53 9731 1550
rect 9731 53 9777 1550
rect 9777 53 9782 1550
rect 9901 53 9902 1550
rect 9902 53 9948 1550
rect 9948 53 9953 1550
rect 10069 53 10070 1550
rect 10070 53 10116 1550
rect 10116 53 10121 1550
rect 10240 53 10241 1550
rect 10241 53 10287 1550
rect 10287 53 10292 1550
rect 10408 53 10409 1550
rect 10409 53 10455 1550
rect 10455 53 10460 1550
rect 10596 53 10597 1550
rect 10597 53 10643 1550
rect 10643 53 10648 1550
rect 10767 53 10768 1550
rect 10768 53 10814 1550
rect 10814 53 10819 1550
rect 10935 53 10936 1550
rect 10936 53 10982 1550
rect 10982 53 10987 1550
rect 11106 53 11107 1550
rect 11107 53 11153 1550
rect 11153 53 11158 1550
rect 11274 53 11275 1550
rect 11275 53 11321 1550
rect 11321 53 11326 1550
rect 11445 53 11446 1550
rect 11446 53 11492 1550
rect 11492 53 11497 1550
rect 11613 53 11614 1550
rect 11614 53 11660 1550
rect 11660 53 11665 1550
rect 11784 53 11785 1550
rect 11785 53 11831 1550
rect 11831 53 11836 1550
rect 11952 53 11953 1550
rect 11953 53 11999 1550
rect 11999 53 12004 1550
rect 12124 53 12125 1550
rect 12125 53 12171 1550
rect 12171 53 12176 1550
rect 12292 53 12293 1550
rect 12293 53 12339 1550
rect 12339 53 12344 1550
rect 12463 53 12464 1550
rect 12464 53 12510 1550
rect 12510 53 12515 1550
rect 12631 53 12632 1550
rect 12632 53 12678 1550
rect 12678 53 12683 1550
rect 12802 53 12803 1550
rect 12803 53 12849 1550
rect 12849 53 12854 1550
rect 12970 53 12971 1550
rect 12971 53 13017 1550
rect 13017 53 13022 1550
rect 13141 53 13142 1550
rect 13142 53 13188 1550
rect 13188 53 13193 1550
rect 13309 53 13310 1550
rect 13310 53 13356 1550
rect 13356 53 13361 1550
rect 13495 53 13496 1550
rect 13496 53 13542 1550
rect 13542 53 13547 1550
rect 13667 53 13668 1550
rect 13668 53 13714 1550
rect 13714 53 13719 1550
rect 13835 53 13836 1550
rect 13836 53 13882 1550
rect 13882 53 13887 1550
rect 14006 53 14007 1550
rect 14007 53 14053 1550
rect 14053 53 14058 1550
rect 14174 53 14175 1550
rect 14175 53 14221 1550
rect 14221 53 14226 1550
rect 14345 53 14346 1550
rect 14346 53 14392 1550
rect 14392 53 14397 1550
rect 14513 53 14514 1550
rect 14514 53 14560 1550
rect 14560 53 14565 1550
rect 14684 53 14685 1550
rect 14685 53 14731 1550
rect 14731 53 14736 1550
rect 14852 53 14853 1550
rect 14853 53 14899 1550
rect 14899 53 14904 1550
rect 15036 53 15037 1550
rect 15037 53 15083 1550
rect 15083 53 15088 1550
rect 15207 53 15208 1550
rect 15208 53 15254 1550
rect 15254 53 15259 1550
rect 15375 53 15376 1550
rect 15376 53 15422 1550
rect 15422 53 15427 1550
rect 15546 53 15547 1550
rect 15547 53 15593 1550
rect 15593 53 15598 1550
rect 15714 53 15715 1550
rect 15715 53 15761 1550
rect 15761 53 15766 1550
rect 15906 53 15907 1550
rect 15907 53 15953 1550
rect 15953 53 15958 1550
rect 16077 53 16078 1550
rect 16078 53 16124 1550
rect 16124 53 16129 1550
rect 16245 53 16246 1550
rect 16246 53 16292 1550
rect 16292 53 16297 1550
rect 16446 53 16447 1545
rect 16447 53 16493 1545
rect 16493 53 16498 1545
rect 16617 53 16618 1545
rect 16618 53 16664 1545
rect 16664 53 16669 1545
rect 16785 53 16786 1545
rect 16786 53 16832 1545
rect 16832 53 16837 1545
rect 16956 53 16957 1545
rect 16957 53 17003 1545
rect 17003 53 17008 1545
rect 17124 53 17125 1545
rect 17125 53 17171 1545
rect 17171 53 17176 1545
rect 17295 53 17296 1545
rect 17296 53 17342 1545
rect 17342 53 17347 1545
rect 17463 53 17464 1545
rect 17464 53 17510 1545
rect 17510 53 17515 1545
rect 17634 53 17635 1545
rect 17635 53 17681 1545
rect 17681 53 17686 1545
rect 17825 830 17826 1545
rect 17826 830 17872 1545
rect 17872 830 17877 1545
rect 17996 830 17997 1545
rect 17997 830 18043 1545
rect 18043 830 18048 1545
rect 18207 1241 18208 1545
rect 18208 1241 18254 1545
rect 18254 1241 18259 1545
rect 18378 1240 18379 1545
rect 18379 1240 18425 1545
rect 18425 1240 18430 1545
rect 18549 1240 18550 1545
rect 18550 1240 18596 1545
rect 18596 1240 18601 1545
rect 18757 1240 18758 1545
rect 18758 1240 18804 1545
rect 18804 1240 18809 1545
rect 18926 1240 18927 1545
rect 18927 1240 18973 1545
rect 18973 1240 18978 1545
rect 19097 1240 19098 1545
rect 19098 1240 19144 1545
rect 19144 1240 19149 1545
rect 19318 1240 19319 1545
rect 19319 1240 19365 1545
rect 19365 1240 19370 1545
rect 19487 1240 19488 1545
rect 19488 1240 19534 1545
rect 19534 1240 19539 1545
rect 19658 1240 19659 1545
rect 19659 1240 19705 1545
rect 19705 1240 19710 1545
rect 19867 1240 19868 1545
rect 19868 1240 19914 1545
rect 19914 1240 19919 1545
rect 20036 1240 20037 1545
rect 20037 1240 20083 1545
rect 20083 1240 20088 1545
rect 20207 1240 20208 1545
rect 20208 1240 20254 1545
rect 20254 1240 20259 1545
rect 20708 1188 20759 1654
rect 20759 1188 20760 1654
rect 20875 1189 20926 1655
rect 20926 1189 20927 1655
rect 21469 1156 21563 1717
rect 18377 874 18440 943
rect 18552 867 18615 936
rect 18893 866 18956 935
rect 19058 867 19121 936
rect 19412 866 19475 935
rect 19577 867 19640 936
rect 19932 866 19995 935
rect 20097 867 20160 936
rect 20464 866 20527 935
rect 20629 867 20692 936
rect 20982 866 21045 935
rect 21147 867 21210 936
rect 18294 19 18295 734
rect 18295 19 18341 734
rect 18341 19 18346 734
rect 18465 19 18466 734
rect 18466 19 18512 734
rect 18512 19 18517 734
rect 18636 19 18637 734
rect 18637 19 18683 734
rect 18683 19 18688 734
rect 18808 19 18809 734
rect 18809 19 18855 734
rect 18855 19 18860 734
rect 18977 19 18978 734
rect 18978 19 19024 734
rect 19024 19 19029 734
rect 19148 19 19149 734
rect 19149 19 19195 734
rect 19195 19 19200 734
rect 19327 718 19328 734
rect 19328 718 19374 734
rect 19326 624 19327 718
rect 19327 624 19374 718
rect 19327 19 19328 624
rect 19328 19 19374 624
rect 19374 19 19379 734
rect 19496 19 19497 734
rect 19497 19 19543 734
rect 19543 19 19548 734
rect 19667 530 19668 734
rect 19668 530 19714 734
rect 19665 430 19666 530
rect 19666 430 19714 530
rect 19667 19 19668 430
rect 19668 19 19714 430
rect 19714 19 19719 734
rect 19847 717 19848 734
rect 19848 717 19894 734
rect 19846 623 19847 717
rect 19847 623 19894 717
rect 19847 19 19848 623
rect 19848 19 19894 623
rect 19894 19 19899 734
rect 20016 19 20017 734
rect 20017 19 20063 734
rect 20063 19 20068 734
rect 20187 530 20188 734
rect 20188 530 20234 734
rect 20184 430 20185 530
rect 20185 430 20234 530
rect 20187 19 20188 430
rect 20188 19 20234 430
rect 20234 19 20239 734
rect 20379 729 20380 734
rect 20380 729 20426 734
rect 20374 635 20375 729
rect 20375 635 20426 729
rect 20379 19 20380 635
rect 20380 19 20426 635
rect 20426 19 20431 734
rect 20548 19 20549 734
rect 20549 19 20595 734
rect 20595 19 20600 734
rect 20719 530 20720 734
rect 20720 530 20766 734
rect 20715 430 20716 530
rect 20716 430 20766 530
rect 20719 19 20720 430
rect 20720 19 20766 430
rect 20766 19 20771 734
rect 20897 724 20898 734
rect 20898 724 20944 734
rect 20944 724 20949 734
rect 20893 630 20894 724
rect 20894 630 20945 724
rect 20945 630 20949 724
rect 20897 19 20898 630
rect 20898 19 20944 630
rect 20944 19 20949 630
rect 21066 19 21067 734
rect 21067 19 21113 734
rect 21113 19 21118 734
rect 21237 530 21238 734
rect 21238 530 21284 734
rect 21232 430 21233 530
rect 21233 430 21284 530
rect 21237 19 21238 430
rect 21238 19 21284 430
rect 21284 19 21289 734
rect 21462 -23 21556 538
rect 2224 -262 2785 -168
rect 3667 -259 4228 -165
rect 5075 -266 5636 -172
rect 6375 -259 6936 -165
rect 7595 -255 8156 -161
rect 9024 -262 9585 -168
rect 10334 -262 10895 -168
rect 11982 -262 12543 -168
rect 13452 -259 14013 -165
rect 15071 -259 15632 -165
rect 16873 -263 17434 -169
rect 18628 -256 19189 -162
rect 20208 -259 20769 -165
<< metal2 >>
rect 11175 2122 11357 2124
rect 16255 2123 16359 2124
rect 17219 2123 18810 2124
rect 13872 2122 20553 2123
rect 10518 2121 20553 2122
rect 21359 2121 21584 2122
rect -10891 2120 1583 2121
rect 1799 2120 4831 2121
rect 6395 2120 6574 2121
rect 7655 2120 21584 2121
rect -10891 2094 1691 2120
rect -10891 2089 -4309 2094
rect -10891 2087 -6214 2089
rect -10891 2024 -10645 2087
rect -10260 2084 -6214 2087
rect -10260 2024 -9736 2084
rect -10891 2021 -9736 2024
rect -9351 2083 -6214 2084
rect -9351 2082 -7244 2083
rect -9351 2021 -8322 2082
rect -10891 2019 -8322 2021
rect -7937 2020 -7244 2082
rect -6859 2026 -6214 2083
rect -5829 2079 -4309 2089
rect -5829 2026 -5186 2079
rect -6859 2020 -5186 2026
rect -7937 2019 -5186 2020
rect -10891 2016 -5186 2019
rect -4801 2031 -4309 2079
rect -3924 2092 1691 2094
rect -3924 2031 -3355 2092
rect -4801 2029 -3355 2031
rect -2970 2091 1691 2092
rect -2970 2029 -2495 2091
rect -4801 2028 -2495 2029
rect -2110 2089 1691 2091
rect -2110 2087 -162 2089
rect -2110 2028 -1528 2087
rect -4801 2024 -1528 2028
rect -1143 2026 -162 2087
rect 223 2026 876 2089
rect 1261 2026 1691 2089
rect -1143 2024 1691 2026
rect -4801 2016 1691 2024
rect -10891 2015 1691 2016
rect -10892 1990 1691 2015
rect -10892 1846 -10768 1990
rect -10892 1461 -10868 1846
rect -10805 1461 -10768 1846
rect -7643 1767 -7538 1792
rect -7643 1703 -7618 1767
rect -7557 1703 -7538 1767
rect -7643 1675 -7538 1703
rect -3654 1770 -3549 1795
rect -3654 1706 -3629 1770
rect -3568 1706 -3549 1770
rect -3654 1678 -3549 1706
rect -1926 1768 -1821 1793
rect -1926 1704 -1901 1768
rect -1840 1704 -1821 1768
rect -1926 1676 -1821 1704
rect -970 1764 -865 1789
rect -970 1700 -945 1764
rect -884 1700 -865 1764
rect -970 1672 -865 1700
rect -476 1757 -371 1782
rect -476 1693 -451 1757
rect -390 1693 -371 1757
rect -476 1665 -371 1693
rect -47 1742 58 1767
rect -47 1678 -22 1742
rect 39 1678 58 1742
rect -47 1650 58 1678
rect 166 1742 271 1767
rect 166 1678 191 1742
rect 252 1678 271 1742
rect 166 1650 271 1678
rect 504 1743 609 1768
rect 504 1679 529 1743
rect 590 1679 609 1743
rect 504 1651 609 1679
rect 719 1742 824 1767
rect 719 1678 744 1742
rect 805 1678 824 1742
rect 719 1650 824 1678
rect 1074 1740 1179 1765
rect 1074 1676 1099 1740
rect 1160 1676 1179 1740
rect 1074 1648 1179 1676
rect 1287 1742 1392 1767
rect 1287 1678 1312 1742
rect 1373 1678 1392 1742
rect 1287 1650 1392 1678
rect 1569 1740 1691 1990
rect -10892 1249 -10768 1461
rect -10892 864 -10860 1249
rect -10797 864 -10768 1249
rect -10892 451 -10768 864
rect -10892 66 -10855 451
rect -10792 66 -10768 451
rect -10892 -148 -10768 66
rect -10570 1549 -10506 1571
rect -10570 1465 -10561 1549
rect -10570 1399 -10565 1465
rect -10570 50 -10561 1399
rect -10509 50 -10506 1549
rect -10570 30 -10506 50
rect -10401 1549 -10337 1571
rect -10401 222 -10394 1549
rect -10341 222 -10337 1549
rect -10401 138 -10396 222
rect -10340 138 -10337 222
rect -10401 48 -10394 138
rect -10341 48 -10337 138
rect -10401 30 -10337 48
rect -10239 1549 -10175 1571
rect -10239 1469 -10230 1549
rect -10239 1403 -10236 1469
rect -10239 50 -10230 1403
rect -10178 50 -10175 1549
rect -10239 30 -10175 50
rect -10070 1549 -10006 1571
rect -10070 48 -10063 1549
rect -10010 236 -10006 1549
rect -9908 1549 -9844 1571
rect -9908 1468 -9899 1549
rect -9908 1402 -9905 1468
rect -10008 222 -10004 236
rect -10007 138 -10004 222
rect -10008 125 -10004 138
rect -10010 48 -10006 125
rect -10070 30 -10006 48
rect -9908 50 -9899 1402
rect -9847 50 -9844 1549
rect -9908 30 -9844 50
rect -9739 1549 -9675 1571
rect -9739 235 -9732 1549
rect -9739 124 -9734 235
rect -9679 221 -9675 1549
rect -9678 137 -9675 221
rect -9739 48 -9732 124
rect -9679 48 -9675 137
rect -9739 30 -9675 48
rect -9577 1549 -9513 1571
rect -9577 1465 -9568 1549
rect -9577 1399 -9573 1465
rect -9577 50 -9568 1399
rect -9516 50 -9513 1549
rect -9577 30 -9513 50
rect -9408 1549 -9344 1571
rect -9408 234 -9401 1549
rect -9408 123 -9403 234
rect -9348 220 -9344 1549
rect -9347 136 -9344 220
rect -9408 48 -9401 123
rect -9348 48 -9344 136
rect -9408 30 -9344 48
rect -9244 1549 -9180 1571
rect -9244 1468 -9235 1549
rect -9183 1468 -9180 1549
rect -9244 1402 -9238 1468
rect -9182 1402 -9180 1468
rect -9244 50 -9235 1402
rect -9183 50 -9180 1402
rect -9244 30 -9180 50
rect -9075 1549 -9011 1571
rect -9075 237 -9068 1549
rect -9075 126 -9070 237
rect -9015 223 -9011 1549
rect -9014 139 -9011 223
rect -9075 48 -9068 126
rect -9015 48 -9011 139
rect -9075 30 -9011 48
rect -8913 1549 -8849 1571
rect -8913 1465 -8904 1549
rect -8852 1465 -8849 1549
rect -8913 1399 -8907 1465
rect -8851 1399 -8849 1465
rect -8913 50 -8904 1399
rect -8852 50 -8849 1399
rect -8913 30 -8849 50
rect -8744 1549 -8680 1571
rect -8744 237 -8737 1549
rect -8744 126 -8739 237
rect -8684 223 -8680 1549
rect -8683 139 -8680 223
rect -8744 48 -8737 126
rect -8684 48 -8680 139
rect -8744 30 -8680 48
rect -8582 1549 -8518 1571
rect -8582 1466 -8573 1549
rect -8582 1400 -8577 1466
rect -8582 50 -8573 1400
rect -8521 50 -8518 1549
rect -8582 30 -8518 50
rect -8413 1549 -8349 1571
rect -8413 239 -8406 1549
rect -8413 128 -8408 239
rect -8353 225 -8349 1549
rect -8352 141 -8349 225
rect -8413 48 -8406 128
rect -8353 48 -8349 141
rect -8413 30 -8349 48
rect -8251 1549 -8187 1571
rect -8251 1467 -8242 1549
rect -8251 1401 -8246 1467
rect -8251 50 -8242 1401
rect -8190 50 -8187 1549
rect -8251 30 -8187 50
rect -8082 1549 -8018 1571
rect -8082 241 -8075 1549
rect -8022 241 -8018 1549
rect -7919 1549 -7855 1571
rect -7919 1467 -7910 1549
rect -7919 1401 -7915 1467
rect -8082 130 -8076 241
rect -8021 227 -8017 241
rect -8020 143 -8017 227
rect -8021 130 -8017 143
rect -8082 48 -8075 130
rect -8022 48 -8018 130
rect -8082 30 -8018 48
rect -7919 50 -7910 1401
rect -7858 50 -7855 1549
rect -7919 30 -7855 50
rect -7750 1549 -7686 1571
rect -7750 241 -7743 1549
rect -7750 130 -7745 241
rect -7690 227 -7686 1549
rect -7689 143 -7686 227
rect -7750 48 -7743 130
rect -7690 48 -7686 143
rect -7750 30 -7686 48
rect -7588 1549 -7524 1571
rect -7588 1466 -7579 1549
rect -7588 1400 -7584 1466
rect -7588 50 -7579 1400
rect -7527 50 -7524 1549
rect -7588 30 -7524 50
rect -7419 1549 -7355 1571
rect -7419 241 -7412 1549
rect -7359 241 -7355 1549
rect -7257 1549 -7193 1571
rect -7257 1465 -7248 1549
rect -7257 1399 -7253 1465
rect -7419 130 -7413 241
rect -7358 227 -7354 241
rect -7357 143 -7354 227
rect -7358 130 -7354 143
rect -7419 48 -7412 130
rect -7359 48 -7355 130
rect -7419 30 -7355 48
rect -7257 50 -7248 1399
rect -7196 50 -7193 1549
rect -7257 30 -7193 50
rect -7088 1549 -7024 1571
rect -7088 241 -7081 1549
rect -7028 241 -7024 1549
rect -6926 1549 -6862 1571
rect -6926 1462 -6917 1549
rect -6926 1396 -6921 1462
rect -7088 130 -7082 241
rect -7027 227 -7023 241
rect -7026 143 -7023 227
rect -7027 130 -7023 143
rect -7088 48 -7081 130
rect -7028 48 -7024 130
rect -7088 30 -7024 48
rect -6926 50 -6917 1396
rect -6865 50 -6862 1549
rect -6926 30 -6862 50
rect -6757 1549 -6693 1571
rect -6757 241 -6750 1549
rect -6757 130 -6752 241
rect -6697 227 -6693 1549
rect -6696 143 -6693 227
rect -6757 48 -6750 130
rect -6697 48 -6693 143
rect -6757 30 -6693 48
rect -6593 1549 -6529 1571
rect -6593 1463 -6584 1549
rect -6593 1397 -6589 1463
rect -6593 50 -6584 1397
rect -6532 50 -6529 1549
rect -6593 30 -6529 50
rect -6424 1549 -6360 1571
rect -6424 241 -6417 1549
rect -6424 130 -6419 241
rect -6364 227 -6360 1549
rect -6363 143 -6360 227
rect -6424 48 -6417 130
rect -6364 48 -6360 143
rect -6424 30 -6360 48
rect -6262 1549 -6198 1571
rect -6262 1462 -6253 1549
rect -6201 1462 -6198 1549
rect -6262 1396 -6256 1462
rect -6200 1396 -6198 1462
rect -6262 50 -6253 1396
rect -6201 50 -6198 1396
rect -6262 30 -6198 50
rect -6093 1549 -6029 1571
rect -6093 241 -6086 1549
rect -6093 130 -6088 241
rect -6033 227 -6029 1549
rect -6032 143 -6029 227
rect -6093 48 -6086 130
rect -6033 48 -6029 143
rect -6093 30 -6029 48
rect -5931 1549 -5867 1571
rect -5931 1464 -5922 1549
rect -5931 1398 -5926 1464
rect -5931 50 -5922 1398
rect -5870 50 -5867 1549
rect -5931 30 -5867 50
rect -5762 1549 -5698 1571
rect -5762 48 -5755 1549
rect -5702 251 -5698 1549
rect -5600 1549 -5536 1571
rect -5600 1462 -5591 1549
rect -5600 1396 -5595 1462
rect -5700 237 -5696 251
rect -5699 153 -5696 237
rect -5700 140 -5696 153
rect -5702 48 -5698 140
rect -5762 30 -5698 48
rect -5600 50 -5591 1396
rect -5539 50 -5536 1549
rect -5600 30 -5536 50
rect -5431 1549 -5367 1571
rect -5431 251 -5424 1549
rect -5431 140 -5426 251
rect -5371 237 -5367 1549
rect -5370 153 -5367 237
rect -5431 48 -5424 140
rect -5371 48 -5367 153
rect -5431 30 -5367 48
rect -5267 1549 -5203 1571
rect -5267 1462 -5258 1549
rect -5267 1396 -5263 1462
rect -5267 50 -5258 1396
rect -5206 50 -5203 1549
rect -5267 30 -5203 50
rect -5098 1549 -5034 1571
rect -5098 240 -5091 1549
rect -5038 240 -5034 1549
rect -5098 161 -5094 240
rect -5037 161 -5034 240
rect -5098 48 -5091 161
rect -5038 48 -5034 161
rect -5098 30 -5034 48
rect -4936 1549 -4872 1571
rect -4936 1462 -4927 1549
rect -4936 1396 -4932 1462
rect -4936 50 -4927 1396
rect -4875 50 -4872 1549
rect -4936 30 -4872 50
rect -4767 1549 -4703 1571
rect -4767 240 -4760 1549
rect -4707 252 -4703 1549
rect -4605 1549 -4541 1571
rect -4605 1463 -4596 1549
rect -4605 1397 -4602 1463
rect -4705 240 -4701 252
rect -4767 161 -4761 240
rect -4704 161 -4701 240
rect -4767 48 -4760 161
rect -4705 150 -4701 161
rect -4707 48 -4703 150
rect -4767 30 -4703 48
rect -4605 50 -4596 1397
rect -4544 50 -4541 1549
rect -4605 30 -4541 50
rect -4436 1549 -4372 1571
rect -4436 252 -4429 1549
rect -4376 252 -4372 1549
rect -4274 1549 -4210 1571
rect -4274 1462 -4265 1549
rect -4274 1396 -4271 1462
rect -4436 240 -4430 252
rect -4375 240 -4371 252
rect -4436 161 -4431 240
rect -4374 161 -4371 240
rect -4436 150 -4430 161
rect -4375 150 -4371 161
rect -4436 48 -4429 150
rect -4376 48 -4372 150
rect -4436 30 -4372 48
rect -4274 50 -4265 1396
rect -4213 50 -4210 1549
rect -4274 30 -4210 50
rect -4105 1549 -4041 1571
rect -4105 252 -4098 1549
rect -4105 240 -4100 252
rect -4045 240 -4041 1549
rect -4105 161 -4101 240
rect -4044 161 -4041 240
rect -4105 150 -4100 161
rect -4105 48 -4098 150
rect -4045 48 -4041 161
rect -4105 30 -4041 48
rect -3941 1549 -3877 1571
rect -3941 1463 -3932 1549
rect -3941 1397 -3936 1463
rect -3941 50 -3932 1397
rect -3880 50 -3877 1549
rect -3941 30 -3877 50
rect -3772 1549 -3708 1571
rect -3772 252 -3765 1549
rect -3712 252 -3708 1549
rect -3610 1549 -3546 1571
rect -3610 1464 -3601 1549
rect -3610 1398 -3606 1464
rect -3772 240 -3766 252
rect -3711 240 -3707 252
rect -3772 161 -3767 240
rect -3710 161 -3707 240
rect -3772 150 -3766 161
rect -3711 150 -3707 161
rect -3772 48 -3765 150
rect -3712 48 -3708 150
rect -3772 30 -3708 48
rect -3610 50 -3601 1398
rect -3549 50 -3546 1549
rect -3610 30 -3546 50
rect -3441 1549 -3377 1571
rect -3441 252 -3434 1549
rect -3381 252 -3377 1549
rect -3279 1549 -3215 1571
rect -3279 1463 -3270 1549
rect -3279 1397 -3275 1463
rect -3441 240 -3435 252
rect -3380 240 -3376 252
rect -3441 161 -3436 240
rect -3379 161 -3376 240
rect -3441 150 -3435 161
rect -3380 150 -3376 161
rect -3441 48 -3434 150
rect -3381 48 -3377 150
rect -3441 30 -3377 48
rect -3279 50 -3270 1397
rect -3218 50 -3215 1549
rect -3279 30 -3215 50
rect -3110 1549 -3046 1571
rect -3110 251 -3103 1549
rect -3110 239 -3105 251
rect -3050 239 -3046 1549
rect -3110 160 -3106 239
rect -3049 160 -3046 239
rect -3110 149 -3105 160
rect -3110 48 -3103 149
rect -3050 48 -3046 160
rect -3110 30 -3046 48
rect -2948 1549 -2884 1571
rect -2948 1464 -2939 1549
rect -2948 1398 -2944 1464
rect -2948 50 -2939 1398
rect -2887 50 -2884 1549
rect -2948 30 -2884 50
rect -2779 1549 -2715 1571
rect -2779 252 -2772 1549
rect -2779 240 -2774 252
rect -2719 240 -2715 1549
rect -2779 161 -2775 240
rect -2718 161 -2715 240
rect -2779 150 -2774 161
rect -2779 48 -2772 150
rect -2719 48 -2715 161
rect -2779 30 -2715 48
rect -2618 1549 -2554 1571
rect -2618 1465 -2609 1549
rect -2618 1399 -2614 1465
rect -2618 50 -2609 1399
rect -2557 50 -2554 1549
rect -2618 30 -2554 50
rect -2449 1549 -2385 1571
rect -2449 252 -2442 1549
rect -2389 252 -2385 1549
rect -2287 1549 -2223 1571
rect -2287 1464 -2278 1549
rect -2287 1398 -2282 1464
rect -2449 240 -2443 252
rect -2388 240 -2384 252
rect -2449 161 -2444 240
rect -2387 161 -2384 240
rect -2449 150 -2443 161
rect -2388 150 -2384 161
rect -2449 48 -2442 150
rect -2389 48 -2385 150
rect -2449 30 -2385 48
rect -2287 50 -2278 1398
rect -2226 50 -2223 1549
rect -2287 30 -2223 50
rect -2118 1549 -2054 1571
rect -2118 252 -2111 1549
rect -2058 252 -2054 1549
rect -1956 1549 -1892 1571
rect -1956 1463 -1947 1549
rect -1956 1397 -1953 1463
rect -2118 240 -2112 252
rect -2057 240 -2053 252
rect -2118 161 -2113 240
rect -2056 161 -2053 240
rect -2118 150 -2112 161
rect -2057 150 -2053 161
rect -2118 48 -2111 150
rect -2058 48 -2054 150
rect -2118 30 -2054 48
rect -1956 50 -1947 1397
rect -1895 50 -1892 1549
rect -1956 30 -1892 50
rect -1787 1549 -1723 1571
rect -1787 252 -1780 1549
rect -1787 240 -1782 252
rect -1727 240 -1723 1549
rect -1787 161 -1783 240
rect -1726 161 -1723 240
rect -1787 150 -1782 161
rect -1787 48 -1780 150
rect -1727 48 -1723 161
rect -1787 30 -1723 48
rect -1625 1549 -1561 1571
rect -1625 1464 -1616 1549
rect -1625 1398 -1621 1464
rect -1625 50 -1616 1398
rect -1564 50 -1561 1549
rect -1625 30 -1561 50
rect -1456 1549 -1392 1571
rect -1456 252 -1449 1549
rect -1396 252 -1392 1549
rect -1293 1549 -1229 1571
rect -1293 1463 -1284 1549
rect -1293 1397 -1289 1463
rect -1456 240 -1450 252
rect -1395 240 -1391 252
rect -1456 161 -1451 240
rect -1394 161 -1391 240
rect -1456 150 -1450 161
rect -1395 150 -1391 161
rect -1456 48 -1449 150
rect -1396 48 -1392 150
rect -1456 30 -1392 48
rect -1293 50 -1284 1397
rect -1232 50 -1229 1549
rect -1293 30 -1229 50
rect -1124 1549 -1060 1571
rect -1124 252 -1117 1549
rect -1124 240 -1119 252
rect -1064 240 -1060 1549
rect -1124 161 -1120 240
rect -1063 161 -1060 240
rect -1124 150 -1119 161
rect -1124 48 -1117 150
rect -1064 48 -1060 161
rect -1124 30 -1060 48
rect -962 1549 -898 1571
rect -962 1465 -953 1549
rect -962 1399 -957 1465
rect -962 50 -953 1399
rect -901 50 -898 1549
rect -962 30 -898 50
rect -793 1549 -729 1571
rect -793 252 -786 1549
rect -733 252 -729 1549
rect -631 1549 -567 1571
rect -631 1467 -622 1549
rect -631 1401 -626 1467
rect -793 240 -787 252
rect -732 240 -728 252
rect -793 161 -788 240
rect -731 161 -728 240
rect -793 150 -787 161
rect -732 150 -728 161
rect -793 48 -786 150
rect -733 48 -729 150
rect -793 30 -729 48
rect -631 50 -622 1401
rect -570 50 -567 1549
rect -631 30 -567 50
rect -462 1549 -398 1571
rect -462 252 -455 1549
rect -402 252 -398 1549
rect -296 1549 -232 1571
rect -296 1468 -289 1549
rect -236 1468 -232 1549
rect -296 1402 -290 1468
rect -233 1402 -232 1468
rect -462 240 -456 252
rect -401 240 -397 252
rect -462 161 -457 240
rect -400 161 -397 240
rect -462 150 -456 161
rect -401 150 -397 161
rect -462 48 -455 150
rect -402 48 -398 150
rect -462 30 -398 48
rect -296 48 -289 1402
rect -236 48 -232 1402
rect -89 1549 -25 1571
rect -89 252 -80 1549
rect -90 240 -85 252
rect -90 161 -86 240
rect -90 150 -85 161
rect -296 30 -232 48
rect -89 50 -80 150
rect -28 50 -25 1549
rect -89 30 -25 50
rect 80 1549 144 1571
rect 80 1451 87 1549
rect 140 1451 144 1549
rect 80 1395 83 1451
rect 142 1395 144 1451
rect 80 48 87 1395
rect 140 48 144 1395
rect 80 30 144 48
rect 246 1549 310 1571
rect 246 252 253 1549
rect 306 252 310 1549
rect 464 1549 528 1571
rect 464 252 473 1549
rect 246 240 251 252
rect 246 161 250 240
rect 246 150 251 161
rect 308 150 310 252
rect 462 240 467 252
rect 462 161 466 240
rect 462 150 467 161
rect 246 48 253 150
rect 306 48 310 150
rect 246 30 310 48
rect 464 50 473 150
rect 525 50 528 1549
rect 464 30 528 50
rect 633 1549 697 1571
rect 633 1452 640 1549
rect 693 1452 697 1549
rect 633 1396 637 1452
rect 696 1396 697 1452
rect 633 48 640 1396
rect 693 48 697 1396
rect 633 30 697 48
rect 799 1549 863 1571
rect 799 244 806 1549
rect 859 244 863 1549
rect 799 158 805 244
rect 862 158 863 244
rect 799 48 806 158
rect 859 48 863 158
rect 799 30 863 48
rect 1033 1549 1097 1571
rect 1033 255 1042 1549
rect 1094 255 1097 1549
rect 1202 1549 1266 1571
rect 1202 1452 1209 1549
rect 1262 1452 1266 1549
rect 1202 1396 1206 1452
rect 1265 1396 1266 1452
rect 1033 245 1041 255
rect 1094 245 1098 255
rect 1033 159 1040 245
rect 1097 159 1098 245
rect 1033 150 1041 159
rect 1094 150 1098 159
rect 1033 50 1042 150
rect 1094 50 1097 150
rect 1033 30 1097 50
rect 1202 48 1209 1396
rect 1262 48 1266 1396
rect 1202 30 1266 48
rect 1368 1549 1432 1571
rect 1368 245 1375 1549
rect 1428 245 1432 1549
rect 1368 159 1374 245
rect 1431 159 1432 245
rect 1368 48 1375 159
rect 1428 48 1432 159
rect 1368 30 1432 48
rect 1569 1355 1600 1740
rect 1663 1355 1691 1740
rect 1569 971 1691 1355
rect 1569 586 1599 971
rect 1662 586 1691 971
rect 1569 379 1691 586
rect 1569 -6 1598 379
rect 1661 -6 1691 379
rect 1569 -148 1691 -6
rect -10893 -175 1691 -148
rect -10893 -182 -8567 -175
rect -10893 -245 -10444 -182
rect -10059 -183 -8567 -182
rect -10059 -245 -9441 -183
rect -10893 -246 -9441 -245
rect -9056 -238 -8567 -183
rect -8182 -179 626 -175
rect -8182 -181 -4325 -179
rect -8182 -238 -7658 -181
rect -9056 -244 -7658 -238
rect -7273 -184 -4325 -181
rect -7273 -186 -5464 -184
rect -7273 -244 -6670 -186
rect -9056 -246 -6670 -244
rect -10893 -249 -6670 -246
rect -6285 -247 -5464 -186
rect -5079 -242 -4325 -184
rect -3940 -185 626 -179
rect -3940 -242 -3208 -185
rect -5079 -247 -3208 -242
rect -6285 -248 -3208 -247
rect -2823 -191 -1140 -185
rect -2823 -248 -2261 -191
rect -6285 -249 -2261 -248
rect -10893 -254 -2261 -249
rect -1876 -248 -1140 -191
rect -755 -248 -270 -185
rect 115 -238 626 -185
rect 1011 -238 1691 -175
rect 115 -248 1691 -238
rect -1876 -254 1691 -248
rect -10893 -280 1691 -254
rect 1799 2110 21584 2120
rect 1799 2107 17623 2110
rect 1799 2106 6883 2107
rect 1799 2101 3780 2106
rect 1799 2007 2184 2101
rect 2745 2012 3780 2101
rect 4341 2099 6883 2106
rect 4341 2012 5230 2099
rect 2745 2007 5230 2012
rect 1799 2005 5230 2007
rect 5791 2013 6883 2099
rect 7444 2104 9727 2107
rect 7444 2013 8198 2104
rect 5791 2010 8198 2013
rect 8759 2013 9727 2104
rect 10288 2106 17623 2107
rect 10288 2102 16308 2106
rect 10288 2013 11480 2102
rect 8759 2010 11480 2013
rect 5791 2008 11480 2010
rect 12041 2100 16308 2102
rect 12041 2098 14532 2100
rect 12041 2008 12864 2098
rect 5791 2005 12864 2008
rect 1799 2004 12864 2005
rect 13425 2006 14532 2098
rect 15093 2012 16308 2100
rect 16869 2016 17623 2106
rect 18184 2107 21584 2110
rect 18184 2016 19309 2107
rect 16869 2013 19309 2016
rect 19870 2100 21584 2107
rect 19870 2013 20507 2100
rect 16869 2012 20507 2013
rect 15093 2006 20507 2012
rect 21068 2006 21584 2100
rect 13425 2004 21584 2006
rect 1799 1991 21584 2004
rect 1799 1990 14000 1991
rect 1799 1716 1919 1990
rect 4800 1989 7665 1990
rect 8848 1989 9027 1990
rect 12591 1989 12773 1990
rect 13819 1989 14000 1990
rect 14507 1989 14688 1991
rect 12591 1988 12769 1989
rect 13820 1988 14000 1989
rect 14508 1988 14688 1989
rect 15140 1988 15319 1991
rect 15478 1988 15657 1991
rect 18757 1990 20553 1991
rect 21359 1990 21584 1991
rect 13820 1987 13998 1988
rect 14508 1987 14686 1988
rect 15140 1987 15317 1988
rect 15478 1987 15655 1988
rect 20768 1857 20880 1872
rect 1799 1361 1827 1716
rect 1899 1361 1919 1716
rect 3221 1782 3399 1801
rect 3221 1712 3258 1782
rect 3370 1712 3399 1782
rect 3221 1690 3399 1712
rect 6396 1782 6574 1801
rect 6396 1712 6433 1782
rect 6545 1712 6574 1782
rect 6396 1690 6574 1712
rect 8849 1781 9027 1800
rect 8849 1711 8886 1781
rect 8998 1711 9027 1781
rect 8849 1689 9027 1711
rect 11175 1784 11353 1803
rect 11175 1714 11212 1784
rect 11324 1714 11353 1784
rect 11175 1692 11353 1714
rect 12591 1780 12769 1799
rect 20768 1798 20781 1857
rect 20865 1798 20880 1857
rect 12591 1710 12628 1780
rect 12740 1710 12769 1780
rect 12591 1688 12769 1710
rect 13820 1779 13998 1798
rect 13820 1709 13857 1779
rect 13969 1709 13998 1779
rect 13820 1687 13998 1709
rect 14508 1779 14686 1798
rect 14508 1709 14545 1779
rect 14657 1709 14686 1779
rect 14508 1687 14686 1709
rect 15140 1779 15317 1798
rect 15140 1709 15176 1779
rect 15288 1709 15317 1779
rect 15140 1688 15317 1709
rect 15478 1779 15655 1798
rect 20768 1781 20880 1798
rect 15478 1709 15514 1779
rect 15626 1709 15655 1779
rect 16725 1771 17612 1773
rect 16725 1770 17616 1771
rect 17789 1770 17978 1771
rect 16725 1769 17978 1770
rect 18259 1769 18348 1771
rect 18431 1770 18520 1771
rect 18803 1770 18892 1771
rect 18954 1770 19482 1771
rect 18431 1769 20175 1770
rect 15478 1688 15655 1709
rect 15930 1748 16043 1763
rect 15930 1689 15943 1748
rect 16027 1689 16043 1748
rect 15930 1670 16043 1689
rect 16153 1748 16265 1763
rect 16153 1689 16166 1748
rect 16250 1689 16265 1748
rect 16153 1670 16265 1689
rect 16725 1752 20175 1769
rect 16725 1695 16751 1752
rect 16870 1746 20175 1752
rect 16870 1695 17262 1746
rect 16725 1692 17262 1695
rect 17380 1741 20175 1746
rect 17380 1692 17542 1741
rect 16725 1677 17542 1692
rect 17236 1674 17397 1677
rect 17527 1673 17542 1677
rect 17599 1678 17904 1741
rect 17599 1673 17616 1678
rect 17789 1677 17904 1678
rect 17527 1648 17616 1673
rect 17889 1673 17904 1677
rect 17961 1679 18274 1741
rect 17961 1673 17978 1679
rect 17889 1648 17978 1673
rect 18259 1673 18274 1679
rect 18331 1679 18446 1741
rect 18331 1673 18348 1679
rect 18259 1648 18348 1673
rect 18431 1673 18446 1679
rect 18503 1678 18818 1741
rect 18503 1673 18520 1678
rect 18431 1648 18520 1673
rect 18803 1673 18818 1678
rect 18875 1678 18991 1741
rect 18875 1673 18892 1678
rect 18803 1648 18892 1673
rect 18976 1673 18991 1678
rect 19048 1678 19379 1741
rect 19048 1673 19065 1678
rect 18976 1648 19065 1673
rect 19364 1673 19379 1678
rect 19436 1678 19552 1741
rect 19436 1673 19453 1678
rect 19364 1648 19453 1673
rect 19537 1673 19552 1678
rect 19609 1679 19928 1741
rect 19609 1673 19626 1679
rect 19912 1678 19928 1679
rect 19537 1648 19626 1673
rect 19913 1673 19928 1678
rect 19985 1678 20101 1741
rect 19985 1673 20002 1678
rect 19913 1648 20002 1673
rect 20086 1673 20101 1678
rect 20158 1673 20175 1741
rect 21427 1717 21584 1990
rect 20086 1648 20175 1673
rect 20698 1654 20771 1713
rect 1799 920 1919 1361
rect 1799 565 1824 920
rect 1896 565 1919 920
rect 1799 352 1919 565
rect 1799 -3 1820 352
rect 1892 -3 1919 352
rect 2058 1550 2121 1572
rect 2058 1531 2067 1550
rect 2058 1457 2061 1531
rect 2058 53 2067 1457
rect 2119 53 2121 1550
rect 2058 30 2121 53
rect 2230 1550 2293 1572
rect 2230 170 2239 1550
rect 2230 53 2239 80
rect 2291 53 2293 1550
rect 2230 30 2293 53
rect 2398 1550 2461 1572
rect 2398 1529 2407 1550
rect 2398 1455 2401 1529
rect 2398 53 2407 1455
rect 2459 53 2461 1550
rect 2398 30 2461 53
rect 2569 1550 2632 1572
rect 2569 170 2578 1550
rect 2569 80 2570 170
rect 2569 53 2578 80
rect 2630 53 2632 1550
rect 2569 30 2632 53
rect 2737 1550 2800 1572
rect 2737 1531 2746 1550
rect 2737 1457 2741 1531
rect 2737 53 2746 1457
rect 2798 53 2800 1550
rect 2737 30 2800 53
rect 2908 1550 2971 1572
rect 2908 170 2917 1550
rect 2969 170 2971 1550
rect 2908 80 2910 170
rect 2970 80 2971 170
rect 2908 53 2917 80
rect 2969 53 2971 80
rect 2908 30 2971 53
rect 3076 1550 3139 1572
rect 3076 1534 3085 1550
rect 3076 1460 3080 1534
rect 3076 53 3085 1460
rect 3137 53 3139 1550
rect 3076 30 3139 53
rect 3247 1550 3310 1572
rect 3247 170 3256 1550
rect 3308 170 3310 1550
rect 3247 80 3250 170
rect 3247 53 3256 80
rect 3308 53 3310 80
rect 3247 30 3310 53
rect 3415 1550 3478 1572
rect 3415 1531 3424 1550
rect 3476 1531 3478 1550
rect 3415 1457 3420 1531
rect 3477 1457 3478 1531
rect 3415 53 3424 1457
rect 3476 53 3478 1457
rect 3415 30 3478 53
rect 3587 1550 3650 1572
rect 3587 170 3596 1550
rect 3648 170 3650 1550
rect 3587 80 3590 170
rect 3587 53 3596 80
rect 3648 53 3650 80
rect 3587 30 3650 53
rect 3755 1550 3818 1572
rect 3755 1532 3764 1550
rect 3755 1458 3759 1532
rect 3755 53 3764 1458
rect 3816 53 3818 1550
rect 3755 30 3818 53
rect 3926 1550 3989 1572
rect 3926 178 3935 1550
rect 3987 178 3989 1550
rect 3926 80 3928 178
rect 3988 170 3989 178
rect 4094 1550 4157 1572
rect 4094 1532 4103 1550
rect 4094 1458 4096 1532
rect 3988 80 3990 170
rect 3926 53 3935 80
rect 3987 53 3989 80
rect 3926 30 3989 53
rect 4094 53 4103 1458
rect 4155 53 4157 1550
rect 4094 30 4157 53
rect 4265 1550 4328 1572
rect 4265 168 4274 1550
rect 4326 168 4328 1550
rect 4265 78 4267 168
rect 4327 78 4328 168
rect 4265 53 4274 78
rect 4326 53 4328 78
rect 4265 30 4328 53
rect 4433 1550 4496 1572
rect 4433 1535 4442 1550
rect 4433 1461 4435 1535
rect 4433 53 4442 1461
rect 4494 53 4496 1550
rect 4433 30 4496 53
rect 4604 1550 4667 1572
rect 4604 172 4613 1550
rect 4665 172 4667 1550
rect 4604 82 4606 172
rect 4666 82 4667 172
rect 4604 53 4613 82
rect 4665 53 4667 82
rect 4604 30 4667 53
rect 4772 1550 4835 1572
rect 4772 1535 4781 1550
rect 4772 1461 4773 1535
rect 4772 53 4781 1461
rect 4833 53 4835 1550
rect 4772 30 4835 53
rect 4972 1550 5035 1572
rect 4972 179 4981 1550
rect 4972 108 4976 179
rect 4972 53 4981 108
rect 5033 53 5035 1550
rect 4972 30 5035 53
rect 5144 1550 5207 1572
rect 5144 1530 5153 1550
rect 5144 1458 5148 1530
rect 5144 53 5153 1458
rect 5205 53 5207 1550
rect 5144 30 5207 53
rect 5312 1550 5375 1572
rect 5312 178 5321 1550
rect 5312 107 5314 178
rect 5312 53 5321 107
rect 5373 53 5375 1550
rect 5312 30 5375 53
rect 5483 1550 5546 1572
rect 5483 1530 5492 1550
rect 5483 1458 5487 1530
rect 5483 53 5492 1458
rect 5544 53 5546 1550
rect 5483 30 5546 53
rect 5651 1550 5714 1572
rect 5651 177 5660 1550
rect 5651 106 5654 177
rect 5651 53 5660 106
rect 5712 53 5714 1550
rect 5651 30 5714 53
rect 5822 1550 5885 1572
rect 5822 1530 5831 1550
rect 5822 1458 5826 1530
rect 5822 53 5831 1458
rect 5883 53 5885 1550
rect 5822 30 5885 53
rect 5990 1550 6053 1572
rect 5990 177 5999 1550
rect 5990 106 5994 177
rect 5990 53 5999 106
rect 6051 53 6053 1550
rect 5990 30 6053 53
rect 6161 1550 6224 1572
rect 6161 1530 6170 1550
rect 6222 1530 6224 1550
rect 6161 1458 6167 1530
rect 6223 1458 6224 1530
rect 6161 53 6170 1458
rect 6222 53 6224 1458
rect 6161 30 6224 53
rect 6329 1550 6392 1572
rect 6329 175 6338 1550
rect 6329 104 6333 175
rect 6329 53 6338 104
rect 6390 53 6392 1550
rect 6329 30 6392 53
rect 6501 1550 6564 1572
rect 6501 1528 6510 1550
rect 6501 1456 6504 1528
rect 6501 53 6510 1456
rect 6562 53 6564 1550
rect 6501 30 6564 53
rect 6669 1550 6732 1572
rect 6669 175 6678 1550
rect 6669 104 6673 175
rect 6669 53 6678 104
rect 6730 53 6732 1550
rect 6669 30 6732 53
rect 6840 1550 6903 1572
rect 6840 1528 6849 1550
rect 6840 1456 6844 1528
rect 6840 53 6849 1456
rect 6901 53 6903 1550
rect 6840 30 6903 53
rect 7008 1550 7071 1572
rect 7008 174 7017 1550
rect 7008 103 7012 174
rect 7008 53 7017 103
rect 7069 53 7071 1550
rect 7008 30 7071 53
rect 7179 1550 7242 1572
rect 7179 1529 7188 1550
rect 7179 1457 7183 1529
rect 7179 53 7188 1457
rect 7240 53 7242 1550
rect 7179 30 7242 53
rect 7347 1550 7410 1572
rect 7347 175 7356 1550
rect 7347 104 7351 175
rect 7347 53 7356 104
rect 7408 53 7410 1550
rect 7347 30 7410 53
rect 7518 1550 7581 1572
rect 7518 1529 7527 1550
rect 7518 1457 7523 1529
rect 7518 53 7527 1457
rect 7579 53 7581 1550
rect 7518 30 7581 53
rect 7686 1550 7749 1572
rect 7686 174 7695 1550
rect 7686 103 7690 174
rect 7686 53 7695 103
rect 7747 53 7749 1550
rect 7686 30 7749 53
rect 7857 1550 7920 1572
rect 7857 1210 7866 1550
rect 7918 1210 7920 1550
rect 7857 1137 7861 1210
rect 7919 1137 7920 1210
rect 7857 53 7866 1137
rect 7918 53 7920 1137
rect 7857 30 7920 53
rect 8025 1550 8088 1572
rect 8025 175 8034 1550
rect 8025 104 8028 175
rect 8025 53 8034 104
rect 8086 53 8088 1550
rect 8025 30 8088 53
rect 8196 1550 8259 1572
rect 8196 1210 8205 1550
rect 8257 1210 8259 1550
rect 8196 1137 8201 1210
rect 8196 53 8205 1137
rect 8257 53 8259 1137
rect 8196 30 8259 53
rect 8364 1550 8427 1572
rect 8364 174 8373 1550
rect 8364 103 8366 174
rect 8364 53 8373 103
rect 8425 53 8427 1550
rect 8364 30 8427 53
rect 8535 1550 8598 1572
rect 8535 1209 8544 1550
rect 8596 1209 8598 1550
rect 8535 1136 8539 1209
rect 8597 1136 8598 1209
rect 8535 53 8544 1136
rect 8596 53 8598 1136
rect 8535 30 8598 53
rect 8703 1550 8766 1572
rect 8703 182 8712 1550
rect 8703 111 8706 182
rect 8703 53 8712 111
rect 8764 53 8766 1550
rect 8703 30 8766 53
rect 8874 1550 8937 1572
rect 8874 1213 8883 1550
rect 8935 1213 8937 1550
rect 8874 1140 8879 1213
rect 8874 53 8883 1140
rect 8935 53 8937 1140
rect 8874 30 8937 53
rect 9042 1550 9105 1572
rect 9042 189 9051 1550
rect 9042 118 9047 189
rect 9042 53 9051 118
rect 9103 53 9105 1550
rect 9042 30 9105 53
rect 9214 1550 9277 1572
rect 9214 1214 9223 1550
rect 9214 1141 9217 1214
rect 9214 53 9223 1141
rect 9275 53 9277 1550
rect 9214 30 9277 53
rect 9382 1550 9445 1572
rect 9382 183 9391 1550
rect 9382 112 9386 183
rect 9382 53 9391 112
rect 9443 53 9445 1550
rect 9382 30 9445 53
rect 9553 1550 9616 1572
rect 9553 1214 9562 1550
rect 9553 1141 9555 1214
rect 9553 53 9562 1141
rect 9614 53 9616 1550
rect 9553 30 9616 53
rect 9721 1550 9784 1572
rect 9721 187 9730 1550
rect 9721 116 9726 187
rect 9721 53 9730 116
rect 9782 53 9784 1550
rect 9721 30 9784 53
rect 9892 1550 9955 1572
rect 9892 1214 9901 1550
rect 9892 1141 9894 1214
rect 9892 53 9901 1141
rect 9953 53 9955 1550
rect 9892 30 9955 53
rect 10060 1550 10123 1572
rect 10060 186 10069 1550
rect 10060 115 10065 186
rect 10060 53 10069 115
rect 10121 53 10123 1550
rect 10060 30 10123 53
rect 10231 1550 10294 1572
rect 10231 1213 10240 1550
rect 10231 1140 10234 1213
rect 10231 53 10240 1140
rect 10292 53 10294 1550
rect 10231 30 10294 53
rect 10399 1550 10462 1572
rect 10399 185 10408 1550
rect 10399 114 10403 185
rect 10399 53 10408 114
rect 10460 53 10462 1550
rect 10399 30 10462 53
rect 10587 1550 10650 1572
rect 10587 179 10596 1550
rect 10587 104 10591 179
rect 10587 53 10596 104
rect 10648 53 10650 1550
rect 10587 30 10650 53
rect 10758 1550 10821 1572
rect 10758 1530 10767 1550
rect 10758 1457 10762 1530
rect 10758 53 10767 1457
rect 10819 53 10821 1550
rect 10758 30 10821 53
rect 10926 1550 10989 1572
rect 10926 173 10935 1550
rect 10926 98 10931 173
rect 10926 53 10935 98
rect 10987 53 10989 1550
rect 10926 30 10989 53
rect 11097 1550 11160 1572
rect 11097 1530 11106 1550
rect 11097 1457 11102 1530
rect 11097 53 11106 1457
rect 11158 53 11160 1550
rect 11097 30 11160 53
rect 11265 1550 11328 1572
rect 11265 176 11274 1550
rect 11265 101 11270 176
rect 11265 53 11274 101
rect 11326 53 11328 1550
rect 11265 30 11328 53
rect 11436 1550 11499 1572
rect 11436 1529 11445 1550
rect 11436 1456 11441 1529
rect 11436 53 11445 1456
rect 11497 53 11499 1550
rect 11436 30 11499 53
rect 11604 1550 11667 1572
rect 11604 182 11613 1550
rect 11604 107 11608 182
rect 11604 53 11613 107
rect 11665 53 11667 1550
rect 11604 30 11667 53
rect 11775 1550 11838 1572
rect 11775 1530 11784 1550
rect 11775 1457 11779 1530
rect 11775 53 11784 1457
rect 11836 53 11838 1550
rect 11775 30 11838 53
rect 11943 1550 12006 1572
rect 11943 181 11952 1550
rect 11943 106 11946 181
rect 11943 53 11952 106
rect 12004 53 12006 1550
rect 11943 30 12006 53
rect 12115 1550 12178 1572
rect 12115 1214 12124 1550
rect 12115 1141 12117 1214
rect 12115 53 12124 1141
rect 12176 53 12178 1550
rect 12115 30 12178 53
rect 12283 1550 12346 1572
rect 12283 182 12292 1550
rect 12283 107 12288 182
rect 12283 53 12292 107
rect 12344 53 12346 1550
rect 12283 30 12346 53
rect 12454 1550 12517 1572
rect 12454 1213 12463 1550
rect 12515 1213 12517 1550
rect 12454 1140 12459 1213
rect 12454 53 12463 1140
rect 12515 53 12517 1140
rect 12454 30 12517 53
rect 12622 1550 12685 1572
rect 12622 182 12631 1550
rect 12622 107 12626 182
rect 12622 53 12631 107
rect 12683 53 12685 1550
rect 12622 30 12685 53
rect 12793 1550 12856 1572
rect 12793 1210 12802 1550
rect 12793 1137 12796 1210
rect 12793 53 12802 1137
rect 12854 53 12856 1550
rect 12793 30 12856 53
rect 12961 1550 13024 1572
rect 12961 183 12970 1550
rect 12961 108 12964 183
rect 12961 53 12970 108
rect 13022 53 13024 1550
rect 12961 30 13024 53
rect 13132 1550 13195 1572
rect 13132 1212 13141 1550
rect 13132 1139 13133 1212
rect 13132 53 13141 1139
rect 13193 53 13195 1550
rect 13132 30 13195 53
rect 13300 1550 13363 1572
rect 13300 189 13309 1550
rect 13300 114 13304 189
rect 13300 53 13309 114
rect 13361 53 13363 1550
rect 13300 30 13363 53
rect 13486 1550 13549 1572
rect 13486 184 13495 1550
rect 13547 184 13549 1550
rect 13486 109 13492 184
rect 13548 109 13549 184
rect 13486 53 13495 109
rect 13547 53 13549 109
rect 13486 30 13549 53
rect 13658 1550 13721 1572
rect 13658 1533 13667 1550
rect 13658 1453 13661 1533
rect 13658 53 13667 1453
rect 13719 53 13721 1550
rect 13658 30 13721 53
rect 13826 1550 13889 1572
rect 13826 185 13835 1550
rect 13826 110 13830 185
rect 13826 53 13835 110
rect 13887 53 13889 1550
rect 13826 30 13889 53
rect 13997 1550 14060 1572
rect 13997 1537 14006 1550
rect 14058 1537 14060 1550
rect 13997 1457 14003 1537
rect 14059 1457 14060 1537
rect 13997 53 14006 1457
rect 14058 53 14060 1457
rect 13997 30 14060 53
rect 14165 1550 14228 1572
rect 14165 185 14174 1550
rect 14165 110 14170 185
rect 14165 53 14174 110
rect 14226 53 14228 1550
rect 14165 30 14228 53
rect 14336 1550 14399 1572
rect 14336 1209 14345 1550
rect 14397 1209 14399 1550
rect 14336 1136 14341 1209
rect 14336 53 14345 1136
rect 14397 53 14399 1136
rect 14336 30 14399 53
rect 14504 1550 14567 1572
rect 14504 187 14513 1550
rect 14504 112 14508 187
rect 14504 53 14513 112
rect 14565 53 14567 1550
rect 14504 30 14567 53
rect 14675 1550 14738 1572
rect 14675 1210 14684 1550
rect 14675 1137 14678 1210
rect 14675 53 14684 1137
rect 14736 53 14738 1550
rect 14675 30 14738 53
rect 14843 1550 14906 1572
rect 14843 190 14852 1550
rect 14843 115 14847 190
rect 14843 53 14852 115
rect 14904 53 14906 1550
rect 14843 30 14906 53
rect 15027 1550 15090 1572
rect 15027 192 15036 1550
rect 15088 192 15090 1550
rect 15027 117 15033 192
rect 15089 117 15090 192
rect 15027 53 15036 117
rect 15088 53 15090 117
rect 15027 30 15090 53
rect 15198 1550 15261 1572
rect 15198 1529 15207 1550
rect 15198 1459 15201 1529
rect 15198 53 15207 1459
rect 15259 53 15261 1550
rect 15198 30 15261 53
rect 15366 1550 15429 1572
rect 15366 198 15375 1550
rect 15366 123 15371 198
rect 15366 53 15375 123
rect 15427 53 15429 1550
rect 15366 30 15429 53
rect 15537 1550 15600 1572
rect 15537 1210 15546 1550
rect 15598 1210 15600 1550
rect 15537 1137 15541 1210
rect 15599 1137 15600 1210
rect 15537 53 15546 1137
rect 15598 53 15600 1137
rect 15537 30 15600 53
rect 15705 1550 15768 1572
rect 15705 204 15714 1550
rect 15705 129 15710 204
rect 15705 53 15714 129
rect 15766 53 15768 1550
rect 15705 30 15768 53
rect 15897 1550 15960 1572
rect 15897 1529 15906 1550
rect 15897 1457 15902 1529
rect 15897 53 15906 1457
rect 15958 53 15960 1550
rect 15897 30 15960 53
rect 16068 1550 16131 1572
rect 16068 200 16077 1550
rect 16068 136 16073 200
rect 16068 53 16077 136
rect 16129 53 16131 1550
rect 16068 30 16131 53
rect 16236 1550 16299 1572
rect 16236 1212 16245 1550
rect 16297 1212 16299 1550
rect 16236 1134 16242 1212
rect 16298 1134 16299 1212
rect 16236 53 16245 1134
rect 16297 53 16299 1134
rect 16236 30 16299 53
rect 16437 1545 16500 1572
rect 16437 1540 16446 1545
rect 16437 1459 16440 1540
rect 16437 53 16446 1459
rect 16498 53 16500 1545
rect 16437 30 16500 53
rect 16608 1545 16671 1572
rect 16608 222 16617 1545
rect 16608 143 16612 222
rect 16608 53 16617 143
rect 16669 53 16671 1545
rect 16608 30 16671 53
rect 16776 1545 16839 1572
rect 16776 1540 16785 1545
rect 16776 1459 16780 1540
rect 16776 53 16785 1459
rect 16837 53 16839 1545
rect 16776 30 16839 53
rect 16947 1545 17010 1572
rect 16947 215 16956 1545
rect 16947 136 16951 215
rect 16947 53 16956 136
rect 17008 53 17010 1545
rect 16947 30 17010 53
rect 17115 1545 17178 1572
rect 17115 1540 17124 1545
rect 17115 1459 17119 1540
rect 17115 53 17124 1459
rect 17176 53 17178 1545
rect 17115 30 17178 53
rect 17286 1545 17349 1572
rect 17286 224 17295 1545
rect 17286 152 17289 224
rect 17286 53 17295 152
rect 17347 53 17349 1545
rect 17286 30 17349 53
rect 17454 1545 17517 1572
rect 17454 1543 17463 1545
rect 17454 1462 17457 1543
rect 17454 53 17463 1462
rect 17515 53 17517 1545
rect 17454 30 17517 53
rect 17625 1545 17688 1572
rect 17625 223 17634 1545
rect 17686 223 17688 1545
rect 17816 1545 17879 1572
rect 17816 1543 17825 1545
rect 17816 1462 17819 1543
rect 17816 830 17825 1462
rect 17877 830 17879 1545
rect 17816 814 17879 830
rect 17987 1545 18050 1572
rect 17987 1367 17996 1545
rect 17987 1293 17991 1367
rect 17987 830 17996 1293
rect 18048 830 18050 1545
rect 18198 1545 18261 1572
rect 18198 1368 18207 1545
rect 18198 1303 18201 1368
rect 18198 1241 18207 1303
rect 18259 1241 18261 1545
rect 18198 1220 18261 1241
rect 18369 1545 18432 1572
rect 18369 1543 18378 1545
rect 18369 1460 18374 1543
rect 18369 1240 18378 1460
rect 18430 1240 18432 1545
rect 18369 1220 18432 1240
rect 18540 1545 18603 1572
rect 18540 1363 18549 1545
rect 18540 1293 18544 1363
rect 18540 1240 18549 1293
rect 18601 1240 18603 1545
rect 18540 1220 18603 1240
rect 18748 1545 18811 1572
rect 18748 1352 18757 1545
rect 18748 1270 18753 1352
rect 18748 1240 18757 1270
rect 18809 1240 18811 1545
rect 18748 1220 18811 1240
rect 18917 1545 18980 1572
rect 18917 1542 18926 1545
rect 18917 1457 18922 1542
rect 18917 1240 18926 1457
rect 18978 1240 18980 1545
rect 18917 1220 18980 1240
rect 19088 1545 19151 1572
rect 19088 1240 19097 1545
rect 19149 1240 19151 1545
rect 19088 1220 19151 1240
rect 19309 1545 19372 1572
rect 19309 1336 19318 1545
rect 19309 1251 19314 1336
rect 19309 1240 19318 1251
rect 19370 1240 19372 1545
rect 19309 1220 19372 1240
rect 19478 1545 19541 1572
rect 19478 1543 19487 1545
rect 19478 1471 19481 1543
rect 19478 1240 19487 1471
rect 19539 1240 19541 1545
rect 19478 1220 19541 1240
rect 19649 1545 19712 1572
rect 19649 1316 19658 1545
rect 19710 1316 19712 1545
rect 19649 1241 19655 1316
rect 19711 1241 19712 1316
rect 19649 1240 19658 1241
rect 19710 1240 19712 1241
rect 19649 1220 19712 1240
rect 19858 1545 19921 1572
rect 19858 1240 19867 1545
rect 19919 1240 19921 1545
rect 19858 1220 19921 1240
rect 20027 1552 20090 1572
rect 20027 1480 20031 1552
rect 20087 1545 20090 1552
rect 20027 1240 20036 1480
rect 20088 1240 20090 1545
rect 20027 1220 20090 1240
rect 20198 1545 20261 1572
rect 20198 1240 20207 1545
rect 20259 1543 20261 1545
rect 20698 1543 20708 1654
rect 20259 1526 20708 1543
rect 20259 1438 20699 1526
rect 20259 1432 20708 1438
rect 20259 1240 20261 1432
rect 20198 1220 20261 1240
rect 19089 1110 19150 1220
rect 18121 1106 19150 1110
rect 17987 814 18050 830
rect 18118 1052 19150 1106
rect 18118 1050 18387 1052
rect 19089 1050 19150 1052
rect 19858 1099 19920 1220
rect 20698 1188 20708 1432
rect 20760 1188 20771 1654
rect 20698 1139 20771 1188
rect 20863 1655 20936 1717
rect 20863 1265 20875 1655
rect 20927 1265 20936 1655
rect 20863 1189 20869 1265
rect 20929 1189 20936 1265
rect 20863 1143 20936 1189
rect 21427 1156 21469 1717
rect 21563 1156 21584 1717
rect 20253 1101 20402 1121
rect 20253 1099 20292 1101
rect 17625 153 17626 223
rect 18118 204 18177 1050
rect 19858 1032 20292 1099
rect 20378 1032 20402 1101
rect 19858 1029 20402 1032
rect 20253 1003 20402 1029
rect 18343 943 18466 974
rect 18534 970 18640 971
rect 18343 874 18377 943
rect 18440 874 18466 943
rect 18343 840 18466 874
rect 18533 936 18640 970
rect 18533 867 18552 936
rect 18615 867 18640 936
rect 18533 838 18640 867
rect 18534 835 18640 838
rect 18883 935 18968 969
rect 18883 866 18893 935
rect 18956 866 18968 935
rect 18883 837 18968 866
rect 19039 936 19133 970
rect 19039 867 19058 936
rect 19121 867 19133 936
rect 19039 838 19133 867
rect 19402 935 19487 969
rect 19402 866 19412 935
rect 19475 866 19487 935
rect 19402 837 19487 866
rect 19558 936 19652 970
rect 19558 867 19577 936
rect 19640 867 19652 936
rect 19558 838 19652 867
rect 19922 935 20007 969
rect 19922 866 19932 935
rect 19995 866 20007 935
rect 19922 837 20007 866
rect 20078 936 20172 970
rect 20078 867 20097 936
rect 20160 867 20172 936
rect 20078 838 20172 867
rect 20454 935 20539 969
rect 20454 866 20464 935
rect 20527 866 20539 935
rect 20454 837 20539 866
rect 20610 936 20704 970
rect 20610 867 20629 936
rect 20692 867 20704 936
rect 20610 838 20704 867
rect 20972 935 21057 969
rect 20972 866 20982 935
rect 21045 866 21057 935
rect 20972 837 21057 866
rect 21128 936 21222 970
rect 21128 867 21147 936
rect 21210 867 21222 936
rect 21128 838 21222 867
rect 17625 53 17634 153
rect 17686 53 17688 153
rect 18055 188 18177 204
rect 18055 131 18079 188
rect 18148 131 18177 188
rect 18055 116 18177 131
rect 18285 734 18348 761
rect 18285 702 18294 734
rect 18285 635 18287 702
rect 18055 115 18150 116
rect 17625 30 17688 53
rect 18285 19 18294 635
rect 18346 19 18348 734
rect 18285 3 18348 19
rect 18456 734 18519 761
rect 18456 131 18465 734
rect 18517 131 18519 734
rect 18456 35 18462 131
rect 18456 19 18465 35
rect 18517 19 18519 35
rect 18456 3 18519 19
rect 18627 734 18690 761
rect 18627 523 18636 734
rect 18688 700 18690 734
rect 18799 734 18862 761
rect 18799 706 18808 734
rect 18688 633 18691 700
rect 18799 635 18804 706
rect 18860 700 18862 734
rect 18968 734 19031 761
rect 18627 447 18630 523
rect 18627 19 18636 447
rect 18688 19 18690 633
rect 18627 3 18690 19
rect 18799 19 18808 635
rect 18860 633 18863 700
rect 18860 19 18862 633
rect 18799 3 18862 19
rect 18968 126 18977 734
rect 18968 30 18972 126
rect 18968 19 18977 30
rect 19029 19 19031 734
rect 18968 3 19031 19
rect 19139 734 19202 761
rect 19139 518 19148 734
rect 19200 700 19202 734
rect 19318 734 19381 761
rect 19318 718 19327 734
rect 19317 706 19326 718
rect 19200 633 19203 700
rect 19317 635 19322 706
rect 19379 700 19381 734
rect 19487 734 19550 761
rect 19139 442 19142 518
rect 19139 19 19148 442
rect 19200 19 19202 633
rect 19317 624 19326 635
rect 19379 633 19382 700
rect 19139 3 19202 19
rect 19318 19 19327 624
rect 19379 19 19381 633
rect 19318 3 19381 19
rect 19487 130 19496 734
rect 19487 34 19490 130
rect 19487 19 19496 34
rect 19548 19 19550 734
rect 19658 734 19721 761
rect 19658 530 19667 734
rect 19719 700 19721 734
rect 19838 734 19901 761
rect 19838 717 19847 734
rect 19837 705 19846 717
rect 19719 633 19722 700
rect 19837 634 19842 705
rect 19899 700 19901 734
rect 20007 734 20070 761
rect 19656 516 19665 530
rect 19656 440 19659 516
rect 19656 430 19665 440
rect 19487 3 19550 19
rect 19658 19 19667 430
rect 19719 19 19721 633
rect 19837 623 19846 634
rect 19899 632 19902 700
rect 19658 3 19721 19
rect 19838 19 19847 623
rect 19899 19 19901 632
rect 19838 3 19901 19
rect 20007 132 20016 734
rect 20007 36 20009 132
rect 20007 19 20016 36
rect 20068 19 20070 734
rect 20178 734 20241 761
rect 20178 530 20187 734
rect 20239 700 20241 734
rect 20370 734 20433 761
rect 20370 729 20379 734
rect 20365 717 20374 729
rect 20239 633 20242 700
rect 20365 646 20370 717
rect 20431 700 20433 734
rect 20539 734 20602 761
rect 20365 635 20374 646
rect 20175 516 20184 530
rect 20175 440 20178 516
rect 20175 430 20184 440
rect 20007 3 20070 19
rect 20178 19 20187 430
rect 20239 19 20241 633
rect 20178 3 20241 19
rect 20370 19 20379 635
rect 20431 633 20434 700
rect 20431 19 20433 633
rect 20370 3 20433 19
rect 20539 134 20548 734
rect 20539 38 20543 134
rect 20539 19 20548 38
rect 20600 19 20602 734
rect 20710 734 20773 761
rect 20710 530 20719 734
rect 20771 700 20773 734
rect 20888 734 20951 761
rect 20888 724 20897 734
rect 20884 712 20893 724
rect 20771 633 20774 700
rect 20884 641 20889 712
rect 20949 700 20951 734
rect 21057 734 21120 761
rect 20706 516 20715 530
rect 20706 440 20709 516
rect 20706 430 20715 440
rect 20539 3 20602 19
rect 20710 19 20719 430
rect 20771 19 20773 633
rect 20884 630 20893 641
rect 20949 633 20952 700
rect 20710 3 20773 19
rect 20888 19 20897 630
rect 20949 19 20951 633
rect 20888 3 20951 19
rect 21057 130 21066 734
rect 21057 34 21061 130
rect 21057 19 21066 34
rect 21118 19 21120 734
rect 21228 734 21291 761
rect 21228 530 21237 734
rect 21289 700 21291 734
rect 21289 633 21292 700
rect 21223 516 21232 530
rect 21223 440 21226 516
rect 21223 430 21232 440
rect 21057 3 21120 19
rect 21228 19 21237 430
rect 21289 19 21291 633
rect 21228 3 21291 19
rect 21427 538 21584 1156
rect 1799 -148 1919 -3
rect 21427 -23 21462 538
rect 21556 -23 21584 538
rect 1799 -149 17252 -148
rect 18821 -149 20526 -147
rect 21427 -149 21584 -23
rect 1799 -161 21584 -149
rect 1799 -165 7595 -161
rect 1799 -168 3667 -165
rect 1799 -262 2224 -168
rect 2785 -259 3667 -168
rect 4228 -172 6375 -165
rect 4228 -259 5075 -172
rect 2785 -262 5075 -259
rect 1799 -266 5075 -262
rect 5636 -259 6375 -172
rect 6936 -255 7595 -165
rect 8156 -162 21584 -161
rect 8156 -165 18628 -162
rect 8156 -168 13452 -165
rect 8156 -255 9024 -168
rect 6936 -259 9024 -255
rect 5636 -262 9024 -259
rect 9585 -262 10334 -168
rect 10895 -262 11982 -168
rect 12543 -259 13452 -168
rect 14013 -259 15071 -165
rect 15632 -169 18628 -165
rect 15632 -259 16873 -169
rect 12543 -262 16873 -259
rect 5636 -263 16873 -262
rect 17434 -256 18628 -169
rect 19189 -165 21584 -162
rect 19189 -256 20208 -165
rect 17434 -259 20208 -256
rect 20769 -259 21584 -165
rect 17434 -263 21584 -259
rect 5636 -266 21584 -263
rect 1799 -279 21584 -266
rect 1799 -280 1919 -279
rect -10893 -281 1690 -280
rect 4844 -281 21584 -279
rect 17245 -282 21435 -281
rect -9502 -460 -9145 -459
rect -9502 -461 6533 -460
rect -9502 -466 19531 -461
rect -9502 -471 21775 -466
rect -9502 -576 -9478 -471
rect -9397 -486 21775 -471
rect -9397 -562 6946 -486
rect 7026 -495 21775 -486
rect 7026 -562 16742 -495
rect -9397 -571 16742 -562
rect 16828 -571 21775 -495
rect -9397 -576 21775 -571
rect -9502 -588 21775 -576
rect 6458 -589 21775 -588
rect -3860 -684 21775 -670
rect -3860 -774 -3839 -684
rect -3775 -704 21775 -684
rect -3775 -767 11915 -704
rect 12004 -705 21775 -704
rect 12004 -767 17270 -705
rect -3775 -774 17270 -767
rect -3860 -775 17270 -774
rect 17332 -775 21775 -705
rect -3860 -793 21775 -775
rect -1801 -915 21775 -900
rect -1801 -1001 -1789 -915
rect -1710 -924 21775 -915
rect -1710 -987 14005 -924
rect 14067 -987 21775 -924
rect -1710 -1001 21775 -987
rect -1801 -1011 21775 -1001
rect -1006 -1148 21775 -1138
rect -1009 -1158 21775 -1148
rect -1009 -1162 15766 -1158
rect -1009 -1241 -996 -1162
rect -924 -1165 15766 -1162
rect -924 -1227 15318 -1165
rect 15378 -1227 15766 -1165
rect -924 -1241 15766 -1227
rect -1009 -1246 15766 -1241
rect 15855 -1246 21775 -1158
rect -1009 -1255 21775 -1246
rect -1006 -1258 21775 -1255
rect -485 -1406 21775 -1385
rect -485 -1488 -469 -1406
rect -399 -1488 16058 -1406
rect -485 -1489 16058 -1488
rect 16128 -1489 21775 -1406
rect -485 -1509 21775 -1489
rect -106 -1642 21775 -1627
rect -106 -1653 18451 -1642
rect -106 -1654 17775 -1653
rect -106 -1728 -92 -1654
rect -22 -1728 17775 -1654
rect -106 -1735 17775 -1728
rect 17836 -1730 18451 -1653
rect 18527 -1730 21775 -1642
rect 17836 -1735 21775 -1730
rect -106 -1753 21775 -1735
rect -106 -1754 725 -1753
rect 222 -1875 958 -1871
rect 220 -1899 21775 -1875
rect 220 -1909 18964 -1899
rect 220 -1984 241 -1909
rect 311 -1973 18964 -1909
rect 19026 -1973 21775 -1899
rect 311 -1984 21775 -1973
rect 220 -2000 21775 -1984
rect 450 -2116 967 -2113
rect 450 -2136 21775 -2116
rect 450 -2226 471 -2136
rect 538 -2140 21775 -2136
rect 538 -2141 19490 -2140
rect 538 -2224 18066 -2141
rect 18137 -2224 19490 -2141
rect 538 -2226 19490 -2224
rect 450 -2231 19490 -2226
rect 19561 -2231 21775 -2140
rect 450 -2245 21775 -2231
rect 771 -2372 21775 -2370
rect 770 -2400 21775 -2372
rect 770 -2403 20014 -2400
rect 770 -2484 783 -2403
rect 861 -2484 20014 -2403
rect 770 -2491 20014 -2484
rect 20085 -2491 21775 -2400
rect 770 -2499 21775 -2491
rect 1011 -2624 1962 -2622
rect 1010 -2635 21775 -2624
rect 1010 -2655 20548 -2635
rect 1010 -2735 1024 -2655
rect 1098 -2726 20548 -2655
rect 20619 -2726 21775 -2635
rect 1098 -2735 21775 -2726
rect 1010 -2752 21775 -2735
rect 1011 -2754 1962 -2752
rect 1348 -2900 1940 -2898
rect 1348 -2923 21775 -2900
rect 1348 -2929 21050 -2923
rect 1348 -3008 1365 -2929
rect 1443 -3008 21050 -2929
rect 1348 -3014 21050 -3008
rect 21121 -3014 21775 -2923
rect 1348 -3031 21775 -3014
rect 2989 -3212 21776 -3176
rect 2989 -3291 3009 -3212
rect 3096 -3291 21776 -3212
rect 2989 -3310 21776 -3291
<< via2 >>
rect -7618 1703 -7557 1767
rect -3629 1706 -3568 1770
rect -1901 1704 -1840 1768
rect -945 1700 -884 1764
rect -451 1693 -390 1757
rect -22 1678 39 1742
rect 191 1678 252 1742
rect 529 1679 590 1743
rect 744 1678 805 1742
rect 1099 1676 1160 1740
rect 1312 1678 1373 1742
rect -10565 1399 -10561 1465
rect -10561 1399 -10509 1465
rect -10396 138 -10394 222
rect -10394 138 -10341 222
rect -10341 138 -10340 222
rect -10236 1403 -10230 1469
rect -10230 1403 -10180 1469
rect -9905 1402 -9899 1468
rect -9899 1402 -9849 1468
rect -10063 138 -10008 222
rect -10008 138 -10007 222
rect -9734 137 -9679 221
rect -9679 137 -9678 221
rect -9573 1399 -9568 1465
rect -9568 1399 -9517 1465
rect -9403 136 -9348 220
rect -9348 136 -9347 220
rect -9238 1402 -9235 1468
rect -9235 1402 -9183 1468
rect -9183 1402 -9182 1468
rect -9070 139 -9015 223
rect -9015 139 -9014 223
rect -8907 1399 -8904 1465
rect -8904 1399 -8852 1465
rect -8852 1399 -8851 1465
rect -8739 139 -8684 223
rect -8684 139 -8683 223
rect -8577 1400 -8573 1466
rect -8573 1400 -8521 1466
rect -8408 141 -8353 225
rect -8353 141 -8352 225
rect -8246 1401 -8242 1467
rect -8242 1401 -8190 1467
rect -7915 1401 -7910 1467
rect -7910 1401 -7859 1467
rect -8076 143 -8021 227
rect -8021 143 -8020 227
rect -7745 143 -7690 227
rect -7690 143 -7689 227
rect -7584 1400 -7579 1466
rect -7579 1400 -7528 1466
rect -7253 1399 -7248 1465
rect -7248 1399 -7197 1465
rect -7413 143 -7358 227
rect -7358 143 -7357 227
rect -6921 1396 -6917 1462
rect -6917 1396 -6865 1462
rect -7082 143 -7027 227
rect -7027 143 -7026 227
rect -6752 143 -6697 227
rect -6697 143 -6696 227
rect -6589 1397 -6584 1463
rect -6584 1397 -6533 1463
rect -6419 143 -6364 227
rect -6364 143 -6363 227
rect -6256 1396 -6253 1462
rect -6253 1396 -6201 1462
rect -6201 1396 -6200 1462
rect -6088 143 -6033 227
rect -6033 143 -6032 227
rect -5926 1398 -5922 1464
rect -5922 1398 -5870 1464
rect -5595 1396 -5591 1462
rect -5591 1396 -5539 1462
rect -5755 153 -5700 237
rect -5700 153 -5699 237
rect -5426 153 -5371 237
rect -5371 153 -5370 237
rect -5263 1396 -5258 1462
rect -5258 1396 -5207 1462
rect -5094 161 -5091 240
rect -5091 161 -5038 240
rect -5038 161 -5037 240
rect -4932 1396 -4927 1462
rect -4927 1396 -4876 1462
rect -4602 1397 -4596 1463
rect -4596 1397 -4546 1463
rect -4761 161 -4760 240
rect -4760 161 -4705 240
rect -4705 161 -4704 240
rect -4271 1396 -4265 1462
rect -4265 1396 -4215 1462
rect -4431 161 -4430 240
rect -4430 161 -4375 240
rect -4375 161 -4374 240
rect -4101 161 -4100 240
rect -4100 161 -4045 240
rect -4045 161 -4044 240
rect -3936 1397 -3932 1463
rect -3932 1397 -3880 1463
rect -3606 1398 -3601 1464
rect -3601 1398 -3550 1464
rect -3767 161 -3766 240
rect -3766 161 -3711 240
rect -3711 161 -3710 240
rect -3275 1397 -3270 1463
rect -3270 1397 -3219 1463
rect -3436 161 -3435 240
rect -3435 161 -3380 240
rect -3380 161 -3379 240
rect -3106 160 -3105 239
rect -3105 160 -3050 239
rect -3050 160 -3049 239
rect -2944 1398 -2939 1464
rect -2939 1398 -2888 1464
rect -2775 161 -2774 240
rect -2774 161 -2719 240
rect -2719 161 -2718 240
rect -2614 1399 -2609 1465
rect -2609 1399 -2558 1465
rect -2282 1398 -2278 1464
rect -2278 1398 -2226 1464
rect -2444 161 -2443 240
rect -2443 161 -2388 240
rect -2388 161 -2387 240
rect -1953 1397 -1947 1463
rect -1947 1397 -1897 1463
rect -2113 161 -2112 240
rect -2112 161 -2057 240
rect -2057 161 -2056 240
rect -1783 161 -1782 240
rect -1782 161 -1727 240
rect -1727 161 -1726 240
rect -1621 1398 -1616 1464
rect -1616 1398 -1565 1464
rect -1289 1397 -1284 1463
rect -1284 1397 -1233 1463
rect -1451 161 -1450 240
rect -1450 161 -1395 240
rect -1395 161 -1394 240
rect -1120 161 -1119 240
rect -1119 161 -1064 240
rect -1064 161 -1063 240
rect -957 1399 -953 1465
rect -953 1399 -901 1465
rect -626 1401 -622 1467
rect -622 1401 -570 1467
rect -788 161 -787 240
rect -787 161 -732 240
rect -732 161 -731 240
rect -290 1402 -289 1468
rect -289 1402 -236 1468
rect -236 1402 -233 1468
rect -457 161 -456 240
rect -456 161 -401 240
rect -401 161 -400 240
rect -86 161 -85 240
rect -85 161 -29 240
rect 83 1395 87 1451
rect 87 1395 140 1451
rect 140 1395 142 1451
rect 250 161 251 240
rect 251 161 307 240
rect 466 161 467 240
rect 467 161 523 240
rect 637 1396 640 1452
rect 640 1396 693 1452
rect 693 1396 696 1452
rect 805 158 806 244
rect 806 158 859 244
rect 859 158 862 244
rect 1206 1396 1209 1452
rect 1209 1396 1262 1452
rect 1262 1396 1265 1452
rect 1040 159 1041 245
rect 1041 159 1094 245
rect 1094 159 1097 245
rect 1374 159 1375 245
rect 1375 159 1428 245
rect 1428 159 1431 245
rect 3258 1712 3370 1782
rect 6433 1712 6545 1782
rect 8886 1711 8998 1781
rect 11212 1714 11324 1784
rect 20781 1798 20865 1857
rect 12628 1710 12740 1780
rect 13857 1709 13969 1779
rect 14545 1709 14657 1779
rect 15176 1709 15288 1779
rect 15514 1709 15626 1779
rect 15943 1689 16027 1748
rect 16166 1689 16250 1748
rect 16751 1750 16870 1752
rect 16751 1696 16752 1750
rect 16752 1696 16870 1750
rect 16751 1695 16870 1696
rect 2061 1457 2067 1531
rect 2067 1457 2118 1531
rect 2230 80 2239 170
rect 2239 80 2290 170
rect 2401 1455 2407 1529
rect 2407 1455 2458 1529
rect 2570 80 2578 170
rect 2578 80 2630 170
rect 2741 1457 2746 1531
rect 2746 1457 2798 1531
rect 2910 80 2917 170
rect 2917 80 2969 170
rect 2969 80 2970 170
rect 3080 1460 3085 1534
rect 3085 1460 3137 1534
rect 3250 80 3256 170
rect 3256 80 3308 170
rect 3308 80 3310 170
rect 3420 1457 3424 1531
rect 3424 1457 3476 1531
rect 3476 1457 3477 1531
rect 3590 80 3596 170
rect 3596 80 3648 170
rect 3648 80 3650 170
rect 3759 1458 3764 1532
rect 3764 1458 3816 1532
rect 3928 80 3935 178
rect 3935 80 3987 178
rect 3987 80 3988 178
rect 4096 1458 4103 1532
rect 4103 1458 4153 1532
rect 4267 78 4274 168
rect 4274 78 4326 168
rect 4326 78 4327 168
rect 4435 1461 4442 1535
rect 4442 1461 4492 1535
rect 4606 82 4613 172
rect 4613 82 4665 172
rect 4665 82 4666 172
rect 4773 1461 4781 1535
rect 4781 1461 4830 1535
rect 4976 108 4981 179
rect 4981 108 5032 179
rect 5148 1458 5153 1530
rect 5153 1458 5204 1530
rect 5314 107 5321 178
rect 5321 107 5370 178
rect 5487 1458 5492 1530
rect 5492 1458 5543 1530
rect 5654 106 5660 177
rect 5660 106 5710 177
rect 5826 1458 5831 1530
rect 5831 1458 5882 1530
rect 5994 106 5999 177
rect 5999 106 6050 177
rect 6167 1458 6170 1530
rect 6170 1458 6222 1530
rect 6222 1458 6223 1530
rect 6333 104 6338 175
rect 6338 104 6389 175
rect 6504 1456 6510 1528
rect 6510 1456 6560 1528
rect 6673 104 6678 175
rect 6678 104 6729 175
rect 6844 1456 6849 1528
rect 6849 1456 6900 1528
rect 7012 103 7017 174
rect 7017 103 7068 174
rect 7183 1457 7188 1529
rect 7188 1457 7239 1529
rect 7351 104 7356 175
rect 7356 104 7407 175
rect 7523 1457 7527 1529
rect 7527 1457 7579 1529
rect 7690 103 7695 174
rect 7695 103 7746 174
rect 7861 1137 7866 1210
rect 7866 1137 7918 1210
rect 7918 1137 7919 1210
rect 8028 104 8034 175
rect 8034 104 8084 175
rect 8201 1137 8205 1210
rect 8205 1137 8257 1210
rect 8257 1137 8259 1210
rect 8366 103 8373 174
rect 8373 103 8422 174
rect 8539 1136 8544 1209
rect 8544 1136 8596 1209
rect 8596 1136 8597 1209
rect 8706 111 8712 182
rect 8712 111 8762 182
rect 8879 1140 8883 1213
rect 8883 1140 8935 1213
rect 8935 1140 8937 1213
rect 9047 118 9051 189
rect 9051 118 9103 189
rect 9217 1141 9223 1214
rect 9223 1141 9275 1214
rect 9386 112 9391 183
rect 9391 112 9442 183
rect 9555 1141 9562 1214
rect 9562 1141 9613 1214
rect 9726 116 9730 187
rect 9730 116 9782 187
rect 9894 1141 9901 1214
rect 9901 1141 9952 1214
rect 10065 115 10069 186
rect 10069 115 10121 186
rect 10234 1140 10240 1213
rect 10240 1140 10292 1213
rect 10403 114 10408 185
rect 10408 114 10459 185
rect 10591 104 10596 179
rect 10596 104 10647 179
rect 10762 1457 10767 1530
rect 10767 1457 10818 1530
rect 10931 98 10935 173
rect 10935 98 10987 173
rect 11102 1457 11106 1530
rect 11106 1457 11158 1530
rect 11270 101 11274 176
rect 11274 101 11326 176
rect 11441 1456 11445 1529
rect 11445 1456 11497 1529
rect 11608 107 11613 182
rect 11613 107 11664 182
rect 11779 1457 11784 1530
rect 11784 1457 11835 1530
rect 11946 106 11952 181
rect 11952 106 12002 181
rect 12117 1141 12124 1214
rect 12124 1141 12175 1214
rect 12288 107 12292 182
rect 12292 107 12344 182
rect 12459 1140 12463 1213
rect 12463 1140 12515 1213
rect 12515 1140 12517 1213
rect 12626 107 12631 182
rect 12631 107 12682 182
rect 12796 1137 12802 1210
rect 12802 1137 12854 1210
rect 12964 108 12970 183
rect 12970 108 13020 183
rect 13133 1139 13141 1212
rect 13141 1139 13191 1212
rect 13304 114 13309 189
rect 13309 114 13360 189
rect 13492 109 13495 184
rect 13495 109 13547 184
rect 13547 109 13548 184
rect 13661 1453 13667 1533
rect 13667 1453 13717 1533
rect 13830 110 13835 185
rect 13835 110 13886 185
rect 14003 1457 14006 1537
rect 14006 1457 14058 1537
rect 14058 1457 14059 1537
rect 14170 110 14174 185
rect 14174 110 14226 185
rect 14341 1136 14345 1209
rect 14345 1136 14397 1209
rect 14397 1136 14399 1209
rect 14508 112 14513 187
rect 14513 112 14564 187
rect 14678 1137 14684 1210
rect 14684 1137 14736 1210
rect 14847 115 14852 190
rect 14852 115 14903 190
rect 15033 117 15036 192
rect 15036 117 15088 192
rect 15088 117 15089 192
rect 15201 1459 15207 1529
rect 15207 1459 15257 1529
rect 15371 123 15375 198
rect 15375 123 15427 198
rect 15541 1137 15546 1210
rect 15546 1137 15598 1210
rect 15598 1137 15599 1210
rect 15710 129 15714 204
rect 15714 129 15766 204
rect 15902 1457 15906 1529
rect 15906 1457 15958 1529
rect 16073 136 16077 200
rect 16077 136 16129 200
rect 16242 1134 16245 1212
rect 16245 1134 16297 1212
rect 16297 1134 16298 1212
rect 16440 1459 16446 1540
rect 16446 1459 16496 1540
rect 16612 143 16617 222
rect 16617 143 16668 222
rect 16780 1459 16785 1540
rect 16785 1459 16836 1540
rect 16951 136 16956 215
rect 16956 136 17007 215
rect 17119 1459 17124 1540
rect 17124 1459 17175 1540
rect 17289 152 17295 224
rect 17295 152 17345 224
rect 17457 1462 17463 1543
rect 17463 1462 17513 1543
rect 17819 1462 17825 1543
rect 17825 1462 17875 1543
rect 17991 1293 17996 1367
rect 17996 1293 18048 1367
rect 18201 1303 18207 1368
rect 18207 1303 18259 1368
rect 18374 1460 18378 1543
rect 18378 1460 18430 1543
rect 18544 1293 18549 1363
rect 18549 1293 18600 1363
rect 18753 1270 18757 1352
rect 18757 1270 18809 1352
rect 18922 1457 18926 1542
rect 18926 1457 18978 1542
rect 19314 1251 19318 1336
rect 19318 1251 19370 1336
rect 19481 1471 19487 1543
rect 19487 1471 19537 1543
rect 19655 1241 19658 1316
rect 19658 1241 19710 1316
rect 19710 1241 19711 1316
rect 20031 1545 20087 1552
rect 20031 1480 20036 1545
rect 20036 1480 20087 1545
rect 20699 1438 20708 1526
rect 20708 1438 20756 1526
rect 20869 1189 20875 1265
rect 20875 1189 20927 1265
rect 20927 1189 20929 1265
rect 17626 153 17634 223
rect 17634 153 17686 223
rect 17686 153 17688 223
rect 20292 1032 20378 1101
rect 18377 874 18440 943
rect 18552 867 18615 936
rect 18893 866 18956 935
rect 19058 867 19121 936
rect 19412 866 19475 935
rect 19577 867 19640 936
rect 19932 866 19995 935
rect 20097 867 20160 936
rect 20464 866 20527 935
rect 20629 867 20692 936
rect 20982 866 21045 935
rect 21147 867 21210 936
rect 18079 131 18148 188
rect 18287 635 18294 702
rect 18294 635 18346 702
rect 18462 35 18465 131
rect 18465 35 18517 131
rect 18517 35 18519 131
rect 18804 635 18808 706
rect 18808 635 18860 706
rect 18630 447 18636 523
rect 18636 447 18686 523
rect 18972 30 18977 126
rect 18977 30 19029 126
rect 19322 635 19326 706
rect 19326 635 19378 706
rect 19142 442 19148 518
rect 19148 442 19198 518
rect 19490 34 19496 130
rect 19496 34 19547 130
rect 19842 634 19846 705
rect 19846 634 19898 705
rect 19659 440 19665 516
rect 19665 440 19715 516
rect 20009 36 20016 132
rect 20016 36 20066 132
rect 20370 646 20374 717
rect 20374 646 20426 717
rect 20178 440 20184 516
rect 20184 440 20234 516
rect 20543 38 20548 134
rect 20548 38 20600 134
rect 20889 641 20893 712
rect 20893 641 20945 712
rect 20709 440 20715 516
rect 20715 440 20765 516
rect 21061 34 21066 130
rect 21066 34 21118 130
rect 21226 440 21232 516
rect 21232 440 21282 516
rect -9478 -576 -9397 -471
rect 6946 -562 7026 -486
rect 16742 -571 16828 -495
rect -3839 -774 -3775 -684
rect 11915 -767 12004 -704
rect 17270 -775 17332 -705
rect -1789 -1001 -1710 -915
rect 14005 -987 14067 -924
rect -996 -1241 -924 -1162
rect 15318 -1227 15378 -1165
rect 15766 -1246 15855 -1158
rect -469 -1488 -399 -1406
rect 16058 -1489 16128 -1406
rect -92 -1728 -22 -1654
rect 17775 -1735 17836 -1653
rect 18451 -1730 18527 -1642
rect 241 -1984 311 -1909
rect 18964 -1973 19026 -1899
rect 471 -2226 538 -2136
rect 18066 -2224 18137 -2141
rect 19490 -2231 19561 -2140
rect 783 -2484 861 -2403
rect 20014 -2491 20085 -2400
rect 1024 -2735 1098 -2655
rect 20548 -2726 20619 -2635
rect 1365 -3008 1443 -2929
rect 21050 -3014 21121 -2923
rect 3009 -3291 3096 -3212
<< metal3 >>
rect -7644 1793 -7535 2411
rect -7645 1767 -7535 1793
rect -7645 1703 -7618 1767
rect -7557 1703 -7535 1767
rect -7645 1674 -7535 1703
rect -3656 1770 -3547 2417
rect -3656 1706 -3629 1770
rect -3568 1706 -3547 1770
rect -3656 1678 -3547 1706
rect -1931 1794 -1822 2412
rect -1931 1768 -1821 1794
rect -971 1790 -862 2410
rect -1931 1704 -1901 1768
rect -1840 1704 -1821 1768
rect -3656 1677 -3549 1678
rect -7644 1672 -7535 1674
rect -1931 1675 -1821 1704
rect -972 1764 -862 1790
rect -972 1700 -945 1764
rect -884 1700 -862 1764
rect -1931 1673 -1822 1675
rect -972 1671 -862 1700
rect -478 1783 -370 2409
rect -478 1757 -369 1783
rect -478 1693 -451 1757
rect -390 1693 -369 1757
rect -478 1665 -369 1693
rect -48 1742 60 2410
rect -48 1678 -22 1742
rect 39 1678 60 1742
rect -478 1664 -370 1665
rect -48 1650 60 1678
rect 165 1742 273 2410
rect 165 1678 191 1742
rect 252 1678 273 1742
rect 165 1650 273 1678
rect 503 1743 611 2411
rect 503 1679 529 1743
rect 590 1679 611 1743
rect 503 1651 611 1679
rect 719 1742 827 2410
rect 719 1678 744 1742
rect 805 1678 827 1742
rect 719 1650 827 1678
rect 1074 1740 1182 2407
rect 1074 1676 1099 1740
rect 1160 1676 1182 1740
rect 1074 1648 1182 1676
rect 1287 1742 1395 2410
rect 3240 1801 3379 2411
rect 6415 1801 6554 2411
rect 1287 1678 1312 1742
rect 1373 1678 1395 1742
rect 3221 1782 3399 1801
rect 3221 1712 3258 1782
rect 3370 1712 3399 1782
rect 3221 1690 3399 1712
rect 6396 1782 6574 1801
rect 8868 1800 9007 2410
rect 11194 1803 11333 2413
rect 6396 1712 6433 1782
rect 6545 1712 6574 1782
rect 6396 1690 6574 1712
rect 8849 1781 9027 1800
rect 8849 1711 8886 1781
rect 8998 1711 9027 1781
rect 8849 1689 9027 1711
rect 11175 1784 11353 1803
rect 12610 1799 12749 2409
rect 11175 1714 11212 1784
rect 11324 1714 11353 1784
rect 11175 1692 11353 1714
rect 12591 1780 12769 1799
rect 13839 1798 13978 2408
rect 14527 1798 14666 2408
rect 15158 1798 15297 2408
rect 15496 1798 15635 2408
rect 12591 1710 12628 1780
rect 12740 1710 12769 1780
rect 12591 1688 12769 1710
rect 13820 1779 13998 1798
rect 13820 1709 13857 1779
rect 13969 1709 13998 1779
rect 13820 1687 13998 1709
rect 14508 1779 14686 1798
rect 14508 1709 14545 1779
rect 14657 1709 14686 1779
rect 14508 1687 14686 1709
rect 15140 1779 15317 1798
rect 15140 1709 15176 1779
rect 15288 1709 15317 1779
rect 15140 1688 15317 1709
rect 15478 1779 15655 1798
rect 15478 1709 15514 1779
rect 15626 1709 15655 1779
rect 15478 1688 15655 1709
rect 15930 1763 16042 2417
rect 15930 1748 16043 1763
rect 15930 1689 15943 1748
rect 16027 1689 16043 1748
rect 1287 1650 1395 1678
rect 15930 1670 16043 1689
rect 16153 1748 16265 2417
rect 16153 1689 16166 1748
rect 16250 1689 16265 1748
rect 16153 1670 16265 1689
rect 16726 1767 16876 2431
rect 20766 1872 20878 2429
rect 20766 1857 20880 1872
rect 20766 1798 20781 1857
rect 20865 1798 20880 1857
rect 20766 1781 20880 1798
rect 16726 1752 16886 1767
rect 16726 1695 16751 1752
rect 16870 1695 16886 1752
rect 16726 1678 16886 1695
rect 19162 1552 19473 1553
rect 16421 1551 17707 1552
rect 17789 1551 18069 1552
rect 18171 1551 20031 1552
rect 16419 1543 20031 1551
rect 4750 1540 7614 1541
rect 16419 1540 17457 1543
rect 4750 1539 12114 1540
rect 13460 1539 13657 1540
rect 4750 1538 16320 1539
rect 1920 1537 16320 1538
rect 1920 1535 14003 1537
rect 1920 1534 4435 1535
rect 1920 1531 3080 1534
rect -11165 1469 547 1475
rect -11165 1465 -10236 1469
rect -11165 1399 -10565 1465
rect -10509 1403 -10236 1465
rect -10180 1468 547 1469
rect -10180 1403 -9905 1468
rect -10509 1402 -9905 1403
rect -9849 1465 -9238 1468
rect -9849 1402 -9573 1465
rect -10509 1399 -9573 1402
rect -9517 1402 -9238 1465
rect -9182 1467 -290 1468
rect -9182 1466 -8246 1467
rect -9182 1465 -8577 1466
rect -9182 1402 -8907 1465
rect -9517 1399 -8907 1402
rect -8851 1400 -8577 1465
rect -8521 1401 -8246 1466
rect -8190 1401 -7915 1467
rect -7859 1466 -626 1467
rect -7859 1401 -7584 1466
rect -8521 1400 -7584 1401
rect -7528 1465 -626 1466
rect -7528 1400 -7253 1465
rect -8851 1399 -7253 1400
rect -7197 1464 -2614 1465
rect -7197 1463 -5926 1464
rect -7197 1462 -6589 1463
rect -7197 1399 -6921 1462
rect -11165 1396 -6921 1399
rect -6865 1397 -6589 1462
rect -6533 1462 -5926 1463
rect -6533 1397 -6256 1462
rect -6865 1396 -6256 1397
rect -6200 1398 -5926 1462
rect -5870 1463 -3606 1464
rect -5870 1462 -4602 1463
rect -5870 1398 -5595 1462
rect -6200 1396 -5595 1398
rect -5539 1396 -5263 1462
rect -5207 1396 -4932 1462
rect -4876 1397 -4602 1462
rect -4546 1462 -3936 1463
rect -4546 1397 -4271 1462
rect -4876 1396 -4271 1397
rect -4215 1397 -3936 1462
rect -3880 1398 -3606 1463
rect -3550 1463 -2944 1464
rect -3550 1398 -3275 1463
rect -3880 1397 -3275 1398
rect -3219 1398 -2944 1463
rect -2888 1399 -2614 1464
rect -2558 1464 -957 1465
rect -2558 1399 -2282 1464
rect -2888 1398 -2282 1399
rect -2226 1463 -1621 1464
rect -2226 1398 -1953 1463
rect -3219 1397 -1953 1398
rect -1897 1398 -1621 1463
rect -1565 1463 -957 1464
rect -1565 1398 -1289 1463
rect -1897 1397 -1289 1398
rect -1233 1399 -957 1463
rect -901 1401 -626 1465
rect -570 1402 -290 1467
rect -233 1466 547 1468
rect -233 1452 1281 1466
rect -233 1451 637 1452
rect -233 1402 83 1451
rect -570 1401 83 1402
rect -901 1399 83 1401
rect -1233 1397 83 1399
rect -4215 1396 83 1397
rect -11165 1395 83 1396
rect 142 1396 637 1451
rect 696 1396 1206 1452
rect 1265 1396 1281 1452
rect 142 1395 1281 1396
rect -11165 1392 1281 1395
rect -11165 1391 -10681 1392
rect 68 1386 1281 1392
rect 1920 1457 2061 1531
rect 2118 1529 2741 1531
rect 2118 1457 2401 1529
rect 1920 1455 2401 1457
rect 2458 1457 2741 1529
rect 2798 1460 3080 1531
rect 3137 1532 4435 1534
rect 3137 1531 3759 1532
rect 3137 1460 3420 1531
rect 2798 1457 3420 1460
rect 3477 1458 3759 1531
rect 3816 1458 4096 1532
rect 4153 1461 4435 1532
rect 4492 1461 4773 1535
rect 4830 1533 14003 1535
rect 4830 1530 13661 1533
rect 4830 1461 5148 1530
rect 4153 1458 5148 1461
rect 5204 1458 5487 1530
rect 5543 1458 5826 1530
rect 5882 1458 6167 1530
rect 6223 1529 10762 1530
rect 6223 1528 7183 1529
rect 6223 1458 6504 1528
rect 3477 1457 6504 1458
rect 2458 1456 6504 1457
rect 6560 1456 6844 1528
rect 6900 1457 7183 1528
rect 7239 1457 7523 1529
rect 7579 1457 10762 1529
rect 10818 1457 11102 1530
rect 11158 1529 11779 1530
rect 11158 1457 11441 1529
rect 6900 1456 11441 1457
rect 11497 1457 11779 1529
rect 11835 1457 13661 1530
rect 11497 1456 13661 1457
rect 2458 1455 13661 1456
rect 1920 1453 13661 1455
rect 13717 1457 14003 1533
rect 14059 1529 16320 1537
rect 14059 1459 15201 1529
rect 15257 1459 15902 1529
rect 14059 1457 15902 1459
rect 15958 1525 16320 1529
rect 15958 1458 16220 1525
rect 16306 1458 16320 1525
rect 15958 1457 16320 1458
rect 13717 1453 16320 1457
rect 1920 1451 16320 1453
rect 1920 1267 2003 1451
rect 7604 1450 16320 1451
rect 16419 1459 16440 1540
rect 16496 1459 16780 1540
rect 16836 1459 17119 1540
rect 17175 1462 17457 1540
rect 17513 1462 17819 1543
rect 17875 1462 18374 1543
rect 17175 1460 18374 1462
rect 18430 1542 19481 1543
rect 18430 1460 18922 1542
rect 17175 1459 18922 1460
rect 16419 1457 18922 1459
rect 18978 1471 19481 1542
rect 19537 1480 20031 1543
rect 20087 1480 20099 1552
rect 19537 1471 20099 1480
rect 18978 1457 20099 1471
rect 16419 1452 20099 1457
rect 20694 1539 21740 1540
rect 20694 1526 21833 1539
rect 16419 1451 19170 1452
rect 2074 1380 2160 1382
rect 16419 1380 16519 1451
rect 18366 1450 19026 1451
rect 18366 1449 18436 1450
rect 18623 1449 18736 1450
rect 18912 1449 18982 1450
rect 20694 1438 20699 1526
rect 20756 1438 21833 1526
rect 20694 1426 21833 1438
rect 2074 1297 16522 1380
rect 16680 1376 16796 1379
rect 18110 1378 18272 1379
rect 17910 1376 18049 1378
rect 16680 1367 18049 1376
rect 16680 1335 17991 1367
rect -11166 1180 2003 1267
rect 2073 1290 16522 1297
rect 16679 1293 17991 1335
rect 18048 1293 18049 1367
rect -4018 1110 -2902 1111
rect -4018 1109 -1202 1110
rect -140 1109 976 1110
rect 2073 1109 2160 1290
rect 16679 1277 18049 1293
rect 4729 1220 6711 1221
rect 4729 1219 7661 1220
rect 13941 1219 16322 1220
rect 3394 1218 16322 1219
rect 2229 1214 16322 1218
rect 2229 1213 9217 1214
rect 2229 1210 8879 1213
rect 2229 1137 7861 1210
rect 7919 1137 8201 1210
rect 8259 1209 8879 1210
rect 8259 1137 8539 1209
rect 2229 1136 8539 1137
rect 8597 1140 8879 1209
rect 8937 1141 9217 1213
rect 9275 1141 9555 1214
rect 9613 1141 9894 1214
rect 9952 1213 12117 1214
rect 9952 1141 10234 1213
rect 8937 1140 10234 1141
rect 10292 1141 12117 1213
rect 12175 1213 16322 1214
rect 12175 1141 12459 1213
rect 10292 1140 12459 1141
rect 12517 1212 16322 1213
rect 12517 1210 13133 1212
rect 12517 1140 12796 1210
rect 8597 1137 12796 1140
rect 12854 1139 13133 1210
rect 13191 1210 16242 1212
rect 13191 1209 14678 1210
rect 13191 1139 14341 1209
rect 12854 1137 14341 1139
rect 8597 1136 14341 1137
rect 14399 1137 14678 1209
rect 14736 1137 15541 1210
rect 15599 1208 16242 1210
rect 15599 1137 16228 1208
rect 14399 1136 16242 1137
rect 2229 1134 16242 1136
rect 16298 1134 16322 1212
rect 2229 1131 16322 1134
rect 2229 1129 5376 1131
rect 5679 1130 16322 1131
rect 7625 1129 16322 1130
rect 2229 1128 4359 1129
rect -4018 1107 2160 1109
rect -4998 1105 2160 1107
rect -11167 1103 -8670 1105
rect -7333 1103 2160 1105
rect -11167 1022 2160 1103
rect -11167 1018 -3882 1022
rect -3072 1021 2160 1022
rect -1220 1020 -104 1021
rect 920 1019 2160 1021
rect -11167 1016 -4949 1018
rect -11167 1011 -6000 1016
rect -8754 1009 -7317 1011
rect -5505 953 -4232 954
rect -11111 952 -9838 953
rect -7263 952 -3188 953
rect -11170 951 -9123 952
rect -8485 951 -3188 952
rect 2230 951 2311 1128
rect 16679 1053 16796 1277
rect 17910 1276 18049 1277
rect 18109 1368 18272 1378
rect 18530 1377 18607 1378
rect 18367 1376 18607 1377
rect 18109 1303 18201 1368
rect 18259 1303 18272 1368
rect 18109 1292 18272 1303
rect 18331 1363 18607 1376
rect 18331 1293 18544 1363
rect 18600 1293 18607 1363
rect 18742 1356 18815 1361
rect 18109 1205 18175 1292
rect 18331 1286 18607 1293
rect 18741 1352 18815 1356
rect 18741 1345 18753 1352
rect 18331 1211 18395 1286
rect 18741 1268 18748 1345
rect 18809 1270 18815 1352
rect 18804 1268 18815 1270
rect 18741 1255 18815 1268
rect 19240 1336 19380 1349
rect 19240 1331 19314 1336
rect 19240 1250 19255 1331
rect 19312 1251 19314 1331
rect 19370 1251 19380 1336
rect 19311 1250 19380 1251
rect 19240 1237 19380 1250
rect 19644 1316 19795 1329
rect 19644 1241 19655 1316
rect 19711 1304 19795 1316
rect 19711 1247 19721 1304
rect 19777 1247 19795 1304
rect 20859 1275 20939 1277
rect 19711 1241 19795 1247
rect 19644 1228 19795 1241
rect 20794 1265 20939 1275
rect 17728 1204 18175 1205
rect 16984 1202 18175 1204
rect 16919 1195 18175 1202
rect 16192 1051 16796 1053
rect -11170 950 -3188 951
rect -90 950 968 951
rect 1809 950 2311 951
rect -11170 949 -2166 950
rect -1318 949 2311 950
rect -11170 891 2311 949
rect 15750 1032 16796 1051
rect 15750 963 15794 1032
rect 15853 1016 16796 1032
rect 16918 1125 18175 1195
rect 18233 1138 18395 1211
rect 20794 1189 20869 1265
rect 20929 1189 20939 1265
rect 20794 1184 20939 1189
rect 20794 1143 20938 1184
rect 16918 1124 18169 1125
rect 16918 1122 17772 1124
rect 16918 1120 17707 1122
rect 15853 972 16795 1016
rect 15853 963 16792 972
rect 15750 950 16792 963
rect 15750 948 16350 950
rect -11170 890 -5077 891
rect -4461 890 2311 891
rect -11170 889 -7212 890
rect -9398 888 -8125 889
rect -3439 887 2311 890
rect -2312 886 -1039 887
rect -90 886 2311 887
rect 919 885 2311 886
rect 16055 881 16404 882
rect 16918 881 16999 1120
rect 17754 1064 18155 1065
rect 18233 1064 18290 1138
rect 17754 1021 18290 1064
rect 20252 1101 20400 1119
rect 20252 1094 20292 1101
rect 20252 1027 20279 1094
rect 20378 1032 20400 1101
rect 20357 1027 20400 1032
rect 17754 999 18289 1021
rect 20252 1003 20400 1027
rect 17754 997 18155 999
rect 16055 873 17001 881
rect 16037 801 17001 873
rect -10411 237 -5350 261
rect -10411 227 -5755 237
rect -10411 225 -8076 227
rect -10411 223 -8408 225
rect -10411 222 -9070 223
rect -10411 138 -10396 222
rect -10340 138 -10063 222
rect -10007 221 -9070 222
rect -10007 138 -9734 221
rect -10411 137 -9734 138
rect -9678 220 -9070 221
rect -9678 137 -9403 220
rect -10411 136 -9403 137
rect -9347 139 -9070 220
rect -9014 139 -8739 223
rect -8683 141 -8408 223
rect -8352 143 -8076 225
rect -8020 143 -7745 227
rect -7689 143 -7413 227
rect -7357 143 -7082 227
rect -7026 143 -6752 227
rect -6696 143 -6419 227
rect -6363 143 -6088 227
rect -6032 153 -5755 227
rect -5699 153 -5426 237
rect -5370 153 -5350 237
rect -6032 143 -5350 153
rect -5112 240 -2697 255
rect -5112 161 -5094 240
rect -5037 161 -4761 240
rect -4704 161 -4431 240
rect -4374 161 -4101 240
rect -4044 161 -3767 240
rect -3710 161 -3436 240
rect -3379 239 -2775 240
rect -3379 161 -3106 239
rect -5112 160 -3106 161
rect -3049 161 -2775 239
rect -2718 161 -2697 240
rect -3049 160 -2697 161
rect -5112 144 -2697 160
rect -2457 240 -1375 260
rect -2457 161 -2444 240
rect -2387 161 -2113 240
rect -2056 161 -1783 240
rect -1726 161 -1451 240
rect -1394 161 -1375 240
rect -2457 152 -1375 161
rect -1142 240 -708 257
rect -1142 161 -1120 240
rect -1063 161 -788 240
rect -731 161 -708 240
rect -1142 153 -708 161
rect -485 240 -376 259
rect -485 161 -457 240
rect -400 161 -376 240
rect -2452 150 -2375 152
rect -2121 150 -2044 152
rect -8352 141 -5350 143
rect -8683 139 -5350 141
rect -9347 136 -5350 139
rect -10411 116 -5350 136
rect -9499 -471 -9385 116
rect -9499 -576 -9478 -471
rect -9397 -576 -9385 -471
rect -9499 -601 -9385 -576
rect -3860 -684 -3750 144
rect -3860 -774 -3839 -684
rect -3775 -774 -3750 -684
rect -3860 -792 -3750 -774
rect -1799 -915 -1694 152
rect -1459 150 -1382 152
rect -1128 150 -907 153
rect -796 150 -719 153
rect -1799 -1001 -1789 -915
rect -1710 -1001 -1694 -915
rect -1799 -1010 -1694 -1001
rect -1007 -1139 -907 150
rect -1008 -1162 -907 -1139
rect -1008 -1241 -996 -1162
rect -924 -1241 -907 -1162
rect -1008 -1257 -907 -1241
rect -485 -1406 -376 161
rect -485 -1428 -469 -1406
rect -484 -1488 -469 -1428
rect -399 -1428 -376 -1406
rect -108 240 1 262
rect -108 161 -86 240
rect -29 161 1 240
rect -399 -1488 -380 -1428
rect -484 -1506 -380 -1488
rect -108 -1493 1 161
rect 227 240 333 258
rect 227 161 250 240
rect 307 161 333 240
rect -106 -1654 0 -1493
rect 227 -1626 333 161
rect -106 -1728 -92 -1654
rect -22 -1728 0 -1654
rect -106 -1754 0 -1728
rect 224 -1751 333 -1626
rect 450 240 559 259
rect 450 161 466 240
rect 523 161 559 240
rect 224 -1909 332 -1751
rect 450 -1872 559 161
rect 769 244 878 256
rect 769 158 805 244
rect 862 158 878 244
rect 224 -1984 241 -1909
rect 311 -1984 332 -1909
rect 224 -1998 332 -1984
rect 449 -2136 561 -1872
rect 769 -2001 878 158
rect 1011 245 1120 256
rect 1011 159 1040 245
rect 1097 159 1120 245
rect 1011 -2001 1120 159
rect 449 -2226 471 -2136
rect 538 -2226 561 -2136
rect 449 -2243 561 -2226
rect 770 -2253 877 -2001
rect 768 -2403 878 -2253
rect 768 -2484 783 -2403
rect 861 -2484 878 -2403
rect 768 -2499 878 -2484
rect 1012 -2500 1120 -2001
rect 1347 245 1456 261
rect 1347 159 1374 245
rect 1431 159 1456 245
rect 15011 204 15778 214
rect 4963 189 10474 196
rect 1347 -1996 1456 159
rect 2220 178 4699 186
rect 2220 170 3928 178
rect 2220 80 2230 170
rect 2290 80 2570 170
rect 2630 80 2910 170
rect 2970 80 3250 170
rect 3310 80 3590 170
rect 3650 80 3928 170
rect 3988 172 4699 178
rect 3988 168 4606 172
rect 3988 80 4267 168
rect 2220 78 4267 80
rect 4327 82 4606 168
rect 4666 82 4699 172
rect 4963 182 9047 189
rect 4963 179 8706 182
rect 4963 108 4976 179
rect 5032 178 8706 179
rect 5032 108 5314 178
rect 4963 107 5314 108
rect 5370 177 8706 178
rect 5370 107 5654 177
rect 4963 106 5654 107
rect 5710 106 5994 177
rect 6050 175 8706 177
rect 6050 106 6333 175
rect 4963 104 6333 106
rect 6389 104 6673 175
rect 6729 174 7351 175
rect 6729 104 7012 174
rect 4963 103 7012 104
rect 7068 104 7351 174
rect 7407 174 8028 175
rect 7407 104 7690 174
rect 7068 103 7690 104
rect 7746 104 8028 174
rect 8084 174 8706 175
rect 8084 104 8366 174
rect 7746 103 8366 104
rect 8422 111 8706 174
rect 8762 118 9047 182
rect 9103 187 10474 189
rect 9103 183 9726 187
rect 9103 118 9386 183
rect 8762 112 9386 118
rect 9442 116 9726 183
rect 9782 186 10474 187
rect 9782 116 10065 186
rect 9442 115 10065 116
rect 10121 185 10474 186
rect 10121 115 10403 185
rect 9442 114 10403 115
rect 10459 114 10474 185
rect 9442 112 10474 114
rect 8762 111 10474 112
rect 8422 103 10474 111
rect 4963 98 10474 103
rect 10581 189 13370 201
rect 10581 183 13304 189
rect 10581 182 12964 183
rect 10581 179 11608 182
rect 10581 104 10591 179
rect 10647 176 11608 179
rect 10647 173 11270 176
rect 10647 104 10931 173
rect 10581 98 10931 104
rect 10987 101 11270 173
rect 11326 107 11608 176
rect 11664 181 12288 182
rect 11664 107 11946 181
rect 11326 106 11946 107
rect 12002 107 12288 181
rect 12344 107 12626 182
rect 12682 108 12964 182
rect 13020 114 13304 183
rect 13360 114 13370 189
rect 13020 108 13370 114
rect 12682 107 13370 108
rect 12002 106 13370 107
rect 11326 101 13370 106
rect 13479 190 14917 202
rect 13479 187 14847 190
rect 13479 185 14508 187
rect 13479 184 13830 185
rect 13479 109 13492 184
rect 13548 110 13830 184
rect 13886 110 14170 185
rect 14226 112 14508 185
rect 14564 115 14847 187
rect 14903 115 14917 190
rect 14564 112 14917 115
rect 15011 198 15710 204
rect 15011 192 15371 198
rect 15011 117 15033 192
rect 15089 123 15371 192
rect 15427 129 15710 198
rect 15766 129 15778 204
rect 16037 210 16145 801
rect 16319 800 17001 801
rect 16588 222 17024 229
rect 16037 200 16146 210
rect 16037 192 16073 200
rect 15427 123 15778 129
rect 15089 117 15778 123
rect 15011 113 15778 117
rect 16040 136 16073 192
rect 16129 136 16146 200
rect 14226 110 14917 112
rect 13548 109 14917 110
rect 13479 102 14917 109
rect 10987 98 13370 101
rect 4327 78 4699 82
rect 2220 76 4699 78
rect 1347 -2468 1455 -1996
rect 1347 -2499 1458 -2468
rect 1349 -2500 1458 -2499
rect 1010 -2655 1121 -2500
rect 1010 -2735 1024 -2655
rect 1098 -2735 1121 -2655
rect 1010 -2753 1121 -2735
rect 1349 -2779 1460 -2500
rect 1349 -2929 1461 -2779
rect 1349 -3001 1365 -2929
rect 1350 -3008 1365 -3001
rect 1443 -3008 1461 -2929
rect 1350 -3030 1461 -3008
rect 2991 -3034 3117 76
rect 6921 -486 7060 98
rect 10581 96 13370 98
rect 6921 -562 6946 -486
rect 7026 -562 7060 -486
rect 6921 -586 7060 -562
rect 11886 -704 12023 96
rect 11886 -767 11915 -704
rect 12004 -767 12023 -704
rect 11886 -796 12023 -767
rect 13987 -924 14086 102
rect 13987 -987 14005 -924
rect 14067 -987 14086 -924
rect 13987 -1013 14086 -987
rect 15303 -1165 15394 113
rect 15303 -1227 15318 -1165
rect 15378 -1227 15394 -1165
rect 15303 -1258 15394 -1227
rect 15744 -1158 15879 -1140
rect 15744 -1246 15766 -1158
rect 15855 -1246 15879 -1158
rect 15744 -1258 15879 -1246
rect 16040 -1406 16146 136
rect 16588 143 16612 222
rect 16668 215 17024 222
rect 16668 143 16951 215
rect 16588 136 16951 143
rect 17007 136 17024 215
rect 16588 132 17024 136
rect 17245 224 17364 238
rect 17245 152 17289 224
rect 17345 152 17364 224
rect 16712 -495 16854 132
rect 16712 -571 16742 -495
rect 16828 -571 16854 -495
rect 16712 -589 16854 -571
rect 17245 -705 17364 152
rect 17245 -775 17270 -705
rect 17332 -775 17364 -705
rect 17245 -792 17364 -775
rect 17598 223 17708 237
rect 17598 153 17626 223
rect 17688 153 17708 223
rect 17598 -1013 17708 153
rect 17769 -1138 17849 997
rect 18343 943 18466 974
rect 18534 970 18640 971
rect 18343 874 18377 943
rect 18440 874 18466 943
rect 18343 840 18466 874
rect 18533 936 18640 970
rect 18533 867 18552 936
rect 18615 867 18640 936
rect 18533 838 18640 867
rect 18534 835 18640 838
rect 18883 935 18968 969
rect 18883 866 18893 935
rect 18956 866 18968 935
rect 18883 837 18968 866
rect 19039 936 19133 970
rect 19039 867 19058 936
rect 19121 867 19133 936
rect 19039 838 19133 867
rect 19402 935 19487 969
rect 19402 866 19412 935
rect 19475 866 19487 935
rect 19402 837 19487 866
rect 19558 936 19652 970
rect 19558 867 19577 936
rect 19640 867 19652 936
rect 19558 838 19652 867
rect 19922 935 20007 969
rect 19922 866 19932 935
rect 19995 866 20007 935
rect 19922 837 20007 866
rect 20078 936 20172 970
rect 20078 867 20097 936
rect 20160 867 20172 936
rect 20078 838 20172 867
rect 20454 935 20539 969
rect 20454 866 20464 935
rect 20527 866 20539 935
rect 20454 837 20539 866
rect 20610 936 20704 970
rect 20610 867 20629 936
rect 20692 867 20704 936
rect 20610 838 20704 867
rect 20794 731 20874 1143
rect 20972 935 21057 969
rect 20972 866 20982 935
rect 21045 866 21057 935
rect 20972 837 21057 866
rect 21128 936 21222 970
rect 21128 867 21147 936
rect 21210 867 21222 936
rect 21128 838 21222 867
rect 20361 725 20431 729
rect 20781 725 20874 731
rect 20361 724 20949 725
rect 18271 702 18360 714
rect 18271 635 18287 702
rect 18347 635 18360 702
rect 18271 625 18360 635
rect 18795 706 18865 718
rect 18795 635 18804 706
rect 18860 635 18865 706
rect 18795 624 18865 635
rect 19313 706 19383 718
rect 20361 717 20950 724
rect 19313 635 19322 706
rect 19378 635 19383 706
rect 19313 624 19383 635
rect 19833 705 19903 717
rect 19833 634 19842 705
rect 19898 634 19903 705
rect 20361 646 20370 717
rect 20426 712 20950 717
rect 20426 646 20889 712
rect 20361 641 20889 646
rect 20945 641 20950 712
rect 20361 635 20950 641
rect 19833 623 19903 634
rect 20365 631 20950 635
rect 20880 630 20950 631
rect 18625 532 18692 536
rect 18624 523 18692 532
rect 19137 527 19203 531
rect 18624 447 18630 523
rect 18686 447 18692 523
rect 18624 440 18692 447
rect 18625 436 18692 440
rect 19136 518 19203 527
rect 19654 525 19720 529
rect 20173 525 20239 529
rect 20704 525 20770 529
rect 21221 525 21287 529
rect 19136 442 19142 518
rect 19198 442 19203 518
rect 19136 435 19203 442
rect 19137 432 19203 435
rect 19653 516 19720 525
rect 19653 440 19659 516
rect 19715 440 19720 516
rect 19653 433 19720 440
rect 20172 516 20239 525
rect 20172 440 20178 516
rect 20234 440 20239 516
rect 20172 433 20239 440
rect 20703 516 20770 525
rect 20703 440 20709 516
rect 20765 440 20770 516
rect 20703 433 20770 440
rect 21220 516 21287 525
rect 21220 440 21226 516
rect 21282 440 21287 516
rect 21220 433 21287 440
rect 19654 430 19720 433
rect 20173 430 20239 433
rect 20704 430 20770 433
rect 21221 430 21287 433
rect 18052 188 18162 200
rect 18052 131 18079 188
rect 18148 131 18162 188
rect 17760 -1210 17853 -1138
rect 16040 -1489 16058 -1406
rect 16128 -1489 16146 -1406
rect 16040 -1508 16146 -1489
rect 17761 -1653 17853 -1210
rect 17761 -1735 17775 -1653
rect 17836 -1735 17853 -1653
rect 17761 -1751 17853 -1735
rect 18052 -2141 18162 131
rect 18439 131 18540 139
rect 18439 35 18462 131
rect 18519 35 18540 131
rect 18439 -1642 18540 35
rect 18439 -1730 18451 -1642
rect 18527 -1730 18540 -1642
rect 18439 -1752 18540 -1730
rect 18948 126 19049 142
rect 18948 30 18972 126
rect 19029 30 19049 126
rect 18948 -1899 19049 30
rect 18948 -1973 18964 -1899
rect 19026 -1973 19049 -1899
rect 18948 -1995 19049 -1973
rect 19473 130 19578 145
rect 19473 34 19490 130
rect 19547 34 19578 130
rect 18052 -2224 18066 -2141
rect 18137 -2224 18162 -2141
rect 18052 -2249 18162 -2224
rect 19473 -2140 19578 34
rect 19473 -2231 19490 -2140
rect 19561 -2231 19578 -2140
rect 19473 -2254 19578 -2231
rect 19995 132 20100 158
rect 19995 36 20009 132
rect 20073 68 20100 132
rect 20066 36 20100 68
rect 19995 -2400 20100 36
rect 19995 -2491 20014 -2400
rect 20085 -2491 20100 -2400
rect 19995 -2500 20100 -2491
rect 20527 134 20627 145
rect 20527 38 20543 134
rect 20600 118 20627 134
rect 20608 48 20627 118
rect 20600 38 20627 48
rect 20527 -2635 20627 38
rect 20527 -2726 20548 -2635
rect 20619 -2726 20627 -2635
rect 20527 -2752 20627 -2726
rect 21038 130 21133 147
rect 21038 112 21061 130
rect 21038 44 21055 112
rect 21038 34 21061 44
rect 21118 34 21133 130
rect 2989 -3212 3117 -3034
rect 21038 -2923 21133 34
rect 21038 -3014 21050 -2923
rect 21121 -3014 21133 -2923
rect 21038 -3035 21133 -3014
rect 2989 -3291 3009 -3212
rect 3096 -3291 3117 -3212
rect 2989 -3310 3117 -3291
<< via3 >>
rect 16220 1458 16306 1525
rect 16228 1137 16242 1208
rect 16242 1137 16297 1208
rect 18748 1270 18753 1345
rect 18753 1270 18804 1345
rect 18748 1268 18804 1270
rect 19255 1251 19312 1331
rect 19255 1250 19311 1251
rect 19721 1247 19777 1304
rect 15794 963 15853 1032
rect 20279 1032 20292 1094
rect 20292 1032 20357 1094
rect 20279 1027 20357 1032
rect 15766 -1246 15855 -1158
rect 18377 874 18440 943
rect 18552 867 18615 936
rect 18893 866 18956 935
rect 19058 867 19121 936
rect 19412 866 19475 935
rect 19577 867 19640 936
rect 19932 866 19995 935
rect 20097 867 20160 936
rect 20464 866 20527 935
rect 20629 867 20692 936
rect 20982 866 21045 935
rect 21147 867 21210 936
rect 18287 635 18346 702
rect 18346 635 18347 702
rect 18804 636 18860 706
rect 19322 636 19378 706
rect 19842 635 19898 705
rect 20370 647 20426 717
rect 20889 642 20945 712
rect 18630 447 18686 523
rect 19142 442 19198 518
rect 19659 440 19715 516
rect 20178 440 20234 516
rect 20709 440 20765 516
rect 21226 440 21282 516
rect 18972 32 19029 119
rect 20015 68 20066 132
rect 20066 68 20073 132
rect 20545 48 20600 118
rect 20600 48 20608 118
rect 21055 44 21061 112
rect 21061 44 21111 112
<< metal4 >>
rect 18184 1542 18280 1547
rect 16207 1525 18280 1542
rect 16207 1458 16220 1525
rect 16306 1458 18280 1525
rect 16207 1449 18280 1458
rect 16211 1208 18106 1226
rect 16211 1137 16228 1208
rect 16297 1137 18106 1208
rect 16211 1126 18106 1137
rect 15755 1044 15881 1051
rect 15743 1032 15881 1044
rect 15743 963 15794 1032
rect 15853 963 15881 1032
rect 15743 946 15881 963
rect 15743 -1158 15879 946
rect 17993 535 18099 1126
rect 18184 717 18280 1449
rect 18343 943 18467 2430
rect 18534 970 18647 2430
rect 18730 1348 18810 1360
rect 18730 1267 18737 1348
rect 18730 1258 18810 1267
rect 18741 1255 18810 1258
rect 18343 874 18377 943
rect 18440 874 18467 943
rect 18343 840 18467 874
rect 18533 936 18647 970
rect 18533 867 18552 936
rect 18615 867 18647 936
rect 18533 838 18647 867
rect 18534 835 18647 838
rect 18866 935 18973 2430
rect 18866 866 18893 935
rect 18956 866 18973 935
rect 18866 833 18973 866
rect 19039 936 19146 2429
rect 19239 1335 19325 1350
rect 19239 1250 19242 1335
rect 19313 1250 19325 1335
rect 19239 1237 19325 1250
rect 19039 867 19058 936
rect 19121 867 19146 936
rect 19039 832 19146 867
rect 19383 935 19490 2429
rect 19383 866 19412 935
rect 19475 866 19490 935
rect 19383 832 19490 866
rect 19557 936 19664 2430
rect 19720 1309 19811 1329
rect 19720 1304 19730 1309
rect 19720 1247 19721 1304
rect 19720 1238 19730 1247
rect 19803 1238 19811 1309
rect 19720 1229 19811 1238
rect 19725 1228 19811 1229
rect 19557 867 19577 936
rect 19640 867 19664 936
rect 19557 833 19664 867
rect 19905 935 20012 2430
rect 19905 866 19932 935
rect 19995 866 20012 935
rect 19905 833 20012 866
rect 20077 936 20184 2430
rect 20251 1105 20382 1121
rect 20251 1012 20262 1105
rect 20371 1012 20382 1105
rect 20251 1003 20382 1012
rect 20077 867 20097 936
rect 20160 867 20184 936
rect 20077 833 20184 867
rect 20442 935 20549 2427
rect 20442 866 20464 935
rect 20527 866 20549 935
rect 20442 830 20549 866
rect 20607 936 20714 2430
rect 20607 867 20629 936
rect 20692 867 20714 936
rect 20607 833 20714 867
rect 20962 935 21069 2429
rect 20962 866 20982 935
rect 21045 866 21069 935
rect 20962 832 21069 866
rect 21128 936 21235 2432
rect 21128 867 21147 936
rect 21210 867 21235 936
rect 21128 835 21235 867
rect 18779 717 20958 729
rect 18184 706 20370 717
rect 18184 702 18804 706
rect 18184 635 18287 702
rect 18347 636 18804 702
rect 18860 636 19322 706
rect 19378 705 20370 706
rect 19378 636 19842 705
rect 18347 635 19842 636
rect 19898 647 20370 705
rect 20426 712 20958 717
rect 20426 647 20889 712
rect 19898 642 20889 647
rect 20945 642 20958 712
rect 19898 635 20958 642
rect 18184 625 20958 635
rect 18184 618 18280 625
rect 18779 624 20958 625
rect 19832 623 19904 624
rect 18936 535 21293 537
rect 17993 523 21293 535
rect 17993 447 18630 523
rect 18686 518 21293 523
rect 18686 447 19142 518
rect 17993 442 19142 447
rect 19198 516 21293 518
rect 19198 442 19659 516
rect 17993 440 19659 442
rect 19715 440 20178 516
rect 20234 440 20709 516
rect 20765 440 21226 516
rect 21282 440 21293 516
rect 17993 438 21293 440
rect 18119 437 21293 438
rect 18936 436 21293 437
rect 19136 432 19203 436
rect 19653 430 19720 436
rect 20172 430 20239 436
rect 20703 430 20770 436
rect 21220 430 21287 436
rect 19995 141 20098 155
rect 18951 119 19042 137
rect 18951 118 18972 119
rect 18951 31 18970 118
rect 19029 32 19042 119
rect 19995 68 20015 141
rect 20080 68 20098 141
rect 19995 50 20098 68
rect 20518 118 20627 147
rect 19027 31 19042 32
rect 18951 13 19042 31
rect 20518 44 20540 118
rect 20614 44 20627 118
rect 20518 12 20627 44
rect 21037 116 21130 141
rect 21037 42 21052 116
rect 21112 42 21130 116
rect 21037 25 21130 42
rect 15743 -1246 15766 -1158
rect 15855 -1246 15879 -1158
rect 15743 -1258 15879 -1246
<< via4 >>
rect 18737 1345 18810 1348
rect 18737 1268 18748 1345
rect 18748 1268 18804 1345
rect 18804 1268 18810 1345
rect 18737 1267 18810 1268
rect 19242 1331 19313 1335
rect 19242 1250 19255 1331
rect 19255 1251 19312 1331
rect 19312 1251 19313 1331
rect 19255 1250 19311 1251
rect 19311 1250 19313 1251
rect 19730 1304 19803 1309
rect 19730 1247 19777 1304
rect 19777 1247 19803 1304
rect 19730 1238 19803 1247
rect 20262 1094 20371 1105
rect 20262 1027 20279 1094
rect 20279 1027 20357 1094
rect 20357 1027 20371 1094
rect 20262 1012 20371 1027
rect 18970 32 18972 118
rect 18972 32 19027 118
rect 20015 132 20080 141
rect 20015 68 20073 132
rect 20073 68 20080 132
rect 18970 31 19027 32
rect 20540 48 20545 118
rect 20545 48 20608 118
rect 20608 48 20614 118
rect 20540 44 20614 48
rect 21052 112 21112 116
rect 21052 44 21055 112
rect 21055 44 21111 112
rect 21111 44 21112 112
rect 21052 42 21112 44
<< metal5 >>
rect 18684 1348 18827 1380
rect 18684 1267 18737 1348
rect 18810 1267 18827 1348
rect 18684 1204 18827 1267
rect 19197 1335 19358 1389
rect 19197 1250 19242 1335
rect 19313 1250 19358 1335
rect 19197 1206 19358 1250
rect 19681 1309 19826 1351
rect 19681 1238 19730 1309
rect 19803 1238 19826 1309
rect 18721 144 18815 1204
rect 19214 155 19309 1206
rect 19681 1194 19826 1238
rect 19726 430 19820 1194
rect 20237 1105 20399 1134
rect 20237 1012 20262 1105
rect 20371 1094 20399 1105
rect 20371 1089 21135 1094
rect 20371 1012 21144 1089
rect 20237 987 21144 1012
rect 19726 416 20640 430
rect 19726 336 20641 416
rect 18721 118 19054 144
rect 18721 31 18970 118
rect 19027 31 19054 118
rect 19214 141 20099 155
rect 19214 68 20015 141
rect 20080 68 20099 141
rect 19214 49 20099 68
rect 20516 118 20641 336
rect 18721 11 19054 31
rect 20516 44 20540 118
rect 20614 44 20641 118
rect 20516 8 20641 44
rect 21034 116 21144 987
rect 21034 42 21052 116
rect 21112 42 21144 116
rect 21034 4 21144 42
<< labels >>
flabel metal3 -11165 1391 -11005 1475 0 FreeSans 320 0 0 0 VREF
port 3 nsew
flabel metal3 1288 2300 1395 2407 0 FreeSans 160 0 0 0 EN_VREF_Z[0]
port 30 nsew
flabel metal3 1074 2301 1181 2407 0 FreeSans 160 0 0 0 EN_VREF_Z[1]
port 29 nsew
flabel metal3 719 2300 826 2407 0 FreeSans 160 0 0 0 EN_VREF_Z[2]
port 28 nsew
flabel metal3 504 2301 611 2408 0 FreeSans 160 0 0 0 EN_VREF_Z[3]
port 27 nsew
flabel metal3 165 2303 271 2410 0 FreeSans 160 0 0 0 EN_VREF_Z[4]
port 26 nsew
flabel metal3 -48 2304 59 2410 0 FreeSans 160 0 0 0 EN_VREF_Z[5]
port 25 nsew
flabel metal3 -478 2297 -370 2409 0 FreeSans 160 0 0 0 EN_VREF_Z[6]
port 24 nsew
flabel metal3 -970 2298 -862 2410 0 FreeSans 160 0 0 0 EN_VREF_Z[7]
port 23 nsew
flabel metal3 -1931 2297 -1822 2412 0 FreeSans 160 0 0 0 EN_VREF_Z[8]
port 22 nsew
flabel metal3 -3656 2300 -3547 2415 0 FreeSans 160 0 0 0 EN_VREF_Z[9]
port 21 nsew
flabel metal3 -7644 2297 -7535 2411 0 FreeSans 160 0 0 0 EN_VREF_Z[10]
port 20 nsew
flabel metal3 3240 2310 3379 2411 0 FreeSans 160 0 0 0 EN_VCM_SW
port 54 nsew
flabel metal3 6415 2307 6554 2408 0 FreeSans 160 0 0 0 EN_VCM[10]
port 42 nsew
flabel metal3 11194 2306 11332 2410 0 FreeSans 160 0 0 0 EN_VCM[9]
port 43 nsew
flabel metal3 13839 2295 13978 2408 0 FreeSans 160 0 0 0 EN_VCM[8]
port 44 nsew
flabel metal3 15158 2286 15297 2406 0 FreeSans 160 0 0 0 EN_VCM[7]
port 45 nsew
flabel metal3 15931 2297 16042 2416 0 FreeSans 160 0 0 0 EN_VCM[6]
port 46 nsew
flabel metal3 8869 2299 9007 2410 0 FreeSans 160 0 0 0 EN_VSS[10]
port 31 nsew
flabel metal3 12610 2294 12749 2407 0 FreeSans 160 0 0 0 EN_VSS[9]
port 32 nsew
flabel metal3 14527 2295 14666 2408 0 FreeSans 160 0 0 0 EN_VSS[8]
port 33 nsew
flabel metal3 15497 2288 15634 2399 0 FreeSans 160 0 0 0 EN_VSS[7]
port 34 nsew
flabel metal3 16155 2299 16263 2411 0 FreeSans 160 0 0 0 EN_VSS[6]
port 35 nsew
flabel metal3 16729 2310 16873 2429 0 FreeSans 160 0 0 0 EN_VIN
port 19 nsew
flabel metal3 -11167 1011 -11029 1105 0 FreeSans 320 0 0 0 VIN
port 4 nsew
flabel metal3 -11163 894 -11016 949 0 FreeSans 160 0 0 0 VREF_GND
port 2 nsew
flabel metal4 18345 2332 18464 2423 0 FreeSans 160 0 0 0 EN_VCM[5]
port 47 nsew
flabel metal4 20967 2328 21058 2420 0 FreeSans 160 0 0 0 EN_VCM[0]
port 52 nsew
flabel metal4 20447 2333 20538 2425 0 FreeSans 160 0 0 0 EN_VCM[1]
port 51 nsew
flabel metal4 19911 2329 20002 2421 0 FreeSans 160 0 0 0 EN_VCM[2]
port 50 nsew
flabel metal4 19390 2329 19481 2421 0 FreeSans 160 0 0 0 EN_VCM[3]
port 49 nsew
flabel metal4 18874 2331 18965 2423 0 FreeSans 160 0 0 0 EN_VCM[4]
port 48 nsew
flabel metal3 -11166 1180 -11013 1267 0 FreeSans 320 0 0 0 VCM
port 1 nsew
flabel metal3 20780 2198 20868 2280 0 FreeSans 160 0 0 0 EN_VCM_DUMMY
port 53 nsew
flabel metal2 21590 -587 21768 -476 0 FreeSans 160 0 0 0 Cbtm_10
port 17 nsew
flabel metal2 21593 -786 21771 -675 0 FreeSans 160 0 0 0 Cbtm_9
port 16 nsew
flabel metal2 21595 -1005 21771 -903 0 FreeSans 160 0 0 0 Cbtm_8
port 15 nsew
flabel metal2 21596 -1251 21772 -1149 0 FreeSans 160 0 0 0 Cbtm_7
port 14 nsew
flabel metal2 21591 -1505 21767 -1403 0 FreeSans 160 0 0 0 Cbtm_6
port 13 nsew
flabel metal2 21590 -1743 21766 -1641 0 FreeSans 160 0 0 0 Cbtm_5
port 12 nsew
flabel metal2 21590 -1990 21766 -1888 0 FreeSans 160 0 0 0 Cbtm_4
port 11 nsew
flabel metal2 21587 -2237 21763 -2135 0 FreeSans 160 0 0 0 Cbtm_3
port 10 nsew
flabel metal2 21589 -2495 21765 -2393 0 FreeSans 160 0 0 0 Cbtm_2
port 9 nsew
flabel metal2 21586 -2745 21762 -2643 0 FreeSans 160 0 0 0 Cbtm_1
port 8 nsew
flabel metal2 21592 -3021 21768 -2919 0 FreeSans 160 0 0 0 Cbtm_0
port 7 nsew
flabel metal3 21687 1428 21740 1540 0 FreeSans 320 0 0 0 Cbtm_0_dummy
port 6 nsew
flabel metal2 16963 2002 17427 2105 0 FreeSans 320 0 0 0 VSS
port 55 nsew
flabel metal3 21588 -3304 21769 -3181 0 FreeSans 160 0 0 0 VDAC
port 18 nsew
flabel metal2 -4756 2003 -4292 2106 0 FreeSans 320 0 0 0 VDD
port 5 nsew
flabel metal4 21136 2325 21229 2425 0 FreeSans 160 0 0 0 EN_VSS[0]
port 41 nsew
flabel metal4 20612 2321 20705 2421 0 FreeSans 160 0 0 0 EN_VSS[1]
port 40 nsew
flabel metal4 20082 2325 20175 2425 0 FreeSans 160 0 0 0 EN_VSS[2]
port 39 nsew
flabel metal4 19564 2323 19657 2423 0 FreeSans 160 0 0 0 EN_VSS[3]
port 38 nsew
flabel metal4 19047 2324 19140 2424 0 FreeSans 160 0 0 0 EN_VSS[4]
port 37 nsew
flabel metal4 18541 2323 18634 2423 0 FreeSans 160 0 0 0 EN_VSS[5]
port 36 nsew
<< end >>
