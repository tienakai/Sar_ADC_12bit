magic
tech gf180mcuD
magscale 1 10
timestamp 1757847982
<< nwell >>
rect -442 -330 442 330
<< pmos >>
rect -268 -200 -212 200
rect -108 -200 -52 200
rect 52 -200 108 200
rect 212 -200 268 200
<< pdiff >>
rect -356 187 -268 200
rect -356 -187 -343 187
rect -297 -187 -268 187
rect -356 -200 -268 -187
rect -212 187 -108 200
rect -212 -187 -183 187
rect -137 -187 -108 187
rect -212 -200 -108 -187
rect -52 187 52 200
rect -52 -187 -23 187
rect 23 -187 52 187
rect -52 -200 52 -187
rect 108 187 212 200
rect 108 -187 137 187
rect 183 -187 212 187
rect 108 -200 212 -187
rect 268 187 356 200
rect 268 -187 297 187
rect 343 -187 356 187
rect 268 -200 356 -187
<< pdiffc >>
rect -343 -187 -297 187
rect -183 -187 -137 187
rect -23 -187 23 187
rect 137 -187 183 187
rect 297 -187 343 187
<< polysilicon >>
rect -268 200 -212 244
rect -108 200 -52 244
rect 52 200 108 244
rect 212 200 268 244
rect -268 -244 -212 -200
rect -108 -244 -52 -200
rect 52 -244 108 -200
rect 212 -244 268 -200
<< metal1 >>
rect -343 187 -297 198
rect -343 -198 -297 -187
rect -183 187 -137 198
rect -183 -198 -137 -187
rect -23 187 23 198
rect -23 -198 23 -187
rect 137 187 183 198
rect 137 -198 183 -187
rect 297 187 343 198
rect 297 -198 343 -187
<< properties >>
string gencell pfet_03v3
string library gf180mcu
string parameters w 2 l 0.280 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {pfet_03v3 pfet_06v0}
<< end >>
