magic
tech gf180mcuD
magscale 1 10
timestamp 1757728064
<< nwell >>
rect 1780 6981 3280 7130
rect 1773 6930 3280 6981
rect 1773 6919 2564 6930
rect 2334 4930 2421 6919
rect 1975 4872 2146 4928
rect 1949 4858 2166 4868
rect 2250 4610 2520 4930
rect 7102 4843 7332 4937
rect 7934 4551 8029 6894
rect 6525 789 6714 790
rect 2724 220 2925 789
rect 6525 751 6612 789
rect 6525 669 6656 751
rect 10313 752 10439 789
rect 2600 90 2925 220
rect 6525 114 6612 669
rect 2642 29 2925 90
rect 6432 33 6680 114
rect 10306 670 10565 752
rect 10313 113 10439 670
rect 2724 -1 2925 29
rect 6525 0 6612 33
rect 10237 31 10496 113
rect 10313 0 10439 31
rect 10313 -1 10485 0
<< pwell >>
rect 909 10430 6786 10593
rect 3292 4552 6377 6995
rect 40 740 420 1160
rect 4602 669 4728 751
rect 8434 749 8468 791
rect 8396 671 8527 749
rect 3831 371 3833 438
rect 773 30 914 112
rect 4627 33 4717 112
rect 8434 113 8468 671
rect 8412 30 8493 113
rect 8434 1 8468 30
<< ndiff >>
rect 3831 371 3833 438
<< psubdiff >>
rect 773 30 914 112
<< nsubdiff >>
rect 2275 4638 2490 4803
<< polysilicon >>
rect 1163 10299 1449 10320
rect 1163 10206 1188 10299
rect 1425 10206 1449 10299
rect 2776 10300 3062 10323
rect 2776 10209 2801 10300
rect 3040 10209 3062 10300
rect 5616 10305 5902 10320
rect 5616 10206 5639 10305
rect 5889 10206 5902 10305
rect 9779 10300 10065 10323
rect 9779 10209 9805 10300
rect 10045 10209 10065 10300
rect 13879 10280 14168 10295
rect 13879 10189 13913 10280
rect 14146 10189 14168 10280
rect 13879 10165 14168 10189
rect 1030 6047 1046 6117
rect 1110 6047 1123 6117
rect 1030 6030 1123 6047
rect 2730 4931 2994 4947
rect 1342 4600 1433 4883
rect 1949 4872 1975 4919
rect 2146 4872 2166 4919
rect 1532 4601 1622 4867
rect 1949 4858 2166 4872
rect 2730 4878 2775 4931
rect 2945 4878 2994 4931
rect 2730 4861 2994 4878
rect 1341 4530 1434 4600
rect 1531 4532 1624 4601
rect 3518 4544 3580 4909
rect 3511 4541 3580 4544
rect 1266 4514 1436 4530
rect 1266 4433 1281 4514
rect 1416 4433 1436 4514
rect 1530 4529 1700 4532
rect 1530 4514 1702 4529
rect 1530 4475 1546 4514
rect 1266 4420 1436 4433
rect 1529 4433 1546 4475
rect 1682 4433 1702 4514
rect 1529 4419 1702 4433
rect 3467 4520 3638 4541
rect 3867 4539 3923 4909
rect 3467 4439 3487 4520
rect 3622 4439 3638 4520
rect 3467 4424 3638 4439
rect 3823 4518 3994 4539
rect 4250 4534 4315 5688
rect 7103 4937 7333 4939
rect 7102 4923 7333 4937
rect 4609 4536 4678 4903
rect 5121 4543 5197 4889
rect 5112 4541 5240 4543
rect 5863 4541 5939 4894
rect 7102 4856 7125 4923
rect 7312 4856 7333 4923
rect 7102 4845 7333 4856
rect 7102 4843 7332 4845
rect 9311 4548 9430 4915
rect 11469 4550 11574 4912
rect 12938 4550 13040 4910
rect 11469 4549 11580 4550
rect 9302 4546 9430 4548
rect 4234 4533 4315 4534
rect 3823 4437 3843 4518
rect 3978 4437 3994 4518
rect 3823 4422 3994 4437
rect 4189 4513 4343 4533
rect 4189 4435 4216 4513
rect 4327 4435 4343 4513
rect 4189 4420 4343 4435
rect 4564 4516 4718 4536
rect 4564 4438 4591 4516
rect 4702 4438 4718 4516
rect 4564 4422 4718 4438
rect 5079 4520 5251 4541
rect 5845 4539 5973 4541
rect 5079 4439 5100 4520
rect 5235 4439 5251 4520
rect 5079 4424 5251 4439
rect 5812 4518 5984 4539
rect 5812 4437 5833 4518
rect 5968 4437 5984 4518
rect 5812 4422 5984 4437
rect 9269 4525 9441 4546
rect 9269 4444 9290 4525
rect 9425 4444 9441 4525
rect 9269 4429 9441 4444
rect 11436 4528 11608 4549
rect 11436 4447 11457 4528
rect 11592 4447 11608 4528
rect 11436 4432 11608 4447
rect 12895 4529 13068 4550
rect 13836 4546 13939 4911
rect 12895 4448 12917 4529
rect 13052 4448 13068 4529
rect 12895 4433 13068 4448
rect 13798 4529 13970 4546
rect 13798 4448 13829 4529
rect 13952 4448 13970 4529
rect 13798 4430 13970 4448
rect 1017 996 1139 1013
rect 1017 919 1033 996
rect 1123 919 1139 996
rect 1017 905 1139 919
rect 1353 986 1474 1003
rect 1353 909 1368 986
rect 1458 909 1474 986
rect 1047 642 1123 905
rect 1353 895 1474 909
rect 1601 985 1722 1002
rect 1601 908 1616 985
rect 1706 908 1722 985
rect 1373 894 1458 895
rect 1601 894 1722 908
rect 2242 986 2363 1003
rect 2242 909 2257 986
rect 2347 909 2363 986
rect 2242 895 2363 909
rect 3166 977 3287 994
rect 3166 900 3181 977
rect 3271 900 3287 977
rect 2269 894 2347 895
rect 1373 642 1449 894
rect 1622 893 1706 894
rect 1622 643 1674 893
rect 2269 644 2321 894
rect 3166 886 3287 900
rect 3807 976 3928 993
rect 3807 899 3822 976
rect 3912 899 3928 976
rect 3195 885 3271 886
rect 3807 885 3928 899
rect 4047 981 4168 998
rect 4047 904 4062 981
rect 4152 904 4168 981
rect 4047 890 4168 904
rect 4387 983 4508 1000
rect 4387 906 4402 983
rect 4492 906 4508 983
rect 4387 892 4508 906
rect 4823 980 4944 997
rect 4823 903 4838 980
rect 4928 903 4944 980
rect 4416 891 4492 892
rect 4076 889 4152 890
rect 3196 641 3248 885
rect 3836 884 3912 885
rect 3849 639 3901 884
rect 4096 640 4148 889
rect 4420 638 4472 891
rect 4823 889 4944 903
rect 5142 988 5263 1005
rect 5142 911 5157 988
rect 5247 911 5263 988
rect 5142 897 5263 911
rect 5391 987 5512 1004
rect 5391 910 5406 987
rect 5496 910 5512 987
rect 5171 896 5247 897
rect 5391 896 5512 910
rect 5992 991 6113 1008
rect 5992 914 6007 991
rect 6097 914 6113 991
rect 5992 900 6113 914
rect 6950 985 7071 1002
rect 6950 908 6965 985
rect 7055 908 7071 985
rect 6021 899 6097 900
rect 4852 888 4928 889
rect 4857 640 4909 888
rect 5180 639 5232 896
rect 5420 895 5496 896
rect 5423 640 5475 895
rect 6027 642 6079 899
rect 6950 894 7071 908
rect 7616 971 7737 988
rect 7616 894 7631 971
rect 7721 894 7737 971
rect 6979 893 7055 894
rect 6990 641 7042 893
rect 7616 880 7737 894
rect 7857 979 7978 996
rect 7857 902 7872 979
rect 7962 902 7978 979
rect 7857 888 7978 902
rect 8161 984 8282 1001
rect 8161 907 8176 984
rect 8266 907 8282 984
rect 8161 893 8282 907
rect 8605 978 8726 995
rect 8605 901 8620 978
rect 8710 901 8726 978
rect 8190 892 8266 893
rect 7886 887 7962 888
rect 7640 879 7721 880
rect 7640 640 7693 879
rect 7887 641 7940 887
rect 8191 640 8244 892
rect 8605 887 8726 901
rect 8938 981 9059 998
rect 8938 904 8953 981
rect 9043 904 9059 981
rect 8938 890 9059 904
rect 9156 980 9277 997
rect 9156 903 9171 980
rect 9261 903 9277 980
rect 8967 889 9043 890
rect 9156 889 9277 903
rect 9766 979 9887 996
rect 9766 902 9781 979
rect 9871 902 9887 979
rect 8634 886 8710 887
rect 8649 639 8702 886
rect 8978 639 9031 889
rect 9185 888 9263 889
rect 9766 888 9887 902
rect 10704 984 10825 1001
rect 10704 907 10719 984
rect 10809 907 10825 984
rect 10704 893 10825 907
rect 11396 989 11517 1006
rect 11396 912 11411 989
rect 11501 912 11517 989
rect 11396 898 11517 912
rect 11633 997 11754 1014
rect 11633 920 11648 997
rect 11738 920 11754 997
rect 11633 906 11754 920
rect 11969 986 12090 1003
rect 11969 909 11984 986
rect 12074 909 12090 986
rect 11662 905 11738 906
rect 11425 897 11501 898
rect 10733 892 10809 893
rect 9210 638 9263 888
rect 9795 887 9871 888
rect 9808 640 9861 887
rect 10748 638 10801 892
rect 11440 640 11493 897
rect 11675 641 11728 905
rect 11969 895 12090 909
rect 11998 894 12074 895
rect 12010 641 12063 894
<< polycontact >>
rect 1188 10198 1425 10299
rect 2801 10206 3040 10300
rect 5639 10196 5889 10305
rect 9805 10198 10045 10300
rect 13913 10189 14146 10280
rect 1046 6047 1110 6117
rect 1975 4872 2146 4928
rect 2775 4878 2945 4931
rect 1281 4433 1416 4514
rect 1546 4433 1682 4514
rect 3487 4439 3622 4520
rect 7125 4856 7312 4923
rect 3843 4437 3978 4518
rect 4216 4435 4327 4513
rect 4591 4438 4702 4516
rect 5100 4439 5235 4520
rect 5833 4437 5968 4518
rect 9290 4444 9425 4525
rect 11457 4447 11592 4528
rect 12917 4448 13052 4529
rect 13829 4448 13952 4529
rect 155 1018 306 1108
rect 1033 919 1123 996
rect 1368 909 1458 986
rect 524 806 689 899
rect 1616 908 1706 985
rect 2257 909 2347 986
rect 3181 900 3271 977
rect 3822 899 3912 976
rect 4062 904 4152 981
rect 4402 906 4492 983
rect 4838 903 4928 980
rect 5157 911 5247 988
rect 5406 910 5496 987
rect 6007 914 6097 991
rect 6965 908 7055 985
rect 7631 894 7721 971
rect 7872 902 7962 979
rect 8176 907 8266 984
rect 8620 901 8710 978
rect 8953 904 9043 981
rect 9171 903 9261 980
rect 9781 902 9871 979
rect 10719 907 10809 984
rect 11411 912 11501 989
rect 11648 920 11738 997
rect 11984 909 12074 986
<< metal1 >>
rect 6739 10593 7306 10594
rect 909 10430 7306 10593
rect 12522 10593 14560 10594
rect 12522 10592 15584 10593
rect 12522 10570 16212 10592
rect 12522 10475 15719 10570
rect 16169 10475 16212 10570
rect 12522 10432 16212 10475
rect 14539 10430 16212 10432
rect 6739 10429 7306 10430
rect 1166 10299 1449 10320
rect 1166 10198 1188 10299
rect 1426 10202 1449 10299
rect 1425 10198 1449 10202
rect 1166 10189 1449 10198
rect 2779 10300 3057 10317
rect 2779 10206 2801 10300
rect 3040 10206 3057 10300
rect 2779 10194 3057 10206
rect 5623 10305 5897 10313
rect 5623 10196 5639 10305
rect 5889 10196 5897 10305
rect 5623 10184 5897 10196
rect 9791 10300 10056 10316
rect 9791 10198 9805 10300
rect 10045 10198 10056 10300
rect 9791 10189 10056 10198
rect 13880 10280 14168 10296
rect 13880 10189 13913 10280
rect 14146 10189 14168 10280
rect 13880 10172 14168 10189
rect -491 10119 675 10120
rect -491 10113 789 10119
rect -491 10049 -479 10113
rect -348 10109 789 10113
rect -348 10051 677 10109
rect 779 10051 789 10109
rect -348 10049 789 10051
rect -491 10040 789 10049
rect 644 10039 789 10040
rect 12513 8371 14560 8374
rect 16204 8373 16430 8375
rect 16204 8372 16435 8373
rect 7047 8369 14560 8371
rect 15567 8369 16963 8372
rect 7047 8349 16963 8369
rect 7047 8246 16480 8349
rect 16937 8246 16963 8349
rect 7047 8213 16963 8246
rect 7047 8212 14560 8213
rect 15567 8210 16963 8213
rect 1652 6723 3381 6870
rect 6275 6695 8189 6847
rect 14078 6808 14560 6814
rect 15567 6811 16211 6812
rect 16407 6811 16966 6812
rect 15567 6808 16966 6811
rect 14078 6773 16966 6808
rect 14078 6678 16496 6773
rect 16910 6678 16966 6773
rect 14078 6642 16966 6678
rect 14496 6639 16966 6642
rect 16191 6638 16416 6639
rect 954 6361 1033 6377
rect 954 6285 956 6361
rect 1030 6285 1033 6361
rect 954 6271 1033 6285
rect 1030 6118 1121 6150
rect 1030 6046 1046 6118
rect 1109 6117 1121 6118
rect 1110 6047 1121 6117
rect 1109 6046 1121 6047
rect 1030 6030 1121 6046
rect 4172 6007 4258 6015
rect 4172 6003 4259 6007
rect 4172 5911 4177 6003
rect 4255 5911 4259 6003
rect 4172 5898 4259 5911
rect 1300 5577 1359 5589
rect 1300 5490 1302 5577
rect 1357 5490 1359 5577
rect 1300 5475 1359 5490
rect 3872 5437 3927 5450
rect 1621 5388 1681 5410
rect 1621 5300 1624 5388
rect 1678 5300 1681 5388
rect 3872 5345 3873 5437
rect 3925 5345 3927 5437
rect 3872 5332 3927 5345
rect 1621 5284 1681 5300
rect 3551 5260 3603 5274
rect 3551 5166 3603 5178
rect -492 5129 -339 5143
rect -492 5054 -465 5129
rect -362 5117 -339 5129
rect -362 5104 229 5117
rect -362 5054 120 5104
rect -492 5039 120 5054
rect 216 5039 229 5104
rect -492 5031 229 5039
rect -492 5029 -339 5031
rect 100 5029 229 5031
rect 1949 4928 2165 4938
rect 1949 4872 1975 4928
rect 2146 4872 2165 4928
rect 1949 4859 2165 4872
rect 2731 4931 2994 4943
rect 2731 4878 2775 4931
rect 2945 4878 2994 4931
rect 2731 4861 2994 4878
rect 7102 4923 7332 4939
rect 7102 4856 7125 4923
rect 7312 4856 7332 4923
rect 7102 4843 7332 4856
rect 14005 4880 14560 4882
rect 14005 4860 16220 4880
rect 914 4642 1862 4800
rect 2275 4638 2490 4803
rect 3229 4633 6524 4761
rect 7864 4599 8247 4761
rect 14005 4740 15680 4860
rect 16170 4740 16220 4860
rect 14005 4711 16220 4740
rect 15567 4710 16220 4711
rect 15567 4709 15649 4710
rect 1265 4514 1437 4528
rect 1265 4433 1281 4514
rect 1416 4433 1437 4514
rect 1530 4514 1702 4529
rect 1530 4475 1546 4514
rect 1265 4421 1437 4433
rect 1529 4433 1546 4475
rect 1682 4433 1702 4514
rect 1529 4419 1702 4433
rect 3467 4520 3639 4540
rect 3467 4439 3487 4520
rect 3622 4439 3639 4520
rect 3467 4424 3639 4439
rect 3823 4518 3995 4538
rect 3823 4437 3843 4518
rect 3978 4437 3995 4518
rect 3823 4422 3995 4437
rect 4189 4513 4343 4533
rect 4189 4435 4216 4513
rect 4327 4435 4343 4513
rect 4189 4420 4343 4435
rect 4564 4516 4718 4536
rect 4564 4438 4591 4516
rect 4702 4438 4718 4516
rect 4564 4422 4718 4438
rect 5079 4520 5252 4540
rect 5079 4439 5100 4520
rect 5235 4439 5252 4520
rect 5079 4424 5252 4439
rect 5812 4518 5985 4538
rect 5812 4437 5833 4518
rect 5968 4437 5985 4518
rect 5812 4422 5985 4437
rect 9269 4525 9442 4545
rect 9269 4444 9290 4525
rect 9425 4444 9442 4525
rect 9269 4428 9442 4444
rect 11436 4528 11609 4548
rect 11436 4447 11457 4528
rect 11592 4447 11609 4528
rect 11436 4431 11609 4447
rect 12896 4529 13069 4549
rect 12896 4448 12917 4529
rect 13052 4448 13069 4529
rect 12896 4432 13069 4448
rect 13799 4529 13971 4547
rect 13799 4448 13829 4529
rect 13952 4448 13971 4529
rect 13799 4429 13971 4448
rect 11965 4357 12096 4359
rect 11963 4348 12097 4357
rect 11962 4346 12097 4348
rect 11962 4267 11980 4346
rect 12084 4267 12097 4346
rect 11962 4177 12097 4267
rect 11634 4172 11765 4174
rect 11632 4163 11767 4172
rect 11631 4161 11767 4163
rect 11631 4082 11649 4161
rect 11753 4082 11767 4161
rect 11631 3991 11767 4082
rect 10701 3977 10834 3990
rect 10701 3898 10716 3977
rect 10820 3898 10834 3977
rect 10701 3855 10834 3898
rect 11631 3880 11766 3991
rect 10700 3812 10834 3855
rect 11630 3860 11766 3880
rect 9763 3810 9888 3811
rect 9760 3797 9893 3810
rect 9760 3718 9775 3797
rect 9879 3718 9893 3797
rect 8935 3621 9060 3635
rect 9760 3632 9893 3718
rect 8935 3542 8947 3621
rect 9051 3542 9060 3621
rect 8935 3458 9060 3542
rect 8599 3442 8731 3456
rect 8599 3363 8611 3442
rect 8715 3433 8731 3442
rect 8715 3363 8732 3433
rect 8154 3266 8286 3280
rect 8154 3187 8166 3266
rect 8270 3187 8286 3266
rect 8154 3105 8286 3187
rect 7857 3088 7983 3101
rect 7857 3075 7866 3088
rect 7855 3009 7866 3075
rect 7970 3075 7983 3088
rect 7970 3009 7984 3075
rect 6950 2908 7076 2922
rect 6950 2829 6959 2908
rect 7063 2829 7076 2908
rect 6950 2775 7076 2829
rect 6949 2746 7076 2775
rect 5990 2730 6116 2744
rect 5990 2651 5999 2730
rect 6103 2651 6116 2730
rect 5142 2568 5266 2571
rect 5139 2567 5266 2568
rect 5138 2554 5266 2567
rect 5138 2475 5150 2554
rect 5254 2475 5266 2554
rect 5138 2394 5266 2475
rect 4820 2390 4944 2391
rect 4819 2377 4944 2390
rect 4819 2298 4831 2377
rect 4935 2364 4944 2377
rect 4935 2298 4945 2364
rect 4389 2212 4513 2213
rect 4387 2199 4513 2212
rect 4387 2120 4400 2199
rect 4504 2120 4513 2199
rect 4387 2033 4513 2120
rect 4387 2031 4512 2033
rect 4049 2015 4173 2029
rect 4049 2005 4060 2015
rect 4048 1936 4060 2005
rect 4164 1936 4173 2015
rect 4048 1875 4173 1936
rect 3165 1801 3292 1814
rect 3165 1736 3179 1801
rect 3164 1723 3179 1736
rect 3279 1723 3292 1801
rect 2239 1620 2367 1633
rect 2239 1542 2254 1620
rect 2354 1542 2367 1620
rect 1600 1445 1722 1457
rect -649 1379 -278 1382
rect 140 1379 310 1380
rect -649 1196 310 1379
rect 1600 1360 1612 1445
rect 1713 1360 1722 1445
rect 1600 1280 1722 1360
rect -454 1194 310 1196
rect 140 1121 310 1194
rect 1351 1261 1473 1276
rect 1351 1181 1362 1261
rect 1461 1181 1473 1261
rect 1351 1171 1473 1181
rect 135 1108 320 1121
rect 135 1018 155 1108
rect 306 1018 320 1108
rect 135 1003 320 1018
rect 1017 1087 1140 1106
rect 1017 1015 1034 1087
rect 1122 1015 1140 1087
rect 1017 996 1140 1015
rect 1017 919 1033 996
rect 1123 919 1140 996
rect 1352 1004 1471 1171
rect 1352 986 1475 1004
rect 1352 977 1368 986
rect 501 899 707 916
rect 1017 905 1140 919
rect 1353 909 1368 977
rect 1458 909 1475 986
rect 501 897 524 899
rect 501 802 523 897
rect 689 806 707 899
rect 1353 895 1475 909
rect 1601 1003 1720 1280
rect 1601 985 1723 1003
rect 1601 908 1616 985
rect 1706 908 1723 985
rect 2239 986 2367 1542
rect 2239 929 2257 986
rect 1601 894 1723 908
rect 2242 909 2257 929
rect 2347 929 2367 986
rect 3164 1632 3292 1723
rect 3164 982 3288 1632
rect 3810 1442 3929 1457
rect 3810 1364 3828 1442
rect 3921 1364 3929 1442
rect 3810 994 3929 1364
rect 4048 999 4172 1875
rect 3166 977 3288 982
rect 2347 909 2364 929
rect 2242 895 2364 909
rect 3166 900 3181 977
rect 3271 900 3288 977
rect 3166 886 3288 900
rect 3807 976 3929 994
rect 3807 899 3822 976
rect 3912 899 3929 976
rect 3807 885 3929 899
rect 4047 981 4172 999
rect 4047 904 4062 981
rect 4152 952 4172 981
rect 4387 983 4510 2031
rect 4152 904 4169 952
rect 4047 890 4169 904
rect 4387 906 4402 983
rect 4492 916 4510 983
rect 4819 980 4945 2298
rect 5143 1006 5263 2394
rect 5390 1434 5509 1455
rect 5390 1361 5397 1434
rect 5501 1361 5509 1434
rect 4819 925 4838 980
rect 4492 906 4509 916
rect 4387 892 4509 906
rect 4823 903 4838 925
rect 4928 903 4945 980
rect 4823 889 4945 903
rect 5142 988 5264 1006
rect 5142 911 5157 988
rect 5247 911 5264 988
rect 5390 1005 5509 1361
rect 5390 987 5513 1005
rect 5390 930 5406 987
rect 5142 897 5264 911
rect 5391 910 5406 930
rect 5496 910 5513 987
rect 5990 991 6116 2651
rect 5990 966 6007 991
rect 5391 896 5513 910
rect 5992 914 6007 966
rect 6097 966 6116 991
rect 6949 985 7073 2746
rect 6097 914 6114 966
rect 5992 900 6114 914
rect 6949 908 6965 985
rect 7055 908 7073 985
rect 6949 894 7073 908
rect 7616 1453 7741 1464
rect 7616 1366 7631 1453
rect 7729 1366 7741 1453
rect 7616 971 7741 1366
rect 7616 894 7631 971
rect 7721 894 7741 971
rect 7616 879 7741 894
rect 7855 979 7984 3009
rect 7855 902 7872 979
rect 7962 902 7984 979
rect 7855 889 7984 902
rect 8155 3034 8285 3105
rect 8155 984 8284 3034
rect 8599 3010 8732 3363
rect 8935 3074 9061 3458
rect 8155 907 8176 984
rect 8266 907 8284 984
rect 8155 890 8284 907
rect 8601 978 8730 3010
rect 8601 901 8620 978
rect 8710 901 8730 978
rect 7857 888 7979 889
rect 8601 884 8730 901
rect 8934 981 9063 3074
rect 9761 3050 9893 3632
rect 8934 904 8953 981
rect 9043 904 9063 981
rect 8934 888 9063 904
rect 9156 1448 9283 1458
rect 9156 1362 9171 1448
rect 9273 1362 9283 1448
rect 9156 980 9283 1362
rect 9156 903 9171 980
rect 9261 903 9283 980
rect 9156 894 9283 903
rect 9762 979 9891 3050
rect 10700 3048 10833 3812
rect 11630 3089 11763 3860
rect 11628 3073 11763 3089
rect 9762 902 9781 979
rect 9871 902 9891 979
rect 9156 889 9278 894
rect 9762 888 9891 902
rect 10701 984 10830 3048
rect 10701 907 10719 984
rect 10809 907 10830 984
rect 10701 890 10830 907
rect 11395 1452 11522 1460
rect 11395 1361 11404 1452
rect 11514 1361 11522 1452
rect 11395 989 11522 1361
rect 11395 912 11411 989
rect 11501 912 11522 989
rect 11395 898 11522 912
rect 11628 997 11757 3073
rect 11628 920 11648 997
rect 11738 920 11757 997
rect 11628 903 11757 920
rect 11968 986 12091 4177
rect 11968 909 11984 986
rect 12074 909 12091 986
rect 11968 897 12091 909
rect 11969 895 12091 897
rect 687 802 707 806
rect 501 790 707 802
rect 2725 668 2806 749
rect 4602 669 4728 751
rect 6530 669 6656 751
rect 8396 671 8527 749
rect 10306 670 10565 752
rect 12207 750 14560 753
rect 15567 750 16209 751
rect 12207 739 16209 750
rect 12207 682 15685 739
rect 16183 682 16209 739
rect 12207 670 16209 682
rect 15567 668 16209 670
rect 15650 667 16208 668
rect 1045 541 1123 554
rect 1045 457 1053 541
rect 1120 457 1123 541
rect 1045 437 1123 457
rect 1364 531 1449 545
rect 1364 463 1375 531
rect 1443 463 1449 531
rect 1364 448 1449 463
rect 1749 449 1759 451
rect 1703 441 1759 449
rect 1703 439 1761 441
rect 1703 379 1704 439
rect 1756 379 1761 439
rect 1703 375 1761 379
rect 1705 367 1761 375
rect 3762 436 3824 448
rect 3762 376 3769 436
rect 3821 376 3824 436
rect 5493 440 5564 450
rect 5493 436 5571 440
rect 3762 363 3824 376
rect 4073 415 4163 431
rect 4073 353 4088 415
rect 4150 353 4163 415
rect 4849 410 4934 421
rect 4073 339 4163 353
rect 4396 401 4480 410
rect 4396 340 4404 401
rect 4471 340 4480 401
rect 4396 332 4480 340
rect 4849 353 4862 410
rect 4924 353 4934 410
rect 4849 339 4934 353
rect 5165 420 5257 433
rect 5165 359 5180 420
rect 5245 359 5257 420
rect 5493 377 5506 436
rect 5558 377 5571 436
rect 5493 371 5571 377
rect 7551 436 7630 441
rect 7551 376 7565 436
rect 7617 376 7630 436
rect 9280 435 9357 441
rect 11350 440 11429 450
rect 7551 371 7630 376
rect 7862 416 7950 428
rect 8183 422 8276 428
rect 5552 365 5564 371
rect 5165 348 5257 359
rect 7862 364 7877 416
rect 7935 364 7950 416
rect 7862 350 7950 364
rect 8182 415 8276 422
rect 8182 353 8199 415
rect 8264 353 8276 415
rect 8955 412 9040 424
rect 8182 346 8276 353
rect 8183 341 8276 346
rect 8636 400 8719 410
rect 8636 339 8646 400
rect 8711 339 8719 400
rect 8955 354 8970 412
rect 9030 354 9040 412
rect 9280 378 9292 435
rect 9345 378 9357 435
rect 9280 371 9357 378
rect 11349 437 11429 440
rect 11349 375 11358 437
rect 11421 375 11429 437
rect 11349 370 11429 375
rect 11350 359 11429 370
rect 11663 415 11752 425
rect 11663 359 11678 415
rect 11740 359 11752 415
rect 8955 345 9040 354
rect 11663 347 11752 359
rect 11982 408 12073 419
rect 8636 326 8719 339
rect 11982 344 11994 408
rect 12061 344 12073 408
rect 11982 334 12073 344
rect 773 30 914 112
rect 2642 29 2890 110
rect 4627 33 4717 112
rect 6432 33 6680 114
rect 8412 30 8493 113
rect 10237 31 10496 113
rect 12201 110 14560 112
rect 16407 110 16967 113
rect 12201 100 16967 110
rect 12201 43 16481 100
rect 16942 43 16967 100
rect 12201 30 16967 43
rect 15567 28 16967 30
rect 16407 26 16967 28
<< via1 >>
rect 15719 10475 16169 10570
rect 1189 10202 1425 10299
rect 1425 10202 1426 10299
rect 2801 10206 3040 10300
rect 5639 10196 5889 10305
rect 9805 10198 10045 10300
rect 13913 10189 14146 10280
rect -479 10049 -348 10113
rect 677 10051 779 10109
rect 16480 8246 16937 8349
rect 16496 6678 16910 6773
rect 956 6285 1030 6361
rect 1046 6117 1109 6118
rect 1046 6047 1109 6117
rect 1046 6046 1109 6047
rect 4177 5911 4255 6003
rect 1302 5490 1357 5577
rect 1624 5300 1678 5388
rect 3873 5345 3925 5437
rect 3551 5178 3603 5260
rect -465 5054 -362 5129
rect 120 5039 216 5104
rect 1975 4872 2146 4928
rect 2775 4878 2945 4931
rect 7125 4856 7312 4923
rect 15680 4740 16170 4860
rect 1281 4433 1416 4514
rect 1546 4433 1681 4514
rect 3487 4439 3622 4520
rect 3843 4437 3978 4518
rect 4216 4435 4327 4513
rect 4591 4438 4702 4516
rect 5100 4439 5235 4520
rect 5833 4437 5968 4518
rect 9290 4444 9425 4525
rect 11457 4447 11592 4528
rect 12917 4448 13052 4529
rect 13829 4448 13952 4529
rect 11980 4267 12084 4346
rect 11649 4082 11753 4161
rect 10716 3898 10820 3977
rect 9775 3718 9879 3797
rect 8947 3542 9051 3621
rect 8611 3363 8715 3442
rect 8166 3187 8270 3266
rect 7866 3009 7970 3088
rect 6959 2829 7063 2908
rect 5999 2651 6103 2730
rect 5150 2475 5254 2554
rect 4831 2298 4935 2377
rect 4400 2120 4504 2199
rect 4060 1936 4164 2015
rect 3179 1723 3279 1801
rect 2254 1542 2354 1620
rect 1612 1360 1713 1445
rect 1362 1181 1461 1261
rect 1034 1015 1122 1087
rect 275 799 335 908
rect 523 806 524 897
rect 524 806 687 897
rect 3828 1364 3921 1442
rect 5397 1361 5501 1434
rect 7631 1366 7729 1453
rect 9171 1362 9273 1448
rect 11404 1361 11514 1452
rect 523 802 687 806
rect 15685 682 16183 739
rect 649 537 714 630
rect 1053 457 1120 541
rect 1375 463 1443 531
rect 1704 379 1756 439
rect 3769 376 3821 436
rect 4088 353 4150 415
rect 4404 340 4471 401
rect 4862 353 4924 410
rect 5180 359 5245 420
rect 5506 377 5558 436
rect 7565 376 7617 436
rect 7877 364 7935 416
rect 8199 353 8264 415
rect 8646 339 8711 400
rect 8970 354 9030 412
rect 9292 378 9345 435
rect 11358 375 11421 437
rect 11678 359 11740 415
rect 11994 344 12061 408
rect 16481 43 16942 100
<< metal2 >>
rect -492 10113 -341 10580
rect -492 10049 -479 10113
rect -348 10049 -341 10113
rect -492 5129 -341 10049
rect -223 10005 -44 10580
rect -224 9961 -44 10005
rect 79 10009 259 10581
rect 79 9976 260 10009
rect 355 9976 538 10583
rect 1187 10319 1424 10321
rect 1167 10299 1450 10319
rect 2800 10317 3040 10767
rect 1167 10202 1189 10299
rect 1426 10292 1450 10299
rect 1427 10204 1450 10292
rect 1426 10202 1450 10204
rect 1167 10190 1450 10202
rect 2779 10300 3057 10317
rect 5640 10313 5879 10745
rect 9823 10316 10033 10820
rect 2779 10206 2801 10300
rect 3040 10206 3057 10300
rect 2779 10194 3057 10206
rect 5623 10305 5897 10313
rect 5623 10196 5639 10305
rect 5889 10196 5897 10305
rect 5623 10184 5897 10196
rect 9791 10300 10056 10316
rect 9791 10198 9805 10300
rect 10045 10198 10056 10300
rect 13899 10296 14145 10800
rect 15652 10570 16218 10593
rect 15652 10475 15719 10570
rect 16169 10475 16218 10570
rect 15652 10426 16218 10475
rect 9791 10189 10056 10198
rect 13880 10280 14168 10296
rect 13880 10189 13913 10280
rect 14146 10189 14168 10280
rect 13880 10172 14168 10189
rect 934 10120 7288 10123
rect 643 10109 7288 10120
rect 643 10051 677 10109
rect 779 10051 7288 10109
rect 643 10044 7288 10051
rect 13142 10047 13291 10073
rect 643 10041 6997 10044
rect 12688 10030 13341 10047
rect -224 9883 -202 9961
rect -65 9883 -44 9961
rect -224 9857 -44 9883
rect 80 9870 260 9976
rect 357 9870 537 9976
rect 4400 9964 4520 9980
rect 12686 9973 13341 10030
rect 4400 9889 4408 9964
rect 4490 9889 4520 9964
rect 4400 9870 4520 9889
rect 7000 9950 13341 9973
rect 7000 9870 13340 9950
rect -223 5606 -44 9857
rect 79 9861 260 9870
rect 79 9777 259 9861
rect 79 9681 107 9777
rect 245 9681 259 9777
rect 79 8050 259 9681
rect 355 9446 538 9870
rect 13219 9869 13340 9870
rect 1700 9765 1810 9790
rect 1700 9681 1715 9765
rect 1787 9681 1810 9765
rect 1700 9660 1810 9681
rect 355 9310 1075 9446
rect 79 5927 261 8050
rect 355 6001 538 9310
rect 8939 8098 9075 8592
rect 13021 8501 13143 8530
rect 8939 8009 8955 8098
rect 9055 8009 9075 8098
rect 8939 7989 9075 8009
rect 8939 7896 9072 7909
rect 8939 7794 8950 7896
rect 9067 7794 9072 7896
rect 5549 7632 5678 7659
rect 8939 7654 9072 7794
rect 5549 7540 5570 7632
rect 5667 7540 5678 7632
rect 5549 7518 5678 7540
rect 3241 7381 3361 7402
rect 3241 7293 3251 7381
rect 3340 7293 3361 7381
rect 1735 7134 1855 7154
rect 1735 7042 1745 7134
rect 1846 7042 1855 7134
rect 1735 6521 1855 7042
rect 3241 7031 3361 7293
rect 3241 6938 3363 7031
rect 3243 6543 3363 6938
rect 4402 6457 4428 6549
rect 4515 6457 4639 6552
rect 5549 6551 5679 7518
rect 8942 6573 9071 7654
rect 13020 6958 13143 8501
rect 16410 8349 16960 8371
rect 16410 8246 16480 8349
rect 16937 8246 16960 8349
rect 16410 8209 16960 8246
rect 12988 6929 13214 6958
rect 12988 6849 13018 6929
rect 13177 6849 13214 6929
rect 12988 6839 13214 6849
rect 16414 6773 16966 6812
rect 16414 6678 16496 6773
rect 16910 6678 16966 6773
rect 16414 6639 16966 6678
rect 5551 6539 5663 6551
rect 4425 6442 4428 6457
rect 906 6376 1033 6377
rect 870 6361 1033 6376
rect 870 6285 956 6361
rect 1030 6285 1033 6361
rect 870 6271 1033 6285
rect 870 6270 949 6271
rect -223 5394 -43 5606
rect 79 5593 263 5927
rect 355 5905 371 6001
rect 507 5905 538 6001
rect 355 5786 538 5905
rect 871 5786 947 6270
rect 1030 6118 1121 6150
rect 1030 6046 1046 6118
rect 1109 6046 1121 6118
rect 1030 6030 1121 6046
rect 354 5780 947 5786
rect 3394 6010 3510 6012
rect 4165 6010 4758 6014
rect 3394 6003 4758 6010
rect 3394 5911 4177 6003
rect 4255 5911 4758 6003
rect 3394 5906 4758 5911
rect 3394 5901 4294 5906
rect 3394 5781 3510 5901
rect 2761 5780 3513 5781
rect 354 5662 3513 5780
rect 354 5661 2774 5662
rect 354 5658 886 5661
rect 4666 5637 4755 5906
rect 1317 5595 1758 5596
rect 924 5594 1758 5595
rect 2072 5594 2424 5595
rect 353 5593 2424 5594
rect 2587 5593 3543 5594
rect 77 5582 3543 5593
rect 77 5479 534 5582
rect 673 5577 3543 5582
rect 673 5490 1302 5577
rect 1357 5490 3543 5577
rect 4664 5515 13974 5637
rect 673 5479 3543 5490
rect 77 5474 3543 5479
rect 77 5473 2885 5474
rect 77 5472 1365 5473
rect 1668 5472 2687 5473
rect 77 5471 1274 5472
rect 1668 5471 2424 5472
rect 79 5469 263 5471
rect 353 5469 852 5471
rect 3423 5446 3543 5474
rect 3423 5437 4929 5446
rect -225 5393 454 5394
rect 1073 5393 1755 5394
rect 2408 5393 3314 5394
rect -225 5392 3314 5393
rect -225 5388 3353 5392
rect -225 5300 1624 5388
rect 1678 5300 3353 5388
rect 3423 5345 3873 5437
rect 3925 5345 4929 5437
rect 3423 5341 4929 5345
rect 5511 5427 11740 5446
rect 5511 5360 11577 5427
rect 11675 5360 11740 5427
rect 5511 5342 11740 5360
rect 3610 5340 4929 5341
rect -225 5297 3353 5300
rect -225 5296 1511 5297
rect 1749 5296 2431 5297
rect -225 5295 865 5296
rect -225 5289 454 5295
rect -492 5054 -465 5129
rect -362 5054 -341 5129
rect -492 5028 -341 5054
rect -492 4063 -342 5028
rect -494 3004 -342 4063
rect -494 2875 -344 3004
rect -494 1777 -339 2875
rect -490 888 -339 1777
rect -491 873 -339 888
rect -491 799 -480 873
rect -353 799 -339 873
rect -221 897 -68 5289
rect 3263 5269 3353 5297
rect 4792 5271 5697 5272
rect 11292 5271 12790 5272
rect 4120 5269 5697 5271
rect 3263 5260 5697 5269
rect 3263 5178 3551 5260
rect 3603 5178 5697 5260
rect 3263 5172 5697 5178
rect 3263 5171 5025 5172
rect 6270 5171 12794 5271
rect 3334 5169 4239 5171
rect 11292 5170 12794 5171
rect 99 5104 1954 5110
rect 99 5039 120 5104
rect 216 5039 1954 5104
rect 99 5028 1954 5039
rect 2240 5025 2514 5108
rect 4982 5100 7761 5101
rect 3054 5052 7761 5100
rect 7807 5052 8147 5053
rect 3054 5013 8147 5052
rect 3054 5012 5833 5013
rect 7736 4987 8147 5013
rect 10692 4987 10705 5053
rect 10871 4987 11032 5053
rect 12690 5049 12794 5170
rect 13846 5031 13971 5515
rect 7736 4986 8076 4987
rect 1949 4928 2165 4938
rect 1949 4872 1975 4928
rect 2146 4872 2165 4928
rect 1949 4858 2165 4872
rect 2731 4934 2994 4943
rect 2731 4878 2775 4934
rect 2945 4878 2994 4934
rect 2731 4861 2994 4878
rect 7102 4923 7332 4939
rect 7102 4856 7125 4923
rect 7312 4856 7332 4923
rect 7102 4843 7332 4856
rect 15650 4860 16220 4880
rect 15650 4740 15680 4860
rect 16170 4740 16220 4860
rect 15650 4710 16220 4740
rect 1019 4532 1126 4535
rect 1019 4521 1128 4532
rect 1019 4439 1035 4521
rect 1117 4439 1128 4521
rect 1019 1460 1128 4439
rect 1265 4514 1437 4528
rect 1265 4433 1281 4514
rect 1416 4433 1437 4514
rect 1530 4514 1702 4529
rect 1530 4475 1546 4514
rect 1265 4421 1437 4433
rect 1529 4433 1546 4475
rect 1681 4433 1702 4514
rect 1529 4419 1702 4433
rect 3467 4520 3639 4540
rect 3467 4439 3487 4520
rect 3622 4439 3639 4520
rect 3467 4424 3639 4439
rect 3823 4518 3995 4538
rect 3823 4437 3843 4518
rect 3978 4437 3995 4518
rect 3823 4422 3995 4437
rect 4189 4513 4343 4533
rect 4189 4435 4216 4513
rect 4327 4435 4343 4513
rect 4189 4420 4343 4435
rect 4564 4516 4718 4536
rect 4564 4438 4591 4516
rect 4702 4438 4718 4516
rect 4564 4422 4718 4438
rect 5079 4520 5252 4540
rect 5079 4439 5100 4520
rect 5235 4439 5252 4520
rect 5079 4424 5252 4439
rect 5812 4518 5985 4538
rect 5812 4437 5833 4518
rect 5968 4437 5985 4518
rect 5812 4422 5985 4437
rect 9269 4525 9442 4545
rect 9269 4444 9290 4525
rect 9425 4444 9442 4525
rect 9269 4428 9442 4444
rect 11436 4528 11609 4548
rect 11436 4447 11457 4528
rect 11592 4447 11609 4528
rect 11436 4431 11609 4447
rect 12896 4529 13069 4549
rect 12896 4448 12917 4529
rect 13052 4448 13069 4529
rect 12896 4432 13069 4448
rect 13799 4529 13971 4547
rect 13799 4448 13829 4529
rect 13952 4448 13971 4529
rect 13799 4429 13971 4448
rect 11962 4359 12166 4360
rect 11962 4346 14177 4359
rect 11962 4267 11980 4346
rect 12084 4267 14177 4346
rect 11962 4241 14177 4267
rect 12751 4178 14175 4181
rect 12368 4175 14175 4178
rect 11882 4174 14175 4175
rect 11635 4161 14175 4174
rect 11635 4082 11649 4161
rect 11753 4082 14175 4161
rect 11635 4061 14175 4082
rect 11635 4059 12390 4061
rect 11751 4058 12390 4059
rect 12751 4060 14175 4061
rect 12751 4058 13329 4060
rect 11751 4057 11893 4058
rect 12265 3991 13326 3993
rect 10819 3990 13326 3991
rect 10702 3989 13326 3990
rect 10702 3977 14166 3989
rect 10702 3898 10716 3977
rect 10820 3898 14166 3977
rect 10702 3876 14166 3898
rect 10702 3875 12290 3876
rect 12749 3875 14166 3876
rect 10819 3874 12290 3875
rect 13311 3873 14166 3875
rect 12746 3812 13323 3813
rect 9761 3797 14180 3812
rect 9761 3718 9775 3797
rect 9879 3718 14180 3797
rect 9761 3695 14180 3718
rect 13304 3694 14180 3695
rect 9060 3635 9207 3636
rect 8936 3632 9376 3635
rect 12743 3633 13320 3636
rect 12743 3632 14160 3633
rect 8936 3621 14160 3632
rect 8936 3542 8947 3621
rect 9051 3542 14160 3621
rect 8936 3519 14160 3542
rect 9060 3518 9176 3519
rect 9316 3518 14160 3519
rect 13305 3517 14160 3518
rect 13303 3457 14151 3460
rect 8600 3453 9244 3456
rect 12733 3453 14151 3457
rect 8600 3442 14151 3453
rect 8600 3363 8611 3442
rect 8715 3363 14151 3442
rect 8600 3340 14151 3363
rect 9240 3339 14151 3340
rect 13299 3282 14147 3283
rect 8761 3281 8976 3282
rect 8272 3279 9243 3281
rect 12732 3279 14147 3282
rect 8158 3266 14147 3279
rect 8158 3187 8166 3266
rect 8270 3187 14147 3266
rect 8158 3169 14147 3187
rect 8172 3168 14147 3169
rect 8251 3167 14147 3168
rect 8272 3166 14147 3167
rect 9235 3165 14147 3166
rect 12732 3164 14147 3165
rect 8982 3103 9252 3104
rect 12731 3103 14151 3107
rect 7985 3101 14151 3103
rect 7858 3088 14151 3101
rect 7858 3009 7866 3088
rect 7970 3009 14151 3088
rect 7858 2991 14151 3009
rect 7872 2990 14151 2991
rect 7951 2989 14151 2990
rect 7985 2986 9252 2989
rect 12732 2925 14147 2928
rect 7159 2922 14147 2925
rect 6951 2908 14147 2922
rect 6951 2829 6959 2908
rect 7063 2829 14147 2908
rect 6951 2811 14147 2829
rect 6965 2810 9062 2811
rect 12732 2810 14147 2811
rect 7044 2809 7215 2810
rect 6105 2744 9528 2746
rect 5991 2743 9528 2744
rect 12730 2743 14147 2748
rect 5991 2730 14147 2743
rect 5991 2651 5999 2730
rect 6103 2651 14147 2730
rect 5991 2633 14147 2651
rect 6005 2632 14147 2633
rect 6084 2631 14147 2632
rect 6116 2630 6172 2631
rect 9299 2630 14147 2631
rect 9299 2629 13266 2630
rect 5139 2554 14145 2568
rect 5139 2475 5150 2554
rect 5254 2475 14145 2554
rect 5139 2457 14145 2475
rect 5156 2456 14145 2457
rect 5235 2455 5640 2456
rect 5366 2392 13277 2393
rect 4928 2391 13277 2392
rect 4820 2377 14144 2391
rect 4820 2298 4831 2377
rect 4935 2298 14144 2377
rect 4820 2281 14144 2298
rect 4820 2280 5726 2281
rect 4837 2279 5726 2280
rect 13261 2279 14144 2281
rect 4406 2214 4513 2215
rect 4406 2213 13280 2214
rect 4389 2199 14143 2213
rect 4389 2120 4400 2199
rect 4504 2120 14143 2199
rect 4389 2102 14143 2120
rect 4406 2101 5832 2102
rect 13260 2101 14143 2102
rect 4389 2031 4513 2034
rect 4066 2030 5671 2031
rect 4066 2029 14143 2030
rect 4049 2015 14143 2029
rect 4049 1936 4060 2015
rect 4164 1936 14143 2015
rect 4049 1918 14143 1936
rect 4066 1917 5671 1918
rect 3809 1817 3966 1822
rect 3168 1816 4711 1817
rect 3168 1814 14149 1816
rect 3165 1801 14149 1814
rect 3165 1723 3179 1801
rect 3279 1723 14149 1801
rect 3165 1709 14149 1723
rect 3165 1708 3809 1709
rect 3168 1707 3809 1708
rect 3938 1707 14149 1709
rect 4699 1706 14149 1707
rect 5422 1704 14149 1706
rect 3800 1638 3957 1644
rect 5463 1638 7006 1641
rect 13263 1638 14146 1641
rect 2237 1633 2480 1635
rect 3165 1634 3293 1636
rect 3800 1634 14146 1638
rect 3165 1633 14146 1634
rect 2237 1620 14146 1633
rect 2237 1542 2254 1620
rect 2354 1542 14146 1620
rect 2237 1531 14146 1542
rect 2237 1528 3809 1531
rect 3938 1528 5464 1531
rect 6628 1529 14146 1531
rect 2237 1527 3207 1528
rect 1019 1457 1656 1460
rect 6929 1459 12502 1461
rect 13265 1459 14148 1461
rect 5390 1458 14148 1459
rect 3938 1457 14148 1458
rect 1019 1455 1916 1457
rect 3849 1455 14148 1457
rect 1019 1453 14148 1455
rect 1019 1445 7631 1453
rect 1019 1360 1612 1445
rect 1713 1442 7631 1445
rect 1713 1364 3828 1442
rect 3921 1434 7631 1442
rect 3921 1364 5397 1434
rect 1713 1361 5397 1364
rect 5501 1366 7631 1434
rect 7729 1452 14148 1453
rect 7729 1448 11404 1452
rect 7729 1366 9171 1448
rect 5501 1362 9171 1366
rect 9273 1362 11404 1448
rect 5501 1361 11404 1362
rect 11514 1361 14148 1452
rect 1713 1360 14148 1361
rect 1019 1350 14148 1360
rect 1019 1349 12502 1350
rect 13265 1349 14148 1350
rect 1019 1348 3127 1349
rect 3849 1348 5392 1349
rect 1019 1347 1916 1348
rect 1019 1346 1656 1347
rect 1019 1315 1195 1346
rect 509 1182 1195 1315
rect 5097 1285 6640 1286
rect 13258 1285 14141 1286
rect 265 908 338 921
rect 265 897 275 908
rect -221 800 275 897
rect -491 780 -339 799
rect 265 799 275 800
rect 335 799 338 908
rect 265 783 338 799
rect 513 897 697 1182
rect 1070 1181 1195 1182
rect 1351 1277 1667 1278
rect 1351 1276 2184 1277
rect 3556 1276 14141 1285
rect 1351 1261 14141 1276
rect 1351 1181 1362 1261
rect 1461 1181 14141 1261
rect 1351 1176 14141 1181
rect 1351 1175 5099 1176
rect 1351 1171 3571 1175
rect 13258 1174 14141 1176
rect 1476 1170 3571 1171
rect 2138 1169 2846 1170
rect 1016 1103 1167 1106
rect 1016 1101 13327 1103
rect 1016 1087 14145 1101
rect 1016 1015 1034 1087
rect 1122 1015 14145 1087
rect 1016 1009 14145 1015
rect 513 802 523 897
rect 687 802 697 897
rect 513 786 697 802
rect 1811 883 1951 897
rect 1811 807 1841 883
rect 1912 830 1951 883
rect 11929 833 12418 834
rect 11929 830 12423 833
rect 1912 807 12423 830
rect -490 775 -339 780
rect 1811 762 12423 807
rect 11929 760 12423 762
rect 636 641 720 644
rect -221 630 720 641
rect -221 621 649 630
rect -221 539 -211 621
rect -89 539 649 621
rect -221 537 649 539
rect 714 537 720 630
rect -221 529 720 537
rect 636 524 720 529
rect 1045 541 1126 554
rect 298 -67 394 399
rect 643 358 719 524
rect 1045 457 1053 541
rect 1120 540 1126 541
rect 1123 457 1126 540
rect 1045 439 1126 457
rect 1364 531 1449 545
rect 1364 530 1375 531
rect 1364 462 1374 530
rect 1443 463 1449 531
rect 2647 500 2960 570
rect 3585 500 5830 571
rect 6441 501 6736 569
rect 7373 499 9618 570
rect 10234 502 10528 568
rect 12341 566 12423 760
rect 15650 739 16208 750
rect 15650 682 15685 739
rect 16183 682 16208 739
rect 15650 667 16208 682
rect 11171 499 12423 566
rect 12341 497 12423 499
rect 1442 462 1449 463
rect 1364 448 1449 462
rect 1690 439 1845 445
rect 5564 440 7631 441
rect 1690 379 1704 439
rect 1756 438 1845 439
rect 1756 436 3835 438
rect 1756 435 3769 436
rect 3821 435 3835 436
rect 1756 379 3768 435
rect 1690 377 3768 379
rect 3825 377 3835 435
rect 5483 436 7631 440
rect 1690 376 3769 377
rect 3821 376 3835 377
rect 1690 372 3835 376
rect 4073 415 4163 431
rect 1690 371 3833 372
rect 1690 369 1845 371
rect 1690 359 1770 369
rect 877 358 1770 359
rect 643 299 1770 358
rect 4073 353 4088 415
rect 4150 353 4163 415
rect 4849 410 4934 421
rect 4073 339 4163 353
rect 4396 401 4482 410
rect 4396 340 4404 401
rect 4472 340 4482 401
rect 4396 331 4482 340
rect 4849 353 4862 410
rect 4924 353 4934 410
rect 4849 339 4934 353
rect 5165 420 5257 433
rect 5165 359 5180 420
rect 5245 359 5257 420
rect 5483 377 5505 436
rect 5562 377 7564 436
rect 7620 377 7631 436
rect 9270 437 11436 441
rect 9270 435 11358 437
rect 5483 376 7565 377
rect 7617 376 7631 377
rect 5483 371 7631 376
rect 7862 420 7950 428
rect 5165 348 5257 359
rect 7862 364 7877 420
rect 7935 364 7950 420
rect 7862 350 7950 364
rect 8183 415 8276 428
rect 8183 353 8199 415
rect 8264 353 8276 415
rect 8955 412 9040 424
rect 8183 341 8276 353
rect 8636 400 8719 410
rect 8636 339 8646 400
rect 8711 339 8719 400
rect 8955 354 8970 412
rect 9030 354 9040 412
rect 9270 377 9292 435
rect 9348 377 11358 435
rect 9270 375 11358 377
rect 11421 375 11436 437
rect 9270 371 11436 375
rect 11663 415 11752 425
rect 8955 345 9040 354
rect 11663 359 11678 415
rect 11740 359 11752 415
rect 11663 347 11752 359
rect 11982 408 12073 419
rect 8636 326 8719 339
rect 11982 344 11994 408
rect 12061 344 12073 408
rect 11982 334 12073 344
rect 643 298 972 299
rect 1767 -39 1836 213
rect 298 -138 312 -67
rect 381 -138 394 -67
rect 298 -149 394 -138
rect 1766 -151 1836 -39
rect 1766 -273 1835 -151
rect 1766 -354 1775 -273
rect 1832 -354 1835 -273
rect 1766 -364 1835 -354
rect 3662 -459 3731 216
rect 3660 -468 3731 -459
rect 3660 -540 3672 -468
rect 3729 -540 3731 -468
rect 3660 -550 3731 -540
rect 5558 -670 5633 195
rect 5558 -671 5570 -670
rect 5558 -730 5567 -671
rect 5626 -702 5633 -670
rect 5558 -731 5570 -730
rect 5626 -731 5632 -702
rect 5558 -737 5632 -731
rect 7466 -739 7549 219
rect 7466 -855 7551 -739
rect 7466 -919 7478 -855
rect 7543 -919 7551 -855
rect 7466 -927 7551 -919
rect 9302 -931 9412 200
rect 9301 -1035 9412 -931
rect 9301 -1107 9320 -1035
rect 9391 -1054 9412 -1035
rect 9391 -1107 9410 -1054
rect 9301 -1123 9410 -1107
rect 11181 -1238 11269 188
rect 16407 100 16967 113
rect 16407 43 16481 100
rect 16942 43 16967 100
rect 16407 26 16967 43
rect 11181 -1307 11193 -1238
rect 11257 -1248 11269 -1238
rect 11257 -1307 11268 -1248
rect 11181 -1315 11268 -1307
<< via2 >>
rect 1191 10204 1426 10292
rect 1426 10204 1427 10292
rect 15719 10475 16169 10570
rect -202 9883 -65 9961
rect 4408 9889 4490 9964
rect 107 9681 245 9777
rect 1715 9681 1787 9765
rect 8955 8009 9055 8098
rect 8950 7794 9067 7896
rect 5570 7540 5667 7632
rect 3251 7293 3340 7381
rect 1745 7042 1846 7134
rect 16480 8246 16937 8349
rect 13018 6849 13177 6929
rect 16496 6678 16910 6773
rect 371 5905 507 6001
rect 1046 6046 1109 6118
rect 534 5479 673 5582
rect 11577 5360 11675 5427
rect -480 799 -353 873
rect 11583 4990 11694 5046
rect 1975 4872 2146 4928
rect 2775 4931 2945 4934
rect 2775 4878 2945 4931
rect 7125 4856 7312 4923
rect 15680 4740 16170 4860
rect 1035 4439 1117 4521
rect 1281 4433 1416 4514
rect 1546 4433 1681 4514
rect 3487 4439 3622 4520
rect 3843 4437 3978 4518
rect 4216 4435 4327 4513
rect 4591 4438 4702 4516
rect 5100 4439 5235 4520
rect 5833 4437 5968 4518
rect 9290 4444 9425 4525
rect 11457 4447 11592 4528
rect 12917 4448 13052 4529
rect 13829 4448 13952 4529
rect 275 800 335 904
rect 1841 807 1912 883
rect -211 539 -89 621
rect 1054 457 1120 540
rect 1120 457 1123 540
rect 1374 463 1375 530
rect 1375 463 1442 530
rect 15685 682 16183 739
rect 1374 462 1442 463
rect 3768 377 3769 435
rect 3769 377 3821 435
rect 3821 377 3825 435
rect 4088 353 4150 415
rect 4405 340 4471 401
rect 4471 340 4472 401
rect 4862 353 4924 410
rect 5180 359 5245 420
rect 5505 377 5506 436
rect 5506 377 5558 436
rect 5558 377 5562 436
rect 7564 377 7565 436
rect 7565 377 7617 436
rect 7617 377 7620 436
rect 7877 416 7935 420
rect 7877 364 7935 416
rect 8200 353 8264 415
rect 8646 339 8711 400
rect 8970 354 9030 412
rect 9292 378 9345 435
rect 9345 378 9348 435
rect 9292 377 9348 378
rect 11678 359 11740 415
rect 11994 344 12061 408
rect 312 -138 381 -67
rect 1775 -354 1832 -273
rect 3672 -540 3729 -468
rect 5570 -671 5626 -670
rect 5567 -730 5626 -671
rect 5570 -731 5626 -730
rect 7478 -919 7543 -855
rect 9320 -1107 9391 -1035
rect 16481 43 16942 100
rect 11193 -1307 11257 -1238
<< metal3 >>
rect 15652 10570 16218 10593
rect 15652 10475 15719 10570
rect 16169 10475 16218 10570
rect 15652 10426 16218 10475
rect 1166 10293 1450 10318
rect 1166 10292 1192 10293
rect 1423 10292 1450 10293
rect 1166 10204 1191 10292
rect 1427 10204 1450 10292
rect 1166 10201 1192 10204
rect 1423 10201 1450 10204
rect 1166 10187 1450 10201
rect 601 9976 696 9977
rect 4401 9976 4500 9977
rect -227 9964 4500 9976
rect -227 9961 4408 9964
rect -227 9883 -202 9961
rect -65 9889 4408 9961
rect 4490 9889 4500 9964
rect -65 9883 4500 9889
rect -227 9873 4500 9883
rect -227 9870 3565 9873
rect 601 9868 696 9870
rect 80 9777 1808 9791
rect 80 9681 107 9777
rect 245 9765 1808 9777
rect 245 9681 1715 9765
rect 1787 9681 1808 9765
rect 80 9653 1808 9681
rect 16410 8349 16960 8371
rect 16410 8246 16480 8349
rect 16937 8246 16960 8349
rect 16410 8209 16960 8246
rect 8937 8117 9517 8118
rect 8937 8098 14116 8117
rect 8937 8009 8955 8098
rect 9055 8009 14116 8098
rect 8937 7989 14116 8009
rect 8936 7896 14107 7907
rect 8936 7794 8950 7896
rect 9067 7794 14107 7896
rect 8936 7779 14107 7794
rect 5552 7656 5878 7657
rect 8937 7656 14108 7657
rect 5551 7632 14108 7656
rect 5551 7540 5570 7632
rect 5667 7540 14108 7632
rect 5551 7529 14108 7540
rect 5551 7526 14107 7529
rect 3241 7381 14103 7407
rect 3241 7293 3251 7381
rect 3340 7293 14103 7381
rect 3241 7281 14103 7293
rect 3241 7277 3574 7281
rect 1732 7155 2287 7156
rect 3239 7155 14101 7156
rect 1732 7134 14101 7155
rect 1732 7042 1745 7134
rect 1846 7042 14101 7134
rect 1732 7030 14101 7042
rect 1732 7029 12278 7030
rect 12988 6959 13405 6960
rect 12988 6929 14103 6959
rect 12988 6849 13018 6929
rect 13177 6849 14103 6929
rect 12988 6839 14103 6849
rect 16414 6773 16966 6812
rect 16414 6678 16496 6773
rect 16910 6678 16966 6773
rect 16414 6639 16966 6678
rect 1030 6148 1121 6150
rect 1020 6118 1125 6148
rect 1020 6117 1046 6118
rect 1109 6117 1125 6118
rect 1020 6048 1045 6117
rect 1111 6048 1125 6117
rect 1020 6046 1046 6048
rect 1109 6046 1125 6048
rect -221 6038 -75 6041
rect -221 6001 538 6038
rect -221 5905 371 6001
rect 507 5905 538 6001
rect -221 5893 538 5905
rect -491 873 -339 888
rect -491 799 -480 873
rect -353 799 -339 873
rect -491 780 -339 799
rect -221 621 -75 5893
rect 523 5582 684 5590
rect 523 5479 534 5582
rect 673 5479 684 5582
rect -221 539 -211 621
rect -89 539 -75 621
rect -221 526 -75 539
rect 262 904 350 926
rect 262 800 275 904
rect 335 800 350 904
rect 262 552 350 800
rect 523 823 684 5479
rect 1020 4522 1125 6046
rect 11560 5427 11704 5458
rect 11560 5360 11577 5427
rect 11675 5412 11704 5427
rect 11675 5360 11706 5412
rect 11560 5338 11706 5360
rect 11561 5046 11706 5338
rect 11561 4990 11583 5046
rect 11694 4990 11706 5046
rect 11561 4981 11706 4990
rect 1949 4928 2165 4938
rect 1949 4872 1975 4928
rect 2146 4872 2165 4928
rect 1949 4858 2165 4872
rect 2731 4934 2994 4943
rect 2731 4878 2775 4934
rect 2945 4878 2994 4934
rect 2731 4861 2994 4878
rect 7102 4923 7332 4939
rect 1020 4521 1037 4522
rect 1115 4521 1125 4522
rect 1020 4439 1035 4521
rect 1117 4439 1125 4521
rect 1020 4422 1125 4439
rect 1265 4514 1437 4528
rect 1265 4433 1281 4514
rect 1416 4433 1437 4514
rect 1530 4514 1702 4529
rect 1530 4475 1546 4514
rect 1529 4433 1546 4475
rect 1681 4433 1702 4514
rect 1265 4421 1440 4433
rect 1269 2106 1440 4421
rect 1529 4419 1702 4433
rect 1529 2216 1700 4419
rect 1966 2450 2152 4858
rect 2772 4213 2959 4861
rect 7102 4856 7125 4923
rect 7312 4856 7332 4923
rect 7102 4843 7332 4856
rect 15650 4860 16220 4880
rect 3467 4520 3641 4541
rect 3467 4440 3487 4520
rect 3465 4439 3487 4440
rect 3622 4440 3641 4520
rect 3823 4518 3997 4539
rect 3823 4513 3843 4518
rect 3622 4439 3643 4440
rect 2772 3143 2961 4213
rect 2774 2565 2961 3143
rect 3465 2912 3643 4439
rect 3822 4437 3843 4513
rect 3978 4437 3997 4518
rect 3822 4420 3997 4437
rect 4189 4513 4343 4533
rect 4189 4435 4216 4513
rect 4327 4435 4343 4513
rect 4189 4420 4343 4435
rect 4564 4516 4718 4536
rect 4564 4438 4591 4516
rect 4702 4438 4718 4516
rect 5079 4520 5254 4543
rect 5079 4462 5100 4520
rect 4564 4422 4718 4438
rect 5075 4439 5100 4462
rect 5235 4462 5254 4520
rect 5811 4518 5988 4541
rect 5235 4439 5257 4462
rect 5811 4453 5833 4518
rect 3822 3141 3995 4420
rect 5075 3242 5257 4439
rect 5808 4437 5833 4453
rect 5968 4437 5988 4518
rect 5808 4422 5988 4437
rect 5808 3582 5986 4422
rect 7120 4275 7287 4843
rect 15650 4740 15680 4860
rect 16170 4740 16220 4860
rect 15650 4710 16220 4740
rect 9269 4525 9442 4545
rect 9269 4444 9290 4525
rect 9425 4444 9442 4525
rect 11436 4528 11609 4548
rect 11436 4457 11457 4528
rect 9269 4440 9442 4444
rect 11435 4447 11457 4457
rect 11592 4447 11609 4528
rect 12896 4529 13069 4549
rect 12896 4512 12917 4529
rect 9269 4428 9445 4440
rect 7116 4209 7287 4275
rect 7116 3793 7283 4209
rect 9272 4002 9445 4428
rect 9271 3889 9445 4002
rect 11435 4215 11609 4447
rect 12895 4448 12917 4512
rect 13052 4448 13069 4529
rect 12895 4323 13069 4448
rect 13799 4529 13971 4547
rect 13799 4448 13829 4529
rect 13952 4448 13971 4529
rect 13799 4429 13971 4448
rect 12895 4225 12913 4323
rect 13054 4225 13069 4323
rect 11435 4100 11611 4215
rect 12895 4214 13069 4225
rect 11435 4017 11463 4100
rect 11591 4017 11611 4100
rect 11435 3997 11611 4017
rect 9271 3805 9301 3889
rect 9427 3805 9445 3889
rect 7115 3695 7289 3793
rect 9271 3787 9445 3805
rect 7115 3598 7142 3695
rect 7281 3598 7289 3695
rect 5808 3468 5990 3582
rect 7115 3581 7289 3598
rect 5808 3440 5847 3468
rect 5810 3379 5847 3440
rect 5975 3379 5990 3468
rect 5810 3362 5990 3379
rect 5075 3155 5102 3242
rect 5227 3155 5257 3242
rect 3818 3016 4003 3141
rect 5075 3134 5257 3155
rect 3818 2940 3850 3016
rect 3983 2940 4003 3016
rect 3818 2915 4003 2940
rect 3462 2795 3646 2912
rect 3462 2707 3483 2795
rect 3635 2707 3646 2795
rect 3462 2685 3646 2707
rect 2774 2471 2794 2565
rect 2941 2478 2961 2565
rect 2941 2471 2956 2478
rect 2774 2453 2956 2471
rect 1961 2329 2148 2450
rect 1961 2234 1979 2329
rect 2134 2234 2148 2329
rect 1961 2220 2148 2234
rect 1270 1984 1439 2106
rect 1526 2102 1701 2216
rect 1526 2004 1549 2102
rect 1673 2004 1701 2102
rect 1526 1989 1701 2004
rect 1269 1874 1441 1984
rect 1269 1767 1290 1874
rect 1421 1767 1441 1874
rect 1269 1751 1441 1767
rect 1812 883 1950 895
rect 523 822 1163 823
rect 523 731 1449 822
rect 1812 807 1841 883
rect 1912 807 1950 883
rect 1812 783 1950 807
rect 809 730 1449 731
rect 1362 650 1449 730
rect 15650 739 16208 750
rect 15650 682 15685 739
rect 16183 682 16208 739
rect 15650 667 16208 682
rect 4268 650 7355 651
rect 10144 650 11805 651
rect 1362 649 7355 650
rect 8073 649 11805 650
rect 1362 603 11805 649
rect 1364 572 11805 603
rect 1364 570 4276 572
rect 1044 552 1125 553
rect 262 540 1125 552
rect 262 457 1054 540
rect 1123 509 1125 540
rect 1364 530 1449 570
rect 1123 457 1126 509
rect 262 439 1126 457
rect 1364 462 1374 530
rect 1442 462 1449 530
rect 1364 448 1449 462
rect 1041 135 1126 439
rect 3754 435 3835 450
rect 3754 377 3768 435
rect 3826 377 3835 435
rect 4079 431 4158 570
rect 5180 433 5254 572
rect 5484 437 5572 452
rect 3754 364 3835 377
rect 4073 415 4163 431
rect 4073 353 4088 415
rect 4150 353 4163 415
rect 4395 410 4482 413
rect 4073 339 4163 353
rect 4393 401 4482 410
rect 4393 340 4405 401
rect 4472 340 4482 401
rect 4393 136 4482 340
rect 4849 410 4934 421
rect 4849 353 4862 410
rect 4924 353 4934 410
rect 4849 339 4934 353
rect 5165 420 5257 433
rect 5165 359 5180 420
rect 5245 359 5257 420
rect 5484 377 5505 437
rect 5562 377 5572 437
rect 5484 366 5572 377
rect 7551 436 7630 448
rect 7551 377 7564 436
rect 7620 435 7630 436
rect 7551 376 7565 377
rect 7621 376 7630 435
rect 7864 428 7943 572
rect 8073 571 11805 572
rect 7551 365 7630 376
rect 7862 420 7950 428
rect 8962 424 9033 571
rect 9273 436 9359 446
rect 5165 348 5257 359
rect 7862 364 7877 420
rect 7935 364 7950 420
rect 7862 350 7950 364
rect 8182 415 8276 422
rect 8182 353 8200 415
rect 8264 353 8276 415
rect 8955 412 9040 424
rect 8182 346 8276 353
rect 8636 400 8719 410
rect 4851 136 4931 339
rect 4393 135 5964 136
rect 1041 134 5964 135
rect 8188 134 8271 346
rect 8636 339 8646 400
rect 8711 339 8719 400
rect 8955 354 8970 412
rect 9030 354 9040 412
rect 9273 377 9292 436
rect 9349 378 9359 436
rect 11669 425 11746 571
rect 9348 377 9359 378
rect 9273 364 9359 377
rect 11663 415 11752 425
rect 8955 345 9040 354
rect 11663 359 11678 415
rect 11740 359 11752 415
rect 11663 347 11752 359
rect 11982 408 12073 419
rect 8636 326 8719 339
rect 11982 344 11994 408
rect 12061 344 12073 408
rect 11982 334 12073 344
rect 1041 132 8300 134
rect 8646 132 8711 326
rect 1041 131 8747 132
rect 11986 131 12070 334
rect 1041 58 12086 131
rect 4497 57 12086 58
rect 5956 55 12086 57
rect 8722 54 12086 55
rect 16407 100 16967 113
rect 16407 43 16481 100
rect 16942 43 16967 100
rect 16407 26 16967 43
rect 299 -56 1233 -55
rect 299 -57 1636 -56
rect 299 -67 14486 -57
rect 299 -138 312 -67
rect 381 -138 14486 -67
rect 299 -149 14486 -138
rect 1766 -273 14475 -258
rect 1766 -354 1775 -273
rect 1832 -354 14475 -273
rect 1766 -364 14475 -354
rect 3661 -457 14477 -456
rect 3659 -468 14477 -457
rect 3659 -540 3672 -468
rect 3729 -536 14477 -468
rect 3729 -540 14475 -536
rect 3659 -552 14475 -540
rect 5559 -670 14473 -640
rect 5559 -671 5570 -670
rect 5559 -678 5567 -671
rect 5558 -730 5567 -678
rect 5558 -731 5570 -730
rect 5626 -731 14473 -670
rect 5558 -737 14473 -731
rect 5559 -738 5759 -737
rect 7464 -830 7691 -829
rect 7464 -855 14464 -830
rect 7464 -919 7478 -855
rect 7543 -919 14464 -855
rect 7464 -929 14464 -919
rect 9301 -1025 10693 -1024
rect 9301 -1035 14461 -1025
rect 9301 -1107 9320 -1035
rect 9391 -1107 14461 -1035
rect 9301 -1123 14461 -1107
rect 11181 -1218 11340 -1217
rect 11181 -1219 12613 -1218
rect 11181 -1238 14459 -1219
rect 11181 -1307 11193 -1238
rect 11257 -1307 14459 -1238
rect 11181 -1317 14459 -1307
<< via3 >>
rect 15719 10475 16169 10570
rect 1192 10292 1423 10293
rect 1192 10204 1423 10292
rect 1192 10201 1423 10204
rect 16480 8246 16937 8349
rect 16496 6678 16910 6773
rect 1045 6048 1046 6117
rect 1046 6048 1109 6117
rect 1109 6048 1111 6117
rect -480 799 -353 873
rect 1037 4521 1115 4522
rect 1037 4440 1115 4521
rect 4216 4435 4327 4513
rect 4591 4438 4702 4516
rect 15680 4740 16170 4860
rect 13829 4448 13952 4529
rect 12913 4225 13054 4323
rect 11463 4017 11591 4100
rect 9301 3805 9427 3889
rect 7142 3598 7281 3695
rect 5847 3379 5975 3468
rect 5102 3155 5227 3242
rect 3850 2940 3983 3016
rect 3483 2707 3635 2795
rect 2794 2471 2941 2565
rect 1979 2234 2134 2329
rect 1549 2004 1673 2102
rect 1290 1767 1421 1874
rect 1841 807 1912 883
rect 15685 682 16183 739
rect 3770 377 3825 435
rect 3825 377 3826 435
rect 5505 436 5562 437
rect 5505 377 5562 436
rect 7565 377 7620 435
rect 7620 377 7621 435
rect 7565 376 7621 377
rect 9292 435 9349 436
rect 9292 378 9348 435
rect 9348 378 9349 435
rect 16481 43 16942 100
<< metal4 >>
rect 15650 10570 16220 11140
rect 15650 10475 15719 10570
rect 16169 10475 16220 10570
rect 1020 10293 1450 10320
rect 1020 10201 1192 10293
rect 1423 10201 1450 10293
rect 1020 10179 1450 10201
rect 1024 7360 1120 10179
rect 1024 6150 1121 7360
rect 1024 6135 1123 6150
rect 1020 6117 1125 6135
rect 1020 6048 1045 6117
rect 1111 6048 1125 6117
rect 1020 4535 1125 6048
rect 15650 4880 16220 10475
rect 15649 4860 16220 4880
rect 15649 4740 15680 4860
rect 16170 4740 16220 4860
rect 15649 4706 16220 4740
rect 13236 4547 13969 4548
rect 13236 4545 13971 4547
rect 12149 4544 13971 4545
rect 8832 4541 10219 4542
rect 11436 4541 11610 4544
rect 11889 4541 13971 4544
rect 8832 4540 13971 4541
rect 989 4533 1682 4535
rect 2314 4533 3152 4535
rect 3467 4534 3641 4539
rect 3465 4533 3642 4534
rect 989 4532 3735 4533
rect 3823 4532 3997 4537
rect 5079 4536 5254 4539
rect 6564 4537 13971 4540
rect 5406 4536 13971 4537
rect 4527 4534 13971 4536
rect 4300 4533 13971 4534
rect 4188 4532 13971 4533
rect 989 4529 13971 4532
rect 989 4522 13829 4529
rect 989 4440 1037 4522
rect 1115 4516 13829 4522
rect 1115 4513 4591 4516
rect 1115 4440 4216 4513
rect 989 4435 4216 4440
rect 4327 4438 4591 4513
rect 4702 4448 13829 4516
rect 13952 4448 13971 4529
rect 4702 4438 13971 4448
rect 4327 4435 13971 4438
rect 989 4431 13971 4435
rect 989 4430 13049 4431
rect 989 4428 9552 4430
rect 9935 4429 12233 4430
rect 13799 4429 13971 4431
rect 989 4425 6793 4428
rect 7469 4427 9552 4428
rect 989 4424 5988 4425
rect 989 4422 5687 4424
rect 5811 4422 5988 4424
rect 989 4420 4344 4422
rect 1515 4418 2353 4420
rect 3102 4419 4333 4420
rect 945 4343 5410 4345
rect 945 4342 12399 4343
rect 945 4341 13065 4342
rect 464 4340 13065 4341
rect 464 4323 13069 4340
rect 464 4225 12913 4323
rect 13054 4225 13069 4323
rect 464 4224 13069 4225
rect 945 4221 13069 4224
rect 5144 4217 13069 4221
rect 10963 4215 13069 4217
rect 12357 4214 13069 4215
rect 5144 4124 11461 4126
rect 3465 4121 11610 4124
rect 461 4100 11610 4121
rect 461 4017 11463 4100
rect 11591 4017 11610 4100
rect 461 4000 11610 4017
rect 991 3997 3685 4000
rect 11414 3998 11610 4000
rect 985 3919 3679 3921
rect 985 3918 5449 3919
rect 985 3917 8473 3918
rect 985 3915 9449 3917
rect 464 3889 9449 3915
rect 464 3805 9301 3889
rect 9427 3805 9449 3889
rect 464 3797 9449 3805
rect 464 3794 1001 3797
rect 3528 3795 9449 3797
rect 5150 3794 9449 3795
rect 8372 3787 9449 3794
rect 6887 3705 7288 3708
rect 985 3699 1211 3701
rect 456 3698 3765 3699
rect 5141 3698 7288 3705
rect 456 3695 7288 3698
rect 456 3598 7142 3695
rect 7281 3598 7288 3695
rect 456 3581 7288 3598
rect 456 3578 5449 3581
rect 985 3575 5449 3578
rect 3528 3574 5449 3575
rect 4082 3491 5717 3492
rect 4082 3490 5988 3491
rect 440 3487 993 3489
rect 440 3485 1207 3487
rect 3542 3485 5988 3490
rect 440 3468 5988 3485
rect 440 3379 5847 3468
rect 5975 3379 5988 3468
rect 440 3364 5988 3379
rect 981 3362 5988 3364
rect 981 3361 5717 3362
rect 3542 3359 5717 3361
rect 3542 3357 5177 3359
rect 4886 3266 5255 3270
rect 982 3262 1208 3264
rect 2230 3262 5255 3266
rect 982 3261 5255 3262
rect 437 3242 5255 3261
rect 437 3155 5102 3242
rect 5227 3155 5255 3242
rect 437 3142 5255 3155
rect 437 3138 3842 3142
rect 437 3136 990 3138
rect 4886 3135 5255 3142
rect 1675 3041 3109 3042
rect 1675 3040 4004 3041
rect 981 3036 4004 3040
rect 441 3016 4004 3036
rect 441 2940 3850 3016
rect 3983 2940 4004 3016
rect 441 2915 4004 2940
rect 441 2911 3109 2915
rect 981 2909 2415 2911
rect 1711 2809 3651 2814
rect 969 2799 3651 2809
rect 427 2795 3651 2799
rect 427 2707 3483 2795
rect 3635 2707 3651 2795
rect 427 2686 3651 2707
rect 427 2683 3145 2686
rect 427 2678 2403 2683
rect 427 2674 980 2678
rect 1814 2585 2967 2587
rect 956 2582 2967 2585
rect 412 2565 2967 2582
rect 412 2471 2794 2565
rect 2941 2471 2967 2565
rect 412 2457 2967 2471
rect 956 2452 2967 2457
rect 956 2447 2319 2452
rect 960 2356 1777 2358
rect 401 2354 1777 2356
rect 401 2329 2154 2354
rect 401 2234 1979 2329
rect 2134 2234 2154 2329
rect 401 2223 2154 2234
rect 401 2221 967 2223
rect 1339 2218 2154 2223
rect 918 2122 1702 2127
rect 366 2102 1702 2122
rect 366 2004 1549 2102
rect 1673 2004 1702 2102
rect 366 1987 1702 2004
rect 918 1983 1702 1987
rect 362 1889 928 1890
rect 362 1874 1444 1889
rect 362 1767 1290 1874
rect 1421 1767 1444 1874
rect 362 1755 1444 1767
rect 857 1745 1444 1755
rect -491 887 1150 888
rect 1812 887 1950 895
rect -491 883 1950 887
rect -491 873 1841 883
rect -491 799 -480 873
rect -353 807 1841 873
rect 1912 807 1950 883
rect -353 799 1950 807
rect -491 791 1950 799
rect -491 780 -339 791
rect 296 790 1950 791
rect 1812 783 1950 790
rect 15650 739 16220 4706
rect 15650 682 15685 739
rect 16183 682 16220 739
rect 3754 437 5570 452
rect 3754 435 5505 437
rect 3754 377 3770 435
rect 3826 377 5505 435
rect 5562 377 5570 437
rect 3754 364 5570 377
rect 7549 436 9360 452
rect 7549 435 9292 436
rect 7549 376 7565 435
rect 7621 378 9292 435
rect 9349 378 9360 436
rect 7621 376 9360 378
rect 7549 362 9360 376
rect 15650 -1310 16220 682
rect 16400 8349 16970 11150
rect 16400 8246 16480 8349
rect 16937 8246 16970 8349
rect 16400 6773 16970 8246
rect 16400 6678 16496 6773
rect 16910 6678 16970 6773
rect 16400 100 16970 6678
rect 16400 43 16481 100
rect 16942 43 16970 100
rect 16400 -1300 16970 43
use switch_C5  switch_C5_0
timestamp 1757325932
transform 1 0 558 0 1 346
box 308 -346 2174 443
use switch_C5  switch_C5_1
timestamp 1757325932
transform -1 0 4965 0 1 346
box 308 -346 2174 443
use switch_C5  switch_C5_2
timestamp 1757325932
transform 1 0 4362 0 1 346
box 308 -346 2174 443
use switch_C5  switch_C5_3
timestamp 1757325932
transform -1 0 8754 0 1 346
box 308 -346 2174 443
use switch_C5  switch_C5_4
timestamp 1757325932
transform 1 0 8150 0 1 346
box 308 -346 2174 443
use switch_C5  switch_C5_5
timestamp 1757325932
transform -1 0 12554 0 1 346
box 308 -346 2174 443
use switch_C9  switch_C9_0
timestamp 1757325240
transform -1 0 16617 0 -1 19638
box 2498 12794 8634 14978
use switch_VCM  switch_VCM_0
timestamp 1757325446
transform 1 0 12188 0 1 7930
box 398 249 3158 2595
use switches_6  switches_6_0
timestamp 1757241197
transform -1 0 5024 0 -1 6808
box 2684 -115 4128 2198
use switches_7  switches_7_0
timestamp 1757239750
transform 1 0 -327 0 -1 9286
box 2088 -262 4831 4676
use switches_8  switches_8_0
timestamp 1757235861
transform -1 0 7972 0 -1 12273
box 27 5379 3480 7722
use switches_10  switches_10_0
timestamp 1757233555
transform -1 0 15289 0 1 8656
box 2730 -483 14380 2010
use switches_dummy  switches_dummy_0
timestamp 1757242206
transform 1 0 232 0 1 342
box -232 -342 634 827
<< labels >>
flabel metal3 14152 -145 14481 -62 0 FreeSans 320 0 0 0 Cbtm_0_dummy
port 6 nsew
flabel metal3 14139 -358 14470 -264 0 FreeSans 320 0 0 0 Cbtm_0
port 7 nsew
flabel metal3 14144 -543 14471 -463 0 FreeSans 320 0 0 0 Cbtm_1
port 8 nsew
flabel metal3 14142 -727 14469 -647 0 FreeSans 320 0 0 0 Cbtm_2
port 9 nsew
flabel metal3 14163 -923 14457 -838 0 FreeSans 320 0 0 0 Cbtm_3
port 10 nsew
flabel metal3 14180 -1118 14454 -1033 0 FreeSans 320 0 0 0 Cbtm_4
port 11 nsew
flabel metal3 14199 -1312 14454 -1227 0 FreeSans 320 0 0 0 Cbtm_5
port 12 nsew
flabel metal3 13761 7040 14086 7142 0 FreeSans 320 0 0 0 Cbtm_6
port 13 nsew
flabel metal3 13768 7291 14093 7393 0 FreeSans 320 0 0 0 Cbtm_7
port 14 nsew
flabel metal3 13750 7534 14075 7636 0 FreeSans 320 0 0 0 Cbtm_8
port 15 nsew
flabel metal3 13743 7795 14068 7897 0 FreeSans 320 0 0 0 Cbtm_9
port 16 nsew
flabel metal3 13740 7997 14065 8099 0 FreeSans 320 0 0 0 Cbtm_10
port 17 nsew
flabel metal2 377 10384 512 10571 0 FreeSans 320 0 0 0 VIN
port 4 nsew
flabel metal2 -483 10383 -348 10570 0 FreeSans 320 0 0 0 VREF
port 3 nsew
flabel metal2 -214 10348 -56 10566 0 FreeSans 320 0 0 0 VCM
port 1 nsew
flabel metal2 94 10370 245 10550 0 FreeSans 320 0 0 0 VREF_GND
port 2 nsew
flabel metal3 13847 6848 14094 6954 0 FreeSans 160 0 0 0 VDAC
port 18 nsew
flabel metal2 13830 1357 14144 1452 0 FreeSans 160 0 0 0 EN_VIN
port 19 nsew
flabel metal2 9830 10700 10021 10809 0 FreeSans 160 0 0 0 EN_VREF_Z[10]
port 20 nsew
flabel metal4 472 3800 750 3906 0 FreeSans 160 0 0 0 EN_VREF_Z[9]
port 21 nsew
flabel metal4 463 3586 769 3694 0 FreeSans 160 0 0 0 EN_VREF_Z[8]
port 22 nsew
flabel metal4 420 2464 763 2576 0 FreeSans 160 0 0 0 EN_VREF_Z[7]
port 23 nsew
flabel metal4 405 2225 753 2354 0 FreeSans 160 0 0 0 EN_VREF_Z[6]
port 24 nsew
flabel metal2 13868 3877 14160 3986 0 FreeSans 160 0 0 0 EN_VREF_Z[5]
port 25 nsew
flabel metal2 13925 3695 14173 3806 0 FreeSans 160 0 0 0 EN_VREF_Z[4]
port 26 nsew
flabel metal2 13869 2819 14141 2923 0 FreeSans 160 0 0 0 EN_VREF_Z[3]
port 27 nsew
flabel metal2 13899 2633 14143 2744 0 FreeSans 160 0 0 0 EN_VREF_Z[2]
port 28 nsew
flabel metal2 13822 1709 14141 1807 0 FreeSans 160 0 0 0 EN_VREF_Z[1]
port 29 nsew
flabel metal2 13838 1535 14140 1633 0 FreeSans 160 0 0 0 EN_VREF_Z[0]
port 30 nsew
flabel metal2 2803 10653 3036 10757 0 FreeSans 160 0 0 0 EN_VSS[10]
port 31 nsew
flabel metal4 469 4005 725 4114 0 FreeSans 160 0 0 0 EN_VSS[9]
port 32 nsew
flabel metal4 446 3142 733 3257 0 FreeSans 160 0 0 0 EN_VSS[8]
port 33 nsew
flabel metal4 450 2918 740 3032 0 FreeSans 160 0 0 0 EN_VSS[7]
port 34 nsew
flabel metal4 378 1764 735 1881 0 FreeSans 160 0 0 0 EN_VSS[6]
port 35 nsew
flabel metal2 13846 4064 14171 4173 0 FreeSans 160 0 0 0 EN_VSS[5]
port 36 nsew
flabel metal2 13915 3526 14149 3625 0 FreeSans 160 0 0 0 EN_VSS[4]
port 37 nsew
flabel metal2 13876 2998 14148 3103 0 FreeSans 160 0 0 0 EN_VSS[3]
port 38 nsew
flabel metal2 13899 2462 14139 2563 0 FreeSans 160 0 0 0 EN_VSS[2]
port 39 nsew
flabel metal2 13885 1922 14136 2024 0 FreeSans 160 0 0 0 EN_VSS[1]
port 40 nsew
flabel metal2 13865 1178 14136 1281 0 FreeSans 160 0 0 0 EN_VSS[0]
port 41 nsew
flabel metal2 5646 10612 5873 10736 0 FreeSans 160 0 0 0 EN_VCM[10]
port 42 nsew
flabel metal4 473 4233 767 4333 0 FreeSans 160 0 0 0 EN_VCM[9]
port 43 nsew
flabel metal4 449 3373 760 3485 0 FreeSans 160 0 0 0 EN_VCM[8]
port 44 nsew
flabel metal4 434 2677 715 2793 0 FreeSans 160 0 0 0 EN_VCM[7]
port 45 nsew
flabel metal4 382 1993 737 2117 0 FreeSans 160 0 0 0 EN_VCM[6]
port 46 nsew
flabel metal2 13845 4252 14167 4349 0 FreeSans 160 0 0 0 EN_VCM[5]
port 47 nsew
flabel metal2 13820 3351 14142 3448 0 FreeSans 160 0 0 0 EN_VCM[4]
port 48 nsew
flabel metal2 13820 3174 14142 3271 0 FreeSans 160 0 0 0 EN_VCM[3]
port 49 nsew
flabel metal2 13865 2290 14141 2385 0 FreeSans 160 0 0 0 EN_VCM[2]
port 50 nsew
flabel metal2 13861 2106 14137 2201 0 FreeSans 160 0 0 0 EN_VCM[1]
port 51 nsew
flabel metal2 13888 1013 14141 1094 0 FreeSans 160 0 0 0 EN_VCM[0]
port 52 nsew
flabel metal1 -621 1213 -278 1360 0 FreeSans 160 0 0 0 EN_VCM_DUMMY
port 53 nsew
flabel metal2 13905 10650 14142 10795 0 FreeSans 160 0 0 0 EN_VCM_SW
port 54 nsew
flabel metal4 15700 -1220 16170 11040 0 FreeSans 480 0 0 0 VDD
port 5 nsew
flabel metal4 16450 -1210 16920 11050 0 FreeSans 480 0 0 0 VSS
port 55 nsew
<< end >>
