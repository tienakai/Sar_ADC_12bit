magic
tech gf180mcuD
magscale 1 10
timestamp 1757233555
<< nwell >>
rect 2730 -311 8149 2002
rect 2730 -483 8150 -311
<< pwell >>
rect 8149 2001 14380 2010
rect 8149 1546 14379 2001
rect 8149 -190 14380 1546
rect 8149 -311 14379 -190
rect 8150 -451 14379 -311
rect 8150 -480 14380 -451
rect 8150 -481 14379 -480
<< nmos >>
rect 8352 -122 8408 1478
rect 8512 -122 8568 1478
rect 8672 -122 8728 1478
rect 8832 -122 8888 1478
rect 8992 -122 9048 1478
rect 9152 -122 9208 1478
rect 9312 -122 9368 1478
rect 9472 -122 9528 1478
rect 9632 -122 9688 1478
rect 9792 -122 9848 1478
rect 9952 -122 10008 1478
rect 10112 -122 10168 1478
rect 10272 -122 10328 1478
rect 10432 -122 10488 1478
rect 10592 -122 10648 1478
rect 10752 -122 10808 1478
rect 11041 -122 11097 1478
rect 11201 -122 11257 1478
rect 11361 -122 11417 1478
rect 11521 -122 11577 1478
rect 11681 -122 11737 1478
rect 11841 -122 11897 1478
rect 12001 -122 12057 1478
rect 12161 -122 12217 1478
rect 12321 -122 12377 1478
rect 12481 -122 12537 1478
rect 12641 -122 12697 1478
rect 12801 -122 12857 1478
rect 12961 -122 13017 1478
rect 13121 -122 13177 1478
rect 13281 -122 13337 1478
rect 13441 -122 13497 1478
rect 13732 -122 13788 1478
rect 13892 -122 13948 1478
rect 14052 -122 14108 1478
rect 14212 -122 14268 1478
<< pmos >>
rect 2914 -120 2970 1480
rect 3074 -120 3130 1480
rect 3234 -120 3290 1480
rect 3394 -120 3450 1480
rect 3554 -120 3610 1480
rect 3714 -120 3770 1480
rect 3874 -120 3930 1480
rect 4034 -120 4090 1480
rect 4194 -120 4250 1480
rect 4354 -120 4410 1480
rect 4514 -120 4570 1480
rect 4674 -120 4730 1480
rect 4834 -120 4890 1480
rect 4994 -120 5050 1480
rect 5154 -120 5210 1480
rect 5314 -120 5370 1480
rect 5474 -120 5530 1480
rect 5634 -120 5690 1480
rect 5794 -120 5850 1480
rect 5954 -120 6010 1480
rect 6114 -120 6170 1480
rect 6274 -120 6330 1480
rect 6434 -120 6490 1480
rect 6594 -120 6650 1480
rect 6754 -120 6810 1480
rect 6914 -120 6970 1480
rect 7074 -120 7130 1480
rect 7234 -120 7290 1480
rect 7394 -120 7450 1480
rect 7554 -120 7610 1480
rect 7714 -120 7770 1480
rect 7874 -120 7930 1480
<< ndiff >>
rect 8264 1465 8352 1478
rect 8264 -109 8277 1465
rect 8323 -109 8352 1465
rect 8264 -122 8352 -109
rect 8408 1465 8512 1478
rect 8408 -109 8437 1465
rect 8483 -109 8512 1465
rect 8408 -122 8512 -109
rect 8568 1465 8672 1478
rect 8568 -109 8597 1465
rect 8643 -109 8672 1465
rect 8568 -122 8672 -109
rect 8728 1465 8832 1478
rect 8728 -109 8757 1465
rect 8803 -109 8832 1465
rect 8728 -122 8832 -109
rect 8888 1465 8992 1478
rect 8888 -109 8917 1465
rect 8963 -109 8992 1465
rect 8888 -122 8992 -109
rect 9048 1465 9152 1478
rect 9048 -109 9077 1465
rect 9123 -109 9152 1465
rect 9048 -122 9152 -109
rect 9208 1465 9312 1478
rect 9208 -109 9237 1465
rect 9283 -109 9312 1465
rect 9208 -122 9312 -109
rect 9368 1465 9472 1478
rect 9368 -109 9397 1465
rect 9443 -109 9472 1465
rect 9368 -122 9472 -109
rect 9528 1465 9632 1478
rect 9528 -109 9557 1465
rect 9603 -109 9632 1465
rect 9528 -122 9632 -109
rect 9688 1465 9792 1478
rect 9688 -109 9717 1465
rect 9763 -109 9792 1465
rect 9688 -122 9792 -109
rect 9848 1465 9952 1478
rect 9848 -109 9877 1465
rect 9923 -109 9952 1465
rect 9848 -122 9952 -109
rect 10008 1465 10112 1478
rect 10008 -109 10037 1465
rect 10083 -109 10112 1465
rect 10008 -122 10112 -109
rect 10168 1465 10272 1478
rect 10168 -109 10197 1465
rect 10243 -109 10272 1465
rect 10168 -122 10272 -109
rect 10328 1465 10432 1478
rect 10328 -109 10357 1465
rect 10403 -109 10432 1465
rect 10328 -122 10432 -109
rect 10488 1465 10592 1478
rect 10488 -109 10517 1465
rect 10563 -109 10592 1465
rect 10488 -122 10592 -109
rect 10648 1465 10752 1478
rect 10648 -109 10677 1465
rect 10723 -109 10752 1465
rect 10648 -122 10752 -109
rect 10808 1465 10896 1478
rect 10808 -109 10837 1465
rect 10883 -109 10896 1465
rect 10808 -122 10896 -109
rect 10953 1465 11041 1478
rect 10953 -109 10966 1465
rect 11012 -109 11041 1465
rect 10953 -122 11041 -109
rect 11097 1465 11201 1478
rect 11097 -109 11126 1465
rect 11172 -109 11201 1465
rect 11097 -122 11201 -109
rect 11257 1465 11361 1478
rect 11257 -109 11286 1465
rect 11332 -109 11361 1465
rect 11257 -122 11361 -109
rect 11417 1465 11521 1478
rect 11417 -109 11446 1465
rect 11492 -109 11521 1465
rect 11417 -122 11521 -109
rect 11577 1465 11681 1478
rect 11577 -109 11606 1465
rect 11652 -109 11681 1465
rect 11577 -122 11681 -109
rect 11737 1465 11841 1478
rect 11737 -109 11766 1465
rect 11812 -109 11841 1465
rect 11737 -122 11841 -109
rect 11897 1465 12001 1478
rect 11897 -109 11926 1465
rect 11972 -109 12001 1465
rect 11897 -122 12001 -109
rect 12057 1465 12161 1478
rect 12057 -109 12086 1465
rect 12132 -109 12161 1465
rect 12057 -122 12161 -109
rect 12217 1465 12321 1478
rect 12217 -109 12246 1465
rect 12292 -109 12321 1465
rect 12217 -122 12321 -109
rect 12377 1465 12481 1478
rect 12377 -109 12406 1465
rect 12452 -109 12481 1465
rect 12377 -122 12481 -109
rect 12537 1465 12641 1478
rect 12537 -109 12566 1465
rect 12612 -109 12641 1465
rect 12537 -122 12641 -109
rect 12697 1465 12801 1478
rect 12697 -109 12726 1465
rect 12772 -109 12801 1465
rect 12697 -122 12801 -109
rect 12857 1465 12961 1478
rect 12857 -109 12886 1465
rect 12932 -109 12961 1465
rect 12857 -122 12961 -109
rect 13017 1465 13121 1478
rect 13017 -109 13046 1465
rect 13092 -109 13121 1465
rect 13017 -122 13121 -109
rect 13177 1465 13281 1478
rect 13177 -109 13206 1465
rect 13252 -109 13281 1465
rect 13177 -122 13281 -109
rect 13337 1465 13441 1478
rect 13337 -109 13366 1465
rect 13412 -109 13441 1465
rect 13337 -122 13441 -109
rect 13497 1465 13585 1478
rect 13497 -109 13526 1465
rect 13572 -109 13585 1465
rect 13497 -122 13585 -109
rect 13644 1465 13732 1478
rect 13644 -109 13657 1465
rect 13703 -109 13732 1465
rect 13644 -122 13732 -109
rect 13788 1465 13892 1478
rect 13788 -109 13817 1465
rect 13863 -109 13892 1465
rect 13788 -122 13892 -109
rect 13948 1465 14052 1478
rect 13948 -109 13977 1465
rect 14023 -109 14052 1465
rect 13948 -122 14052 -109
rect 14108 1465 14212 1478
rect 14108 -109 14137 1465
rect 14183 -109 14212 1465
rect 14108 -122 14212 -109
rect 14268 1465 14356 1478
rect 14268 -109 14297 1465
rect 14343 -109 14356 1465
rect 14268 -122 14356 -109
<< pdiff >>
rect 2826 1467 2914 1480
rect 2826 -107 2839 1467
rect 2885 -107 2914 1467
rect 2826 -120 2914 -107
rect 2970 1467 3074 1480
rect 2970 -107 2999 1467
rect 3045 -107 3074 1467
rect 2970 -120 3074 -107
rect 3130 1467 3234 1480
rect 3130 -107 3159 1467
rect 3205 -107 3234 1467
rect 3130 -120 3234 -107
rect 3290 1467 3394 1480
rect 3290 -107 3319 1467
rect 3365 -107 3394 1467
rect 3290 -120 3394 -107
rect 3450 1467 3554 1480
rect 3450 -107 3479 1467
rect 3525 -107 3554 1467
rect 3450 -120 3554 -107
rect 3610 1467 3714 1480
rect 3610 -107 3639 1467
rect 3685 -107 3714 1467
rect 3610 -120 3714 -107
rect 3770 1467 3874 1480
rect 3770 -107 3799 1467
rect 3845 -107 3874 1467
rect 3770 -120 3874 -107
rect 3930 1467 4034 1480
rect 3930 -107 3959 1467
rect 4005 -107 4034 1467
rect 3930 -120 4034 -107
rect 4090 1467 4194 1480
rect 4090 -107 4119 1467
rect 4165 -107 4194 1467
rect 4090 -120 4194 -107
rect 4250 1467 4354 1480
rect 4250 -107 4279 1467
rect 4325 -107 4354 1467
rect 4250 -120 4354 -107
rect 4410 1467 4514 1480
rect 4410 -107 4439 1467
rect 4485 -107 4514 1467
rect 4410 -120 4514 -107
rect 4570 1467 4674 1480
rect 4570 -107 4599 1467
rect 4645 -107 4674 1467
rect 4570 -120 4674 -107
rect 4730 1467 4834 1480
rect 4730 -107 4759 1467
rect 4805 -107 4834 1467
rect 4730 -120 4834 -107
rect 4890 1467 4994 1480
rect 4890 -107 4919 1467
rect 4965 -107 4994 1467
rect 4890 -120 4994 -107
rect 5050 1467 5154 1480
rect 5050 -107 5079 1467
rect 5125 -107 5154 1467
rect 5050 -120 5154 -107
rect 5210 1467 5314 1480
rect 5210 -107 5239 1467
rect 5285 -107 5314 1467
rect 5210 -120 5314 -107
rect 5370 1467 5474 1480
rect 5370 -107 5399 1467
rect 5445 -107 5474 1467
rect 5370 -120 5474 -107
rect 5530 1467 5634 1480
rect 5530 -107 5559 1467
rect 5605 -107 5634 1467
rect 5530 -120 5634 -107
rect 5690 1467 5794 1480
rect 5690 -107 5719 1467
rect 5765 -107 5794 1467
rect 5690 -120 5794 -107
rect 5850 1467 5954 1480
rect 5850 -107 5879 1467
rect 5925 -107 5954 1467
rect 5850 -120 5954 -107
rect 6010 1467 6114 1480
rect 6010 -107 6039 1467
rect 6085 -107 6114 1467
rect 6010 -120 6114 -107
rect 6170 1467 6274 1480
rect 6170 -107 6199 1467
rect 6245 -107 6274 1467
rect 6170 -120 6274 -107
rect 6330 1467 6434 1480
rect 6330 -107 6359 1467
rect 6405 -107 6434 1467
rect 6330 -120 6434 -107
rect 6490 1467 6594 1480
rect 6490 -107 6519 1467
rect 6565 -107 6594 1467
rect 6490 -120 6594 -107
rect 6650 1467 6754 1480
rect 6650 -107 6679 1467
rect 6725 -107 6754 1467
rect 6650 -120 6754 -107
rect 6810 1467 6914 1480
rect 6810 -107 6839 1467
rect 6885 -107 6914 1467
rect 6810 -120 6914 -107
rect 6970 1467 7074 1480
rect 6970 -107 6999 1467
rect 7045 -107 7074 1467
rect 6970 -120 7074 -107
rect 7130 1467 7234 1480
rect 7130 -107 7159 1467
rect 7205 -107 7234 1467
rect 7130 -120 7234 -107
rect 7290 1467 7394 1480
rect 7290 -107 7319 1467
rect 7365 -107 7394 1467
rect 7290 -120 7394 -107
rect 7450 1467 7554 1480
rect 7450 -107 7479 1467
rect 7525 -107 7554 1467
rect 7450 -120 7554 -107
rect 7610 1467 7714 1480
rect 7610 -107 7639 1467
rect 7685 -107 7714 1467
rect 7610 -120 7714 -107
rect 7770 1467 7874 1480
rect 7770 -107 7799 1467
rect 7845 -107 7874 1467
rect 7770 -120 7874 -107
rect 7930 1467 8018 1480
rect 7930 -107 7959 1467
rect 8005 -107 8018 1467
rect 7930 -120 8018 -107
<< ndiffc >>
rect 8277 -109 8323 1465
rect 8437 -109 8483 1465
rect 8597 -109 8643 1465
rect 8757 -109 8803 1465
rect 8917 -109 8963 1465
rect 9077 -109 9123 1465
rect 9237 -109 9283 1465
rect 9397 -109 9443 1465
rect 9557 -109 9603 1465
rect 9717 -109 9763 1465
rect 9877 -109 9923 1465
rect 10037 -109 10083 1465
rect 10197 -109 10243 1465
rect 10357 -109 10403 1465
rect 10517 -109 10563 1465
rect 10677 -109 10723 1465
rect 10837 -109 10883 1465
rect 10966 -109 11012 1465
rect 11126 -109 11172 1465
rect 11286 -109 11332 1465
rect 11446 -109 11492 1465
rect 11606 -109 11652 1465
rect 11766 -109 11812 1465
rect 11926 -109 11972 1465
rect 12086 -109 12132 1465
rect 12246 -109 12292 1465
rect 12406 -109 12452 1465
rect 12566 -109 12612 1465
rect 12726 -109 12772 1465
rect 12886 -109 12932 1465
rect 13046 -109 13092 1465
rect 13206 -109 13252 1465
rect 13366 -109 13412 1465
rect 13526 -109 13572 1465
rect 13657 -109 13703 1465
rect 13817 -109 13863 1465
rect 13977 -109 14023 1465
rect 14137 -109 14183 1465
rect 14297 -109 14343 1465
<< pdiffc >>
rect 2839 -107 2885 1467
rect 2999 -107 3045 1467
rect 3159 -107 3205 1467
rect 3319 -107 3365 1467
rect 3479 -107 3525 1467
rect 3639 -107 3685 1467
rect 3799 -107 3845 1467
rect 3959 -107 4005 1467
rect 4119 -107 4165 1467
rect 4279 -107 4325 1467
rect 4439 -107 4485 1467
rect 4599 -107 4645 1467
rect 4759 -107 4805 1467
rect 4919 -107 4965 1467
rect 5079 -107 5125 1467
rect 5239 -107 5285 1467
rect 5399 -107 5445 1467
rect 5559 -107 5605 1467
rect 5719 -107 5765 1467
rect 5879 -107 5925 1467
rect 6039 -107 6085 1467
rect 6199 -107 6245 1467
rect 6359 -107 6405 1467
rect 6519 -107 6565 1467
rect 6679 -107 6725 1467
rect 6839 -107 6885 1467
rect 6999 -107 7045 1467
rect 7159 -107 7205 1467
rect 7319 -107 7365 1467
rect 7479 -107 7525 1467
rect 7639 -107 7685 1467
rect 7799 -107 7845 1467
rect 7959 -107 8005 1467
<< psubdiff >>
rect 10803 -281 14379 -280
rect 8240 -301 14379 -281
rect 8240 -302 11861 -301
rect 8240 -308 9298 -302
rect 8240 -431 8323 -308
rect 8788 -425 9298 -308
rect 9763 -303 11861 -302
rect 9763 -425 10175 -303
rect 8788 -426 10175 -425
rect 10640 -307 11861 -303
rect 10640 -426 10886 -307
rect 8788 -430 10886 -426
rect 11351 -424 11861 -307
rect 12326 -302 14379 -301
rect 12326 -424 12738 -302
rect 11351 -425 12738 -424
rect 13203 -307 14379 -302
rect 13203 -425 13449 -307
rect 11351 -430 13449 -425
rect 13914 -430 14379 -307
rect 8788 -431 14379 -430
rect 8240 -450 14379 -431
rect 8240 -451 10803 -450
<< nsubdiff >>
rect 4740 1940 6191 1942
rect 2761 1926 7990 1940
rect 2761 1924 3752 1926
rect 2761 1788 2940 1924
rect 3385 1789 3752 1924
rect 4197 1789 4599 1926
rect 5044 1789 5560 1926
rect 6005 1789 6551 1926
rect 6996 1789 7483 1926
rect 7928 1789 7990 1926
rect 3385 1788 7990 1789
rect 2761 1776 7990 1788
rect 2761 1775 4778 1776
rect 6163 1775 7990 1776
<< psubdiffcont >>
rect 8323 -431 8788 -308
rect 9298 -425 9763 -302
rect 10175 -426 10640 -303
rect 10886 -430 11351 -307
rect 11861 -424 12326 -301
rect 12738 -425 13203 -302
rect 13449 -430 13914 -307
<< nsubdiffcont >>
rect 2940 1788 3385 1924
rect 3752 1789 4197 1926
rect 4599 1789 5044 1926
rect 5560 1789 6005 1926
rect 6551 1789 6996 1926
rect 7483 1789 7928 1926
<< polysilicon >>
rect 2914 1524 7930 1566
rect 2914 1480 2970 1524
rect 3074 1480 3130 1524
rect 3234 1480 3290 1524
rect 3394 1480 3450 1524
rect 3554 1480 3610 1524
rect 3714 1480 3770 1524
rect 3874 1480 3930 1524
rect 4034 1480 4090 1524
rect 4194 1480 4250 1524
rect 4354 1480 4410 1524
rect 4514 1480 4570 1524
rect 4674 1480 4730 1524
rect 4834 1480 4890 1524
rect 4994 1480 5050 1524
rect 5154 1480 5210 1524
rect 5314 1480 5370 1524
rect 5474 1480 5530 1524
rect 5634 1480 5690 1524
rect 5794 1480 5850 1524
rect 5954 1480 6010 1524
rect 6114 1480 6170 1524
rect 6274 1480 6330 1524
rect 6434 1480 6490 1524
rect 6594 1480 6650 1524
rect 6754 1480 6810 1524
rect 6914 1480 6970 1524
rect 7074 1480 7130 1524
rect 7234 1480 7290 1524
rect 7394 1480 7450 1524
rect 7554 1480 7610 1524
rect 7714 1480 7770 1524
rect 7874 1480 7930 1524
rect 8351 1519 10808 1560
rect 8352 1478 8408 1519
rect 8512 1478 8568 1519
rect 8672 1478 8728 1519
rect 8832 1478 8888 1519
rect 8992 1478 9048 1519
rect 9152 1478 9208 1519
rect 9312 1478 9368 1519
rect 9472 1478 9528 1519
rect 9632 1478 9688 1519
rect 9792 1478 9848 1519
rect 9952 1478 10008 1519
rect 10112 1478 10168 1519
rect 10272 1478 10328 1519
rect 10432 1478 10488 1519
rect 10592 1478 10648 1519
rect 10752 1478 10808 1519
rect 11040 1517 13497 1561
rect 11041 1478 11097 1517
rect 11201 1478 11257 1517
rect 11361 1478 11417 1517
rect 11521 1478 11577 1517
rect 11681 1478 11737 1517
rect 11841 1478 11897 1517
rect 12001 1478 12057 1517
rect 12161 1478 12217 1517
rect 12321 1478 12377 1517
rect 12481 1478 12537 1517
rect 12641 1478 12697 1517
rect 12801 1478 12857 1517
rect 12961 1478 13017 1517
rect 13121 1478 13177 1517
rect 13281 1478 13337 1517
rect 13441 1478 13497 1517
rect 13732 1513 14270 1561
rect 13732 1478 13788 1513
rect 13892 1478 13948 1513
rect 14052 1478 14108 1513
rect 14212 1478 14268 1513
rect 2914 -164 2970 -120
rect 3074 -164 3130 -120
rect 3234 -164 3290 -120
rect 3394 -164 3450 -120
rect 3554 -164 3610 -120
rect 3714 -164 3770 -120
rect 3874 -164 3930 -120
rect 4034 -164 4090 -120
rect 4194 -164 4250 -120
rect 4354 -164 4410 -120
rect 4514 -164 4570 -120
rect 4674 -164 4730 -120
rect 4834 -164 4890 -120
rect 4994 -164 5050 -120
rect 5154 -164 5210 -120
rect 5314 -164 5370 -120
rect 5474 -164 5530 -120
rect 5634 -164 5690 -120
rect 5794 -164 5850 -120
rect 5954 -164 6010 -120
rect 6114 -164 6170 -120
rect 6274 -164 6330 -120
rect 6434 -164 6490 -120
rect 6594 -164 6650 -120
rect 6754 -164 6810 -120
rect 6914 -164 6970 -120
rect 7074 -164 7130 -120
rect 7234 -164 7290 -120
rect 7394 -164 7450 -120
rect 7554 -164 7610 -120
rect 7714 -164 7770 -120
rect 7874 -164 7930 -120
rect 8352 -166 8408 -122
rect 8512 -166 8568 -122
rect 8672 -166 8728 -122
rect 8832 -166 8888 -122
rect 8992 -166 9048 -122
rect 9152 -166 9208 -122
rect 9312 -166 9368 -122
rect 9472 -166 9528 -122
rect 9632 -166 9688 -122
rect 9792 -166 9848 -122
rect 9952 -166 10008 -122
rect 10112 -166 10168 -122
rect 10272 -166 10328 -122
rect 10432 -166 10488 -122
rect 10592 -166 10648 -122
rect 10752 -166 10808 -122
rect 11041 -166 11097 -122
rect 11201 -166 11257 -122
rect 11361 -166 11417 -122
rect 11521 -166 11577 -122
rect 11681 -166 11737 -122
rect 11841 -166 11897 -122
rect 12001 -166 12057 -122
rect 12161 -166 12217 -122
rect 12321 -166 12377 -122
rect 12481 -166 12537 -122
rect 12641 -166 12697 -122
rect 12801 -166 12857 -122
rect 12961 -166 13017 -122
rect 13121 -166 13177 -122
rect 13281 -166 13337 -122
rect 13441 -166 13497 -122
rect 13732 -166 13788 -122
rect 13892 -166 13948 -122
rect 14052 -166 14108 -122
rect 14212 -166 14268 -122
<< metal1 >>
rect 2761 1926 7990 1940
rect 2761 1924 3752 1926
rect 2761 1788 2940 1924
rect 3385 1789 3752 1924
rect 4197 1789 4599 1926
rect 5044 1789 5560 1926
rect 6005 1789 6551 1926
rect 6996 1789 7483 1926
rect 7928 1789 7990 1926
rect 3385 1788 7990 1789
rect 2761 1775 7990 1788
rect 2839 1468 2885 1478
rect 2839 1467 2892 1468
rect 2885 1455 2892 1467
rect 2885 1386 2892 1400
rect 2999 1467 3045 1478
rect 2839 -118 2885 -107
rect 3159 1467 3205 1478
rect 3319 1467 3365 1478
rect 3205 1451 3212 1465
rect 3045 -4 3052 9
rect 3045 -89 3052 -76
rect 2999 -118 3045 -107
rect 3205 1382 3212 1396
rect 3159 -118 3205 -107
rect 3479 1467 3525 1478
rect 3639 1467 3685 1478
rect 3525 1447 3534 1462
rect 3533 1392 3534 1447
rect 3365 -2 3372 11
rect 3371 -74 3372 -2
rect 3365 -87 3372 -74
rect 3319 -118 3365 -107
rect 3525 1379 3534 1392
rect 3479 -118 3525 -107
rect 3799 1467 3845 1478
rect 3959 1467 4005 1478
rect 3845 1452 3852 1466
rect 3851 1397 3852 1452
rect 3685 -3 3692 10
rect 3685 -88 3692 -75
rect 3639 -118 3685 -107
rect 3845 1383 3852 1397
rect 3799 -118 3845 -107
rect 4119 1467 4165 1478
rect 4279 1467 4325 1478
rect 4165 1452 4172 1467
rect 4171 1397 4172 1452
rect 4005 -4 4012 9
rect 4005 -89 4012 -76
rect 3959 -118 4005 -107
rect 4165 1384 4172 1397
rect 4119 -118 4165 -107
rect 4439 1467 4485 1478
rect 4599 1467 4645 1478
rect 4485 1450 4492 1465
rect 4491 1395 4492 1450
rect 4325 -4 4333 8
rect 4332 -76 4333 -4
rect 4325 -90 4333 -76
rect 4279 -118 4325 -107
rect 4485 1382 4492 1395
rect 4439 -118 4485 -107
rect 4759 1467 4805 1478
rect 4919 1467 4965 1478
rect 4805 1449 4812 1462
rect 4811 1394 4812 1449
rect 4645 -4 4653 9
rect 4652 -76 4653 -4
rect 4645 -89 4653 -76
rect 4599 -118 4645 -107
rect 4805 1379 4812 1394
rect 4759 -118 4805 -107
rect 5079 1467 5125 1478
rect 5239 1467 5285 1478
rect 5125 1450 5132 1464
rect 4965 8 4971 9
rect 4965 -3 4973 8
rect 4971 -75 4973 -3
rect 4965 -90 4973 -75
rect 4919 -118 4965 -107
rect 5125 1381 5132 1395
rect 5079 -118 5125 -107
rect 5399 1467 5445 1478
rect 5559 1467 5605 1478
rect 5445 1449 5452 1462
rect 5451 1394 5452 1449
rect 5285 -1 5294 12
rect 5291 -73 5294 -1
rect 5285 -86 5294 -73
rect 5239 -118 5285 -107
rect 5445 1379 5452 1394
rect 5399 -118 5445 -107
rect 5719 1467 5765 1478
rect 5879 1467 5925 1478
rect 5765 1451 5772 1464
rect 5605 -3 5613 12
rect 5612 -75 5613 -3
rect 5605 -86 5613 -75
rect 5605 -87 5612 -86
rect 5559 -118 5605 -107
rect 5765 1381 5772 1396
rect 5719 -118 5765 -107
rect 6039 1467 6085 1478
rect 6199 1467 6245 1478
rect 6085 1450 6092 1462
rect 5925 -3 5933 11
rect 5931 -75 5933 -3
rect 5925 -87 5933 -75
rect 5879 -118 5925 -107
rect 6085 1379 6092 1395
rect 6039 -118 6085 -107
rect 6359 1467 6405 1478
rect 6519 1467 6565 1478
rect 6405 1449 6412 1463
rect 6245 -2 6253 10
rect 6251 -74 6253 -2
rect 6245 -88 6253 -74
rect 6199 -118 6245 -107
rect 6405 1380 6412 1394
rect 6359 -118 6405 -107
rect 6679 1467 6725 1478
rect 6839 1467 6885 1478
rect 6725 1449 6733 1462
rect 6732 1394 6733 1449
rect 6565 -2 6572 11
rect 6565 -87 6572 -74
rect 6519 -118 6565 -107
rect 6725 1379 6733 1394
rect 6679 -118 6725 -107
rect 6999 1467 7045 1478
rect 7159 1467 7205 1478
rect 7045 1448 7052 1463
rect 6885 -2 6893 12
rect 6892 -74 6893 -2
rect 6885 -86 6893 -74
rect 6839 -118 6885 -107
rect 7045 1380 7052 1393
rect 7158 -86 7159 12
rect 7319 1467 7365 1478
rect 7479 1467 7525 1478
rect 7365 1449 7372 1464
rect 7205 -3 7211 12
rect 6999 -118 7045 -107
rect 7205 -87 7211 -75
rect 7159 -118 7205 -107
rect 7365 1381 7372 1394
rect 7319 -118 7365 -107
rect 7639 1467 7685 1478
rect 7799 1467 7845 1478
rect 7685 1447 7692 1463
rect 7525 -4 7533 10
rect 7531 -76 7533 -4
rect 7525 -88 7533 -76
rect 7479 -118 7525 -107
rect 7685 1380 7692 1392
rect 7639 -118 7685 -107
rect 7959 1467 8005 1478
rect 8005 1448 8012 1466
rect 7845 -2 7853 12
rect 7851 -74 7853 -2
rect 7845 -86 7853 -74
rect 7799 -118 7845 -107
rect 8005 1381 8012 1393
rect 8277 1465 8323 1476
rect 7959 -118 8005 -107
rect 8437 1465 8483 1476
rect 8323 1308 8331 1320
rect 8323 1216 8331 1228
rect 8277 -120 8323 -109
rect 8597 1465 8643 1476
rect 8757 1465 8803 1476
rect 8643 1308 8651 1320
rect 8649 1228 8651 1308
rect 8483 -7 8492 5
rect 8491 -79 8492 -7
rect 8483 -90 8492 -79
rect 8483 -91 8491 -90
rect 8437 -120 8483 -109
rect 8643 1216 8651 1228
rect 8597 -120 8643 -109
rect 8917 1465 8963 1476
rect 9077 1465 9123 1476
rect 8963 1308 8971 1320
rect 8969 1228 8971 1308
rect 8803 -8 8812 6
rect 8810 -80 8812 -8
rect 8803 -94 8812 -80
rect 8757 -120 8803 -109
rect 8963 1216 8971 1228
rect 8917 -120 8963 -109
rect 9237 1465 9283 1476
rect 9397 1465 9443 1476
rect 9283 1308 9291 1320
rect 9290 1228 9291 1308
rect 9123 -10 9134 5
rect 9131 -82 9134 -10
rect 9123 -95 9134 -82
rect 9077 -120 9123 -109
rect 9283 1216 9291 1228
rect 9237 -120 9283 -109
rect 9557 1465 9603 1476
rect 9717 1465 9763 1476
rect 9603 1306 9611 1318
rect 9610 1226 9611 1306
rect 9443 -8 9452 6
rect 9450 -80 9452 -8
rect 9443 -94 9452 -80
rect 9397 -120 9443 -109
rect 9603 1213 9611 1226
rect 9557 -120 9603 -109
rect 9877 1465 9923 1476
rect 10037 1465 10083 1476
rect 9923 1306 9931 1318
rect 9930 1226 9931 1306
rect 9763 -8 9773 6
rect 9772 -80 9773 -8
rect 9763 -94 9773 -80
rect 9717 -120 9763 -109
rect 9923 1213 9931 1226
rect 10032 -8 10037 5
rect 10197 1465 10243 1476
rect 10357 1465 10403 1476
rect 10243 1307 10251 1319
rect 10250 1227 10251 1307
rect 10083 -8 10092 5
rect 10032 -80 10036 -8
rect 10089 -80 10092 -8
rect 10032 -95 10037 -80
rect 9877 -120 9923 -109
rect 10083 -95 10092 -80
rect 10037 -120 10083 -109
rect 10243 1214 10251 1227
rect 10197 -120 10243 -109
rect 10517 1465 10563 1476
rect 10677 1465 10723 1476
rect 10563 1307 10571 1319
rect 10570 1227 10571 1307
rect 10403 -9 10413 6
rect 10412 -81 10413 -9
rect 10403 -96 10413 -81
rect 10357 -120 10403 -109
rect 10563 1214 10571 1227
rect 10517 -120 10563 -109
rect 10837 1465 10883 1476
rect 10966 1465 11012 1476
rect 10883 1307 10891 1320
rect 10889 1227 10891 1307
rect 10723 -9 10735 6
rect 10730 -81 10735 -9
rect 10723 -96 10735 -81
rect 10677 -120 10723 -109
rect 10883 1215 10891 1227
rect 10837 -120 10883 -109
rect 11126 1465 11172 1476
rect 11012 1120 11020 1133
rect 11012 1015 11020 1030
rect 10966 -120 11012 -109
rect 11286 1465 11332 1476
rect 11446 1465 11492 1476
rect 11332 1110 11343 1123
rect 11340 1020 11343 1110
rect 11172 -8 11189 7
rect 11181 -80 11189 -8
rect 11172 -95 11189 -80
rect 11126 -120 11172 -109
rect 11332 1005 11343 1020
rect 11286 -120 11332 -109
rect 11606 1465 11652 1476
rect 11766 1465 11812 1476
rect 11652 1109 11666 1123
rect 11660 1019 11666 1109
rect 11492 -8 11509 7
rect 11500 -80 11509 -8
rect 11492 -95 11509 -80
rect 11446 -120 11492 -109
rect 11652 1005 11666 1019
rect 11606 -120 11652 -109
rect 11926 1465 11972 1476
rect 12086 1465 12132 1476
rect 11972 1109 11982 1123
rect 11980 1019 11982 1109
rect 11812 -9 11832 7
rect 11819 -81 11832 -9
rect 11812 -95 11832 -81
rect 11766 -120 11812 -109
rect 11972 1005 11982 1019
rect 12081 -10 12086 4
rect 12246 1465 12292 1476
rect 12406 1465 12452 1476
rect 12292 1110 12303 1123
rect 12301 1020 12303 1110
rect 12132 -10 12141 4
rect 12081 -82 12085 -10
rect 12138 -82 12141 -10
rect 12081 -94 12086 -82
rect 11926 -120 11972 -109
rect 12132 -94 12141 -82
rect 12086 -120 12132 -109
rect 12292 1005 12303 1020
rect 12246 -120 12292 -109
rect 12566 1465 12612 1476
rect 12726 1465 12772 1476
rect 12612 1109 12624 1123
rect 12620 1019 12624 1109
rect 12452 -7 12461 9
rect 12459 -79 12461 -7
rect 12452 -93 12461 -79
rect 12406 -120 12452 -109
rect 12612 1005 12624 1019
rect 12566 -120 12612 -109
rect 12886 1465 12932 1476
rect 13046 1465 13092 1476
rect 12932 1111 12944 1126
rect 12941 1021 12944 1111
rect 12772 -8 12787 8
rect 12781 -80 12787 -8
rect 12772 -94 12787 -80
rect 12726 -120 12772 -109
rect 12932 1008 12944 1021
rect 12886 -120 12932 -109
rect 13206 1465 13252 1476
rect 13366 1465 13412 1476
rect 13252 1111 13265 1125
rect 13261 1021 13265 1111
rect 13092 -8 13107 6
rect 13100 -80 13107 -8
rect 13092 -96 13107 -80
rect 13046 -120 13092 -109
rect 13252 1007 13265 1021
rect 13206 -120 13252 -109
rect 13526 1465 13572 1476
rect 13657 1465 13703 1476
rect 13572 1110 13582 1123
rect 13581 1020 13582 1110
rect 13412 -8 13421 6
rect 13419 -80 13421 -8
rect 13412 -96 13421 -80
rect 13366 -120 13412 -109
rect 13572 1005 13582 1020
rect 13526 -120 13572 -109
rect 13817 1465 13863 1476
rect 13703 769 13714 787
rect 13711 666 13714 769
rect 13703 652 13714 666
rect 13657 -120 13703 -109
rect 13977 1465 14023 1476
rect 14137 1465 14183 1476
rect 14023 769 14038 789
rect 14030 666 14038 769
rect 13863 -7 13874 6
rect 13870 -79 13874 -7
rect 13863 -96 13874 -79
rect 13817 -120 13863 -109
rect 14023 654 14038 666
rect 13977 -120 14023 -109
rect 14297 1465 14343 1476
rect 14343 778 14356 795
rect 14350 675 14356 778
rect 14183 -5 14195 8
rect 14192 -77 14195 -5
rect 14183 -94 14195 -77
rect 14137 -120 14183 -109
rect 14343 660 14356 675
rect 14297 -120 14343 -109
rect 10803 -281 14379 -280
rect 8240 -301 14379 -281
rect 8240 -302 11861 -301
rect 8240 -308 9298 -302
rect 8240 -431 8323 -308
rect 8788 -425 9298 -308
rect 9763 -303 11861 -302
rect 9763 -425 10175 -303
rect 8788 -426 10175 -425
rect 10640 -307 11861 -303
rect 10640 -426 10886 -307
rect 8788 -430 10886 -426
rect 11351 -424 11861 -307
rect 12326 -302 14379 -301
rect 12326 -424 12738 -302
rect 11351 -425 12738 -424
rect 13203 -307 14379 -302
rect 13203 -425 13449 -307
rect 11351 -430 13449 -425
rect 13914 -430 14379 -307
rect 8788 -431 14379 -430
rect 8240 -450 14379 -431
rect 8240 -451 10803 -450
<< via1 >>
rect 2840 1400 2885 1455
rect 2885 1400 2892 1455
rect 3160 1396 3205 1451
rect 3205 1396 3212 1451
rect 3000 -76 3045 -4
rect 3045 -76 3052 -4
rect 3481 1392 3525 1447
rect 3525 1392 3533 1447
rect 3319 -74 3365 -2
rect 3365 -74 3371 -2
rect 3799 1397 3845 1452
rect 3845 1397 3851 1452
rect 3640 -75 3685 -3
rect 3685 -75 3692 -3
rect 4119 1397 4165 1452
rect 4165 1397 4171 1452
rect 3960 -76 4005 -4
rect 4005 -76 4012 -4
rect 4439 1395 4485 1450
rect 4485 1395 4491 1450
rect 4280 -76 4325 -4
rect 4325 -76 4332 -4
rect 4759 1394 4805 1449
rect 4805 1394 4811 1449
rect 4600 -76 4645 -4
rect 4645 -76 4652 -4
rect 5080 1395 5125 1450
rect 5125 1395 5132 1450
rect 4919 -75 4965 -3
rect 4965 -75 4971 -3
rect 5399 1394 5445 1449
rect 5445 1394 5451 1449
rect 5239 -73 5285 -1
rect 5285 -73 5291 -1
rect 5720 1396 5765 1451
rect 5765 1396 5772 1451
rect 5560 -75 5605 -3
rect 5605 -75 5612 -3
rect 6040 1395 6085 1450
rect 6085 1395 6092 1450
rect 5879 -75 5925 -3
rect 5925 -75 5931 -3
rect 6360 1394 6405 1449
rect 6405 1394 6412 1449
rect 6199 -74 6245 -2
rect 6245 -74 6251 -2
rect 6680 1394 6725 1449
rect 6725 1394 6732 1449
rect 6520 -74 6565 -2
rect 6565 -74 6572 -2
rect 7000 1393 7045 1448
rect 7045 1393 7052 1448
rect 6840 -74 6885 -2
rect 6885 -74 6892 -2
rect 7320 1394 7365 1449
rect 7365 1394 7372 1449
rect 7159 -75 7205 -3
rect 7205 -75 7211 -3
rect 7640 1392 7685 1447
rect 7685 1392 7692 1447
rect 7479 -76 7525 -4
rect 7525 -76 7531 -4
rect 7960 1393 8005 1448
rect 8005 1393 8012 1448
rect 7799 -74 7845 -2
rect 7845 -74 7851 -2
rect 8279 1228 8323 1308
rect 8323 1228 8331 1308
rect 8597 1228 8643 1308
rect 8643 1228 8649 1308
rect 8438 -79 8483 -7
rect 8483 -79 8491 -7
rect 8917 1228 8963 1308
rect 8963 1228 8969 1308
rect 8757 -80 8803 -8
rect 8803 -80 8810 -8
rect 9238 1228 9283 1308
rect 9283 1228 9290 1308
rect 9078 -82 9123 -10
rect 9123 -82 9131 -10
rect 9558 1226 9603 1306
rect 9603 1226 9610 1306
rect 9397 -80 9443 -8
rect 9443 -80 9450 -8
rect 9878 1226 9923 1306
rect 9923 1226 9930 1306
rect 9719 -80 9763 -8
rect 9763 -80 9772 -8
rect 10198 1227 10243 1307
rect 10243 1227 10250 1307
rect 10036 -80 10037 -8
rect 10037 -80 10083 -8
rect 10083 -80 10089 -8
rect 10518 1227 10563 1307
rect 10563 1227 10570 1307
rect 10359 -81 10403 -9
rect 10403 -81 10412 -9
rect 10837 1227 10883 1307
rect 10883 1227 10889 1307
rect 10677 -81 10723 -9
rect 10723 -81 10730 -9
rect 10966 1030 11012 1120
rect 11012 1030 11020 1120
rect 11286 1020 11332 1110
rect 11332 1020 11340 1110
rect 11128 -80 11172 -8
rect 11172 -80 11181 -8
rect 11606 1019 11652 1109
rect 11652 1019 11660 1109
rect 11447 -80 11492 -8
rect 11492 -80 11500 -8
rect 11926 1019 11972 1109
rect 11972 1019 11980 1109
rect 11766 -81 11812 -9
rect 11812 -81 11819 -9
rect 12247 1020 12292 1110
rect 12292 1020 12301 1110
rect 12085 -82 12086 -10
rect 12086 -82 12132 -10
rect 12132 -82 12138 -10
rect 12566 1019 12612 1109
rect 12612 1019 12620 1109
rect 12406 -79 12452 -7
rect 12452 -79 12459 -7
rect 12887 1021 12932 1111
rect 12932 1021 12941 1111
rect 12728 -80 12772 -8
rect 12772 -80 12781 -8
rect 13207 1021 13252 1111
rect 13252 1021 13261 1111
rect 13047 -80 13092 -8
rect 13092 -80 13100 -8
rect 13527 1020 13572 1110
rect 13572 1020 13581 1110
rect 13366 -80 13412 -8
rect 13412 -80 13419 -8
rect 13659 666 13703 769
rect 13703 666 13711 769
rect 13978 666 14023 769
rect 14023 666 14030 769
rect 13817 -79 13863 -7
rect 13863 -79 13870 -7
rect 14298 675 14343 778
rect 14343 675 14350 778
rect 14139 -77 14183 -5
rect 14183 -77 14192 -5
<< metal2 >>
rect 2833 1455 8024 1467
rect 2833 1400 2840 1455
rect 2892 1452 8024 1455
rect 2892 1451 3799 1452
rect 2892 1400 3160 1451
rect 2833 1396 3160 1400
rect 3212 1447 3799 1451
rect 3212 1396 3481 1447
rect 2833 1392 3481 1396
rect 3533 1397 3799 1447
rect 3851 1397 4119 1452
rect 4171 1451 8024 1452
rect 4171 1450 5720 1451
rect 4171 1397 4439 1450
rect 3533 1395 4439 1397
rect 4491 1449 5080 1450
rect 4491 1395 4759 1449
rect 3533 1394 4759 1395
rect 4811 1395 5080 1449
rect 5132 1449 5720 1450
rect 5132 1395 5399 1449
rect 4811 1394 5399 1395
rect 5451 1396 5720 1449
rect 5772 1450 8024 1451
rect 5772 1396 6040 1450
rect 5451 1395 6040 1396
rect 6092 1449 8024 1450
rect 6092 1395 6360 1449
rect 5451 1394 6360 1395
rect 6412 1394 6680 1449
rect 6732 1448 7320 1449
rect 6732 1394 7000 1448
rect 3533 1393 7000 1394
rect 7052 1394 7320 1448
rect 7372 1448 8024 1449
rect 7372 1447 7960 1448
rect 7372 1394 7640 1447
rect 7052 1393 7640 1394
rect 3533 1392 7640 1393
rect 7692 1393 7960 1447
rect 8012 1393 8024 1448
rect 7692 1392 8024 1393
rect 2833 1387 8024 1392
rect 8274 1308 10893 1321
rect 8274 1228 8279 1308
rect 8331 1228 8597 1308
rect 8649 1228 8917 1308
rect 8969 1228 9238 1308
rect 9290 1307 10893 1308
rect 9290 1306 10198 1307
rect 9290 1228 9558 1306
rect 8274 1226 9558 1228
rect 9610 1226 9878 1306
rect 9930 1227 10198 1306
rect 10250 1227 10518 1307
rect 10570 1227 10837 1307
rect 10889 1227 10893 1307
rect 9930 1226 10893 1227
rect 8274 1215 10893 1226
rect 10954 1120 13593 1123
rect 10954 1030 10966 1120
rect 11020 1111 13593 1120
rect 11020 1110 12887 1111
rect 11020 1030 11286 1110
rect 10954 1020 11286 1030
rect 11340 1109 12247 1110
rect 11340 1020 11606 1109
rect 10954 1019 11606 1020
rect 11660 1019 11926 1109
rect 11980 1020 12247 1109
rect 12301 1109 12887 1110
rect 12301 1020 12566 1109
rect 11980 1019 12566 1020
rect 12620 1021 12887 1109
rect 12941 1021 13207 1111
rect 13261 1110 13593 1111
rect 13261 1021 13527 1110
rect 12620 1020 13527 1021
rect 13581 1020 13593 1110
rect 12620 1019 13593 1020
rect 10954 1017 13593 1019
rect 13651 778 14361 789
rect 13651 769 14298 778
rect 13651 666 13659 769
rect 13711 666 13978 769
rect 14030 675 14298 769
rect 14350 675 14361 778
rect 14030 666 14361 675
rect 13651 652 14361 666
rect 2982 3 7882 5
rect 2982 -1 14358 3
rect 2982 -2 5239 -1
rect 2982 -4 3319 -2
rect 2982 -76 3000 -4
rect 3052 -74 3319 -4
rect 3371 -3 5239 -2
rect 3371 -74 3640 -3
rect 3052 -75 3640 -74
rect 3692 -4 4919 -3
rect 3692 -75 3960 -4
rect 3052 -76 3960 -75
rect 4012 -76 4280 -4
rect 4332 -76 4600 -4
rect 4652 -75 4919 -4
rect 4971 -73 5239 -3
rect 5291 -2 14358 -1
rect 5291 -3 6199 -2
rect 5291 -73 5560 -3
rect 4971 -75 5560 -73
rect 5612 -75 5879 -3
rect 5931 -74 6199 -3
rect 6251 -74 6520 -2
rect 6572 -74 6840 -2
rect 6892 -3 7799 -2
rect 6892 -74 7159 -3
rect 5931 -75 7159 -74
rect 7211 -4 7799 -3
rect 7211 -75 7479 -4
rect 4652 -76 7479 -75
rect 7531 -74 7799 -4
rect 7851 -5 14358 -2
rect 7851 -7 14139 -5
rect 7851 -74 8438 -7
rect 7531 -76 8438 -74
rect 2982 -79 8438 -76
rect 8491 -8 12406 -7
rect 8491 -79 8757 -8
rect 2982 -80 8757 -79
rect 8810 -10 9397 -8
rect 8810 -80 9078 -10
rect 2982 -82 9078 -80
rect 9131 -80 9397 -10
rect 9450 -80 9719 -8
rect 9772 -80 10036 -8
rect 10089 -9 11128 -8
rect 10089 -80 10359 -9
rect 9131 -81 10359 -80
rect 10412 -81 10677 -9
rect 10730 -80 11128 -9
rect 11181 -80 11447 -8
rect 11500 -9 12406 -8
rect 11500 -80 11766 -9
rect 10730 -81 11766 -80
rect 11819 -10 12406 -9
rect 11819 -81 12085 -10
rect 9131 -82 12085 -81
rect 12138 -79 12406 -10
rect 12459 -8 13817 -7
rect 12459 -79 12728 -8
rect 12138 -80 12728 -79
rect 12781 -80 13047 -8
rect 13100 -80 13366 -8
rect 13419 -79 13817 -8
rect 13870 -77 14139 -7
rect 14192 -77 14358 -5
rect 13870 -79 14358 -77
rect 13419 -80 14358 -79
rect 12138 -82 14358 -80
rect 2982 -89 14358 -82
rect 7874 -91 14358 -89
<< labels >>
flabel metal1 9581 -406 12346 -309 0 FreeSans 320 0 0 0 VSS
port 11 nsew
flabel metal1 4295 1806 7060 1903 0 FreeSans 320 0 0 0 VDD
port 8 nsew
flabel metal2 13802 678 14267 760 0 FreeSans 320 0 0 0 VIN
port 3 nsew
flabel metal2 11223 1040 13113 1097 0 FreeSans 320 0 0 0 VREF_GND
port 2 nsew
flabel metal2 8931 1235 10821 1292 0 FreeSans 320 0 0 0 VCM
port 1 nsew
flabel metal2 4732 -85 10945 -25 0 FreeSans 320 0 0 0 Cbtm
port 7 nsew
flabel metal2 2834 1390 7951 1464 0 FreeSans 320 0 0 0 VREF
port 4 nsew
flabel polysilicon 13740 1516 14266 1557 0 FreeSans 320 0 0 0 EN_VIN
port 10 nsew
flabel polysilicon 11048 1520 13493 1557 0 FreeSans 320 0 0 0 EN_VSS
port 9 nsew
flabel polysilicon 8351 1520 10806 1558 0 FreeSans 320 0 0 0 EN_VCM
port 5 nsew
flabel polysilicon 2914 1524 7930 1566 0 FreeSans 320 0 0 0 EN_VREF_Z
port 6 nsew
<< end >>
