magic
tech gf180mcuD
timestamp 1756801411
<< metal2 >>
rect 0 42 40 43
rect 0 36 1 42
rect 7 36 33 42
rect 39 36 40 42
rect 0 7 40 36
rect 0 1 1 7
rect 7 1 33 7
rect 39 1 40 7
rect 0 0 40 1
<< via2 >>
rect 1 36 7 42
rect 33 36 39 42
rect 1 1 7 7
rect 33 1 39 7
<< metal3 >>
rect 0 42 40 43
rect 0 36 1 42
rect 7 37 33 42
rect 7 36 8 37
rect 0 35 8 36
rect 32 36 33 37
rect 39 36 40 42
rect 32 35 40 36
rect 0 8 6 35
rect 33 34 40 35
rect 14 29 17 31
rect 12 25 17 29
rect 23 29 26 31
rect 23 25 28 29
rect 12 18 28 25
rect 12 14 17 18
rect 14 12 17 14
rect 23 14 28 18
rect 23 12 26 14
rect 34 8 40 34
rect 0 7 8 8
rect 0 1 1 7
rect 7 6 8 7
rect 32 7 40 8
rect 32 6 33 7
rect 7 1 33 6
rect 39 1 40 7
rect 0 0 40 1
<< via3 >>
rect 17 25 23 31
rect 17 12 23 18
<< metal4 >>
rect 17 31 23 44
rect 16 25 17 30
rect 23 25 24 30
rect 16 18 24 25
rect 16 12 17 18
rect 23 12 24 18
rect 17 -2 23 12
<< end >>
