magic
tech gf180mcuD
magscale 1 10
timestamp 1757727097
<< nwell >>
rect -778 -930 778 930
<< pmos >>
rect -604 -800 -544 800
rect -440 -800 -380 800
rect -276 -800 -216 800
rect -112 -800 -52 800
rect 52 -800 112 800
rect 216 -800 276 800
rect 380 -800 440 800
rect 544 -800 604 800
<< pdiff >>
rect -692 787 -604 800
rect -692 -787 -679 787
rect -633 -787 -604 787
rect -692 -800 -604 -787
rect -544 787 -440 800
rect -544 -787 -515 787
rect -469 -787 -440 787
rect -544 -800 -440 -787
rect -380 787 -276 800
rect -380 -787 -351 787
rect -305 -787 -276 787
rect -380 -800 -276 -787
rect -216 787 -112 800
rect -216 -787 -187 787
rect -141 -787 -112 787
rect -216 -800 -112 -787
rect -52 787 52 800
rect -52 -787 -23 787
rect 23 -787 52 787
rect -52 -800 52 -787
rect 112 787 216 800
rect 112 -787 141 787
rect 187 -787 216 787
rect 112 -800 216 -787
rect 276 787 380 800
rect 276 -787 305 787
rect 351 -787 380 787
rect 276 -800 380 -787
rect 440 787 544 800
rect 440 -787 469 787
rect 515 -787 544 787
rect 440 -800 544 -787
rect 604 787 692 800
rect 604 -787 633 787
rect 679 -787 692 787
rect 604 -800 692 -787
<< pdiffc >>
rect -679 -787 -633 787
rect -515 -787 -469 787
rect -351 -787 -305 787
rect -187 -787 -141 787
rect -23 -787 23 787
rect 141 -787 187 787
rect 305 -787 351 787
rect 469 -787 515 787
rect 633 -787 679 787
<< polysilicon >>
rect -604 800 -544 844
rect -440 800 -380 844
rect -276 800 -216 844
rect -112 800 -52 844
rect 52 800 112 844
rect 216 800 276 844
rect 380 800 440 844
rect 544 800 604 844
rect -604 -844 -544 -800
rect -440 -844 -380 -800
rect -276 -844 -216 -800
rect -112 -844 -52 -800
rect 52 -844 112 -800
rect 216 -844 276 -800
rect 380 -844 440 -800
rect 544 -844 604 -800
<< metal1 >>
rect -679 787 -633 798
rect -679 -798 -633 -787
rect -515 787 -469 798
rect -515 -798 -469 -787
rect -351 787 -305 798
rect -351 -798 -305 -787
rect -187 787 -141 798
rect -187 -798 -141 -787
rect -23 787 23 798
rect -23 -798 23 -787
rect 141 787 187 798
rect 141 -798 187 -787
rect 305 787 351 798
rect 305 -798 351 -787
rect 469 787 515 798
rect 469 -798 515 -787
rect 633 787 679 798
rect 633 -798 679 -787
<< properties >>
string gencell pfet_03v3
string library gf180mcu
string parameters w 8 l 0.3 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {pfet_03v3 pfet_06v0}
<< end >>
