magic
tech gf180mcuD
magscale 1 10
timestamp 1757859342
<< nwell >>
rect 441 724 521 844
<< pwell >>
rect 436 -44 522 59
rect 3 -101 968 -44
rect 3 -104 522 -101
rect 436 -210 522 -104
<< psubdiff >>
rect 434 21 524 60
rect 434 -60 449 21
rect 436 -176 449 -60
rect 508 -60 524 21
rect 508 -176 522 -60
rect 436 -210 522 -176
<< nsubdiff >>
rect 441 826 521 844
rect 441 737 455 826
rect 504 737 521 826
rect 441 724 521 737
rect 430 -894 544 -876
rect 430 -981 450 -894
rect 513 -981 544 -894
rect 430 -996 544 -981
<< psubdiffcont >>
rect 449 -176 508 21
<< nsubdiffcont >>
rect 455 737 504 826
rect 450 -981 513 -894
<< metal1 >>
rect 441 826 521 844
rect 441 737 455 826
rect 504 737 521 826
rect 441 724 521 737
rect 260 248 313 383
rect 318 353 560 430
rect 1197 223 1280 239
rect 1197 141 1208 223
rect 1269 141 1280 223
rect 1197 132 1280 141
rect 863 107 935 114
rect 434 21 524 60
rect 434 -44 449 21
rect 3 -104 449 -44
rect 436 -176 449 -104
rect 508 -44 524 21
rect 962 -44 1290 -22
rect 508 -101 1290 -44
rect 508 -176 522 -101
rect 436 -210 522 -176
rect 962 -212 1290 -101
rect 259 -372 267 -307
rect 259 -387 318 -372
rect 614 -459 685 -439
rect 614 -560 624 -459
rect 676 -560 685 -459
rect 614 -574 685 -560
rect 430 -894 544 -876
rect 430 -981 450 -894
rect 513 -981 544 -894
rect 430 -996 544 -981
<< via1 >>
rect 872 120 930 225
rect 1208 141 1269 223
rect 267 -372 319 -272
rect 624 -560 676 -459
<< metal2 >>
rect 863 235 935 238
rect 855 225 935 235
rect 855 200 872 225
rect 256 129 872 200
rect 256 12 324 129
rect 855 120 872 129
rect 930 120 935 225
rect 1197 223 1280 239
rect 1197 141 1208 223
rect 1269 141 1280 223
rect 1197 135 1280 141
rect 855 103 935 120
rect 1195 33 1280 135
rect 256 -272 322 12
rect 614 -36 1290 33
rect 256 -372 267 -272
rect 319 -372 322 -272
rect 256 -384 322 -372
rect 615 -439 683 -36
rect 1195 -38 1280 -36
rect 613 -459 686 -439
rect 613 -560 624 -459
rect 676 -560 686 -459
rect 613 -574 686 -560
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gf180mcu_fd_sc_mcu7t5v0__inv_1_0 ~/conda-gf180mcu-env/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1757859342
transform 1 0 0 0 1 0
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gf180mcu_fd_sc_mcu7t5v0__inv_1_1
timestamp 1757859342
transform 1 0 3 0 -1 -152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gf180mcu_fd_sc_mcu7t5v0__inv_1_2
timestamp 1757859342
transform 1 0 518 0 -1 -152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  gf180mcu_fd_sc_mcu7t5v0__nand3_1_0 ~/conda-gf180mcu-env/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1757859342
transform 1 0 507 0 1 0
box -86 -86 870 870
<< end >>
