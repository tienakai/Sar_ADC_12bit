magic
tech gf180mcuD
magscale 1 10
timestamp 1757226667
<< nwell >>
rect -2682 -930 2682 930
<< pmos >>
rect -2508 -800 -2452 800
rect -2348 -800 -2292 800
rect -2188 -800 -2132 800
rect -2028 -800 -1972 800
rect -1868 -800 -1812 800
rect -1708 -800 -1652 800
rect -1548 -800 -1492 800
rect -1388 -800 -1332 800
rect -1228 -800 -1172 800
rect -1068 -800 -1012 800
rect -908 -800 -852 800
rect -748 -800 -692 800
rect -588 -800 -532 800
rect -428 -800 -372 800
rect -268 -800 -212 800
rect -108 -800 -52 800
rect 52 -800 108 800
rect 212 -800 268 800
rect 372 -800 428 800
rect 532 -800 588 800
rect 692 -800 748 800
rect 852 -800 908 800
rect 1012 -800 1068 800
rect 1172 -800 1228 800
rect 1332 -800 1388 800
rect 1492 -800 1548 800
rect 1652 -800 1708 800
rect 1812 -800 1868 800
rect 1972 -800 2028 800
rect 2132 -800 2188 800
rect 2292 -800 2348 800
rect 2452 -800 2508 800
<< pdiff >>
rect -2596 787 -2508 800
rect -2596 -787 -2583 787
rect -2537 -787 -2508 787
rect -2596 -800 -2508 -787
rect -2452 787 -2348 800
rect -2452 -787 -2423 787
rect -2377 -787 -2348 787
rect -2452 -800 -2348 -787
rect -2292 787 -2188 800
rect -2292 -787 -2263 787
rect -2217 -787 -2188 787
rect -2292 -800 -2188 -787
rect -2132 787 -2028 800
rect -2132 -787 -2103 787
rect -2057 -787 -2028 787
rect -2132 -800 -2028 -787
rect -1972 787 -1868 800
rect -1972 -787 -1943 787
rect -1897 -787 -1868 787
rect -1972 -800 -1868 -787
rect -1812 787 -1708 800
rect -1812 -787 -1783 787
rect -1737 -787 -1708 787
rect -1812 -800 -1708 -787
rect -1652 787 -1548 800
rect -1652 -787 -1623 787
rect -1577 -787 -1548 787
rect -1652 -800 -1548 -787
rect -1492 787 -1388 800
rect -1492 -787 -1463 787
rect -1417 -787 -1388 787
rect -1492 -800 -1388 -787
rect -1332 787 -1228 800
rect -1332 -787 -1303 787
rect -1257 -787 -1228 787
rect -1332 -800 -1228 -787
rect -1172 787 -1068 800
rect -1172 -787 -1143 787
rect -1097 -787 -1068 787
rect -1172 -800 -1068 -787
rect -1012 787 -908 800
rect -1012 -787 -983 787
rect -937 -787 -908 787
rect -1012 -800 -908 -787
rect -852 787 -748 800
rect -852 -787 -823 787
rect -777 -787 -748 787
rect -852 -800 -748 -787
rect -692 787 -588 800
rect -692 -787 -663 787
rect -617 -787 -588 787
rect -692 -800 -588 -787
rect -532 787 -428 800
rect -532 -787 -503 787
rect -457 -787 -428 787
rect -532 -800 -428 -787
rect -372 787 -268 800
rect -372 -787 -343 787
rect -297 -787 -268 787
rect -372 -800 -268 -787
rect -212 787 -108 800
rect -212 -787 -183 787
rect -137 -787 -108 787
rect -212 -800 -108 -787
rect -52 787 52 800
rect -52 -787 -23 787
rect 23 -787 52 787
rect -52 -800 52 -787
rect 108 787 212 800
rect 108 -787 137 787
rect 183 -787 212 787
rect 108 -800 212 -787
rect 268 787 372 800
rect 268 -787 297 787
rect 343 -787 372 787
rect 268 -800 372 -787
rect 428 787 532 800
rect 428 -787 457 787
rect 503 -787 532 787
rect 428 -800 532 -787
rect 588 787 692 800
rect 588 -787 617 787
rect 663 -787 692 787
rect 588 -800 692 -787
rect 748 787 852 800
rect 748 -787 777 787
rect 823 -787 852 787
rect 748 -800 852 -787
rect 908 787 1012 800
rect 908 -787 937 787
rect 983 -787 1012 787
rect 908 -800 1012 -787
rect 1068 787 1172 800
rect 1068 -787 1097 787
rect 1143 -787 1172 787
rect 1068 -800 1172 -787
rect 1228 787 1332 800
rect 1228 -787 1257 787
rect 1303 -787 1332 787
rect 1228 -800 1332 -787
rect 1388 787 1492 800
rect 1388 -787 1417 787
rect 1463 -787 1492 787
rect 1388 -800 1492 -787
rect 1548 787 1652 800
rect 1548 -787 1577 787
rect 1623 -787 1652 787
rect 1548 -800 1652 -787
rect 1708 787 1812 800
rect 1708 -787 1737 787
rect 1783 -787 1812 787
rect 1708 -800 1812 -787
rect 1868 787 1972 800
rect 1868 -787 1897 787
rect 1943 -787 1972 787
rect 1868 -800 1972 -787
rect 2028 787 2132 800
rect 2028 -787 2057 787
rect 2103 -787 2132 787
rect 2028 -800 2132 -787
rect 2188 787 2292 800
rect 2188 -787 2217 787
rect 2263 -787 2292 787
rect 2188 -800 2292 -787
rect 2348 787 2452 800
rect 2348 -787 2377 787
rect 2423 -787 2452 787
rect 2348 -800 2452 -787
rect 2508 787 2596 800
rect 2508 -787 2537 787
rect 2583 -787 2596 787
rect 2508 -800 2596 -787
<< pdiffc >>
rect -2583 -787 -2537 787
rect -2423 -787 -2377 787
rect -2263 -787 -2217 787
rect -2103 -787 -2057 787
rect -1943 -787 -1897 787
rect -1783 -787 -1737 787
rect -1623 -787 -1577 787
rect -1463 -787 -1417 787
rect -1303 -787 -1257 787
rect -1143 -787 -1097 787
rect -983 -787 -937 787
rect -823 -787 -777 787
rect -663 -787 -617 787
rect -503 -787 -457 787
rect -343 -787 -297 787
rect -183 -787 -137 787
rect -23 -787 23 787
rect 137 -787 183 787
rect 297 -787 343 787
rect 457 -787 503 787
rect 617 -787 663 787
rect 777 -787 823 787
rect 937 -787 983 787
rect 1097 -787 1143 787
rect 1257 -787 1303 787
rect 1417 -787 1463 787
rect 1577 -787 1623 787
rect 1737 -787 1783 787
rect 1897 -787 1943 787
rect 2057 -787 2103 787
rect 2217 -787 2263 787
rect 2377 -787 2423 787
rect 2537 -787 2583 787
<< polysilicon >>
rect -2508 800 -2452 844
rect -2348 800 -2292 844
rect -2188 800 -2132 844
rect -2028 800 -1972 844
rect -1868 800 -1812 844
rect -1708 800 -1652 844
rect -1548 800 -1492 844
rect -1388 800 -1332 844
rect -1228 800 -1172 844
rect -1068 800 -1012 844
rect -908 800 -852 844
rect -748 800 -692 844
rect -588 800 -532 844
rect -428 800 -372 844
rect -268 800 -212 844
rect -108 800 -52 844
rect 52 800 108 844
rect 212 800 268 844
rect 372 800 428 844
rect 532 800 588 844
rect 692 800 748 844
rect 852 800 908 844
rect 1012 800 1068 844
rect 1172 800 1228 844
rect 1332 800 1388 844
rect 1492 800 1548 844
rect 1652 800 1708 844
rect 1812 800 1868 844
rect 1972 800 2028 844
rect 2132 800 2188 844
rect 2292 800 2348 844
rect 2452 800 2508 844
rect -2508 -844 -2452 -800
rect -2348 -844 -2292 -800
rect -2188 -844 -2132 -800
rect -2028 -844 -1972 -800
rect -1868 -844 -1812 -800
rect -1708 -844 -1652 -800
rect -1548 -844 -1492 -800
rect -1388 -844 -1332 -800
rect -1228 -844 -1172 -800
rect -1068 -844 -1012 -800
rect -908 -844 -852 -800
rect -748 -844 -692 -800
rect -588 -844 -532 -800
rect -428 -844 -372 -800
rect -268 -844 -212 -800
rect -108 -844 -52 -800
rect 52 -844 108 -800
rect 212 -844 268 -800
rect 372 -844 428 -800
rect 532 -844 588 -800
rect 692 -844 748 -800
rect 852 -844 908 -800
rect 1012 -844 1068 -800
rect 1172 -844 1228 -800
rect 1332 -844 1388 -800
rect 1492 -844 1548 -800
rect 1652 -844 1708 -800
rect 1812 -844 1868 -800
rect 1972 -844 2028 -800
rect 2132 -844 2188 -800
rect 2292 -844 2348 -800
rect 2452 -844 2508 -800
<< metal1 >>
rect -2583 787 -2537 798
rect -2583 -798 -2537 -787
rect -2423 787 -2377 798
rect -2423 -798 -2377 -787
rect -2263 787 -2217 798
rect -2263 -798 -2217 -787
rect -2103 787 -2057 798
rect -2103 -798 -2057 -787
rect -1943 787 -1897 798
rect -1943 -798 -1897 -787
rect -1783 787 -1737 798
rect -1783 -798 -1737 -787
rect -1623 787 -1577 798
rect -1623 -798 -1577 -787
rect -1463 787 -1417 798
rect -1463 -798 -1417 -787
rect -1303 787 -1257 798
rect -1303 -798 -1257 -787
rect -1143 787 -1097 798
rect -1143 -798 -1097 -787
rect -983 787 -937 798
rect -983 -798 -937 -787
rect -823 787 -777 798
rect -823 -798 -777 -787
rect -663 787 -617 798
rect -663 -798 -617 -787
rect -503 787 -457 798
rect -503 -798 -457 -787
rect -343 787 -297 798
rect -343 -798 -297 -787
rect -183 787 -137 798
rect -183 -798 -137 -787
rect -23 787 23 798
rect -23 -798 23 -787
rect 137 787 183 798
rect 137 -798 183 -787
rect 297 787 343 798
rect 297 -798 343 -787
rect 457 787 503 798
rect 457 -798 503 -787
rect 617 787 663 798
rect 617 -798 663 -787
rect 777 787 823 798
rect 777 -798 823 -787
rect 937 787 983 798
rect 937 -798 983 -787
rect 1097 787 1143 798
rect 1097 -798 1143 -787
rect 1257 787 1303 798
rect 1257 -798 1303 -787
rect 1417 787 1463 798
rect 1417 -798 1463 -787
rect 1577 787 1623 798
rect 1577 -798 1623 -787
rect 1737 787 1783 798
rect 1737 -798 1783 -787
rect 1897 787 1943 798
rect 1897 -798 1943 -787
rect 2057 787 2103 798
rect 2057 -798 2103 -787
rect 2217 787 2263 798
rect 2217 -798 2263 -787
rect 2377 787 2423 798
rect 2377 -798 2423 -787
rect 2537 787 2583 798
rect 2537 -798 2583 -787
<< properties >>
string gencell pfet_03v3
string library gf180mcu
string parameters w 8 l 0.280 m 1 nf 32 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {pfet_03v3 pfet_06v0}
<< end >>
