* SPICE3 file created from CADC_12bit.ext - technology: gf180mcuD

.option scale=5n

C0 C3 Ctop 6.53425f
C1 C3 VSS 0.80455f
C2 C3 C4 9.03513f
C3 C1 Ctop 1.63151f
C4 C2 C3 2.543f
C5 C6 C7 24.8148f
C6 C1 VSS 0.80509f
C7 C6 C5 18.8713f
C8 C2 C1 0.49308f
C9 C8 Ctop 0.20953p
C10 VSS Ctop 12.58842f
C11 C4 Ctop 13.06933f
C12 C0_dummy Ctop 0.81454f
C13 C2 Ctop 3.26508f
C14 C8 VSS 8.01912f
C15 C1 C0 1.01398f
C16 C4 VSS 2.40734f
C17 C0_dummy VSS 0.80437f
C18 C2 VSS 0.80437f
C19 C0_dummy C4 0
C20 C2 C4 1.96397f
C21 C3 C5 0
C22 C0_dummy C2 2.24296f
C23 C0 Ctop 0.81584f
C24 C9 Ctop 0.42017p
C25 C10 Ctop 0.84269p
C26 VSS C0 0.80567f
C27 C9 C8 51.1857f
C28 C9 VSS 9.62097f
C29 C4 C0 0
C30 VSS C10 16.12827f
C31 C0_dummy C0 1.22151f
C32 C2 C0 0.80983f
C33 Ctop C7 0.10473p
C34 C5 Ctop 26.16638f
C35 C8 C7 33.4464f
C36 VSS C7 4.8113f
C37 C6 Ctop 52.34919f
C38 VSS C5 1.60626f
C39 C6 VSS 3.20887f
C40 C4 C5 12.4366f
C41 C2 C5 0
C42 C3 C1 2.98144f
C43 C9 C10 71.4828f
C44 C7 0 16.13945f
C45 Ctop 0 0.3306p
C46 C5 0 4.159f
C47 C0 0 0.38811f
C48 C10 0 0.22588p
C49 VSS 0 77.72894f
C50 C1 0 0.49878f
C51 C8 0 29.74999f
C52 C4 0 2.561f
C53 C9 0 61.18403f
C54 C3 0 1.19934f
C55 C6 0 8.31239f
C56 C2 0 0.72683f
C57 C0_dummy 0 0.3817f
