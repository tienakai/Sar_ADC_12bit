magic
tech gf180mcuD
magscale 1 10
timestamp 1757727608
<< error_p >>
rect -227 -48 -181 48
rect -23 -48 23 48
rect 181 -48 227 48
<< pwell >>
rect -264 -118 264 118
<< nmos >>
rect -152 -50 -52 50
rect 52 -50 152 50
<< ndiff >>
rect -240 37 -152 50
rect -240 -37 -227 37
rect -181 -37 -152 37
rect -240 -50 -152 -37
rect -52 37 52 50
rect -52 -37 -23 37
rect 23 -37 52 37
rect -52 -50 52 -37
rect 152 37 240 50
rect 152 -37 181 37
rect 227 -37 240 37
rect 152 -50 240 -37
<< ndiffc >>
rect -227 -37 -181 37
rect -23 -37 23 37
rect 181 -37 227 37
<< polysilicon >>
rect -152 50 -52 94
rect 52 50 152 94
rect -152 -94 -52 -50
rect 52 -94 152 -50
<< metal1 >>
rect -227 37 -181 48
rect -227 -48 -181 -37
rect -23 37 23 48
rect -23 -48 23 -37
rect 181 37 227 48
rect 181 -48 227 -37
<< properties >>
string gencell nfet_03v3
string library gf180mcu
string parameters w 0.5 l 0.5 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt}
<< end >>
