magic
tech gf180mcuD
magscale 1 10
timestamp 1757388344
<< nwell >>
rect 1886 720 2003 840
rect 1992 569 2048 625
<< psubdiff >>
rect 1877 42 2008 56
rect 1877 -51 1901 42
rect 1987 -51 2008 42
rect 1877 -64 2008 -51
<< nsubdiff >>
rect 1886 826 2003 840
rect 1886 734 1906 826
rect 1985 734 2003 826
rect 1886 720 2003 734
<< psubdiffcont >>
rect 1901 -51 1987 42
<< nsubdiffcont >>
rect 1906 734 1985 826
<< metal1 >>
rect 1886 826 2003 840
rect 1886 734 1906 826
rect 1985 734 2003 826
rect 1886 720 2003 734
rect 3672 643 3682 658
rect 3672 531 3682 556
rect 1877 42 2008 56
rect 1877 -51 1901 42
rect 1987 -51 2008 42
rect 1877 -64 2008 -51
<< via1 >>
rect 1506 541 1568 631
rect 3629 556 3682 643
rect 624 367 711 420
rect 2368 357 2438 416
rect 2791 380 2843 467
rect 260 244 347 297
<< metal2 >>
rect -108 631 1581 691
rect 3621 643 3698 654
rect 3621 632 3629 643
rect 2788 631 3629 632
rect -108 611 1506 631
rect 1499 541 1506 611
rect 1568 605 1581 631
rect 2113 630 3629 631
rect 1978 625 3629 630
rect 1739 605 1807 606
rect 1568 541 1807 605
rect 1978 569 1992 625
rect 2048 569 3629 625
rect 1978 561 3629 569
rect 1978 560 2797 561
rect 1978 559 2662 560
rect 3621 556 3629 561
rect 3682 630 3698 643
rect 3682 560 4101 630
rect 3682 556 3698 560
rect 3621 545 3698 556
rect 1499 526 1807 541
rect 610 428 1510 435
rect 610 420 1410 428
rect 610 367 624 420
rect 711 367 1410 420
rect 610 361 1410 367
rect 1487 361 1510 428
rect 610 355 1510 361
rect 1739 420 1807 526
rect 2775 467 2854 479
rect 2334 420 2451 423
rect 1739 416 2451 420
rect 1739 357 2368 416
rect 2438 357 2451 416
rect 2775 380 2791 467
rect 2843 433 2854 467
rect 2843 432 2927 433
rect 2843 380 4099 432
rect 2775 370 4099 380
rect 612 353 724 355
rect 1739 352 2451 357
rect 2334 351 2451 352
rect 248 309 360 310
rect -112 297 364 309
rect -112 244 260 297
rect 347 244 364 297
rect -112 240 364 244
rect 248 232 360 240
<< via2 >>
rect 1992 569 2048 625
rect 1410 361 1487 428
<< metal3 >>
rect 1979 625 2056 639
rect 1979 569 1992 625
rect 2048 569 2056 625
rect 1979 557 2056 569
rect 1398 437 1506 438
rect 1980 437 2055 557
rect 1398 433 2055 437
rect 1398 428 2051 433
rect 1398 361 1410 428
rect 1487 361 2051 428
rect 1398 350 2051 361
use gf180mcu_fd_sc_mcu7t5v0__and2_4  gf180mcu_fd_sc_mcu7t5v0__and2_4_0 ~/conda-gf180mcu-env/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 -4 0 1 -4
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__or2_4  gf180mcu_fd_sc_mcu7t5v0__or2_4_0 ~/conda-gf180mcu-env/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 1991 0 1 -4
box -86 -86 2102 870
<< end >>
