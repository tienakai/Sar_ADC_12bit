magic
tech gf180mcuD
magscale 1 10
timestamp 1757325240
<< nwell >>
rect 5830 12794 8634 14978
<< pwell >>
rect 2498 12794 5830 14978
<< nmos >>
rect 2610 13054 2666 14654
rect 2770 13054 2826 14654
rect 3062 13054 3118 14654
rect 3222 13054 3278 14654
rect 3382 13054 3438 14654
rect 3542 13054 3598 14654
rect 3702 13054 3758 14654
rect 3862 13054 3918 14654
rect 4022 13054 4078 14654
rect 4182 13054 4238 14654
rect 4480 13054 4536 14654
rect 4640 13054 4696 14654
rect 4800 13054 4856 14654
rect 4960 13054 5016 14654
rect 5120 13054 5176 14654
rect 5280 13054 5336 14654
rect 5440 13054 5496 14654
rect 5600 13054 5656 14654
<< pmos >>
rect 6004 13054 6060 14654
rect 6164 13054 6220 14654
rect 6324 13054 6380 14654
rect 6484 13054 6540 14654
rect 6644 13054 6700 14654
rect 6804 13054 6860 14654
rect 6964 13054 7020 14654
rect 7124 13054 7180 14654
rect 7284 13054 7340 14654
rect 7444 13054 7500 14654
rect 7604 13054 7660 14654
rect 7764 13054 7820 14654
rect 7924 13054 7980 14654
rect 8084 13054 8140 14654
rect 8244 13054 8300 14654
rect 8404 13054 8460 14654
<< ndiff >>
rect 2522 14641 2610 14654
rect 2522 13067 2535 14641
rect 2581 13067 2610 14641
rect 2522 13054 2610 13067
rect 2666 14641 2770 14654
rect 2666 13067 2695 14641
rect 2741 13067 2770 14641
rect 2666 13054 2770 13067
rect 2826 14641 2914 14654
rect 2826 13067 2855 14641
rect 2901 13067 2914 14641
rect 2826 13054 2914 13067
rect 2974 14641 3062 14654
rect 2974 13067 2987 14641
rect 3033 13067 3062 14641
rect 2974 13054 3062 13067
rect 3118 14641 3222 14654
rect 3118 13067 3147 14641
rect 3193 13067 3222 14641
rect 3118 13054 3222 13067
rect 3278 14641 3382 14654
rect 3278 13067 3307 14641
rect 3353 13067 3382 14641
rect 3278 13054 3382 13067
rect 3438 14641 3542 14654
rect 3438 13067 3467 14641
rect 3513 13067 3542 14641
rect 3438 13054 3542 13067
rect 3598 14641 3702 14654
rect 3598 13067 3627 14641
rect 3673 13067 3702 14641
rect 3598 13054 3702 13067
rect 3758 14641 3862 14654
rect 3758 13067 3787 14641
rect 3833 13067 3862 14641
rect 3758 13054 3862 13067
rect 3918 14641 4022 14654
rect 3918 13067 3947 14641
rect 3993 13067 4022 14641
rect 3918 13054 4022 13067
rect 4078 14641 4182 14654
rect 4078 13067 4107 14641
rect 4153 13067 4182 14641
rect 4078 13054 4182 13067
rect 4238 14641 4326 14654
rect 4238 13067 4267 14641
rect 4313 13067 4326 14641
rect 4238 13054 4326 13067
rect 4392 14641 4480 14654
rect 4392 13067 4405 14641
rect 4451 13067 4480 14641
rect 4392 13054 4480 13067
rect 4536 14641 4640 14654
rect 4536 13067 4565 14641
rect 4611 13067 4640 14641
rect 4536 13054 4640 13067
rect 4696 14641 4800 14654
rect 4696 13067 4725 14641
rect 4771 13067 4800 14641
rect 4696 13054 4800 13067
rect 4856 14641 4960 14654
rect 4856 13067 4885 14641
rect 4931 13067 4960 14641
rect 4856 13054 4960 13067
rect 5016 14641 5120 14654
rect 5016 13067 5045 14641
rect 5091 13067 5120 14641
rect 5016 13054 5120 13067
rect 5176 14641 5280 14654
rect 5176 13067 5205 14641
rect 5251 13067 5280 14641
rect 5176 13054 5280 13067
rect 5336 14641 5440 14654
rect 5336 13067 5365 14641
rect 5411 13067 5440 14641
rect 5336 13054 5440 13067
rect 5496 14641 5600 14654
rect 5496 13067 5525 14641
rect 5571 13067 5600 14641
rect 5496 13054 5600 13067
rect 5656 14641 5744 14654
rect 5656 13067 5685 14641
rect 5731 13067 5744 14641
rect 5656 13054 5744 13067
<< pdiff >>
rect 5916 14641 6004 14654
rect 5916 13067 5929 14641
rect 5975 13067 6004 14641
rect 5916 13054 6004 13067
rect 6060 14641 6164 14654
rect 6060 13067 6089 14641
rect 6135 13067 6164 14641
rect 6060 13054 6164 13067
rect 6220 14641 6324 14654
rect 6220 13067 6249 14641
rect 6295 13067 6324 14641
rect 6220 13054 6324 13067
rect 6380 14641 6484 14654
rect 6380 13067 6409 14641
rect 6455 13067 6484 14641
rect 6380 13054 6484 13067
rect 6540 14641 6644 14654
rect 6540 13067 6569 14641
rect 6615 13067 6644 14641
rect 6540 13054 6644 13067
rect 6700 14641 6804 14654
rect 6700 13067 6729 14641
rect 6775 13067 6804 14641
rect 6700 13054 6804 13067
rect 6860 14641 6964 14654
rect 6860 13067 6889 14641
rect 6935 13067 6964 14641
rect 6860 13054 6964 13067
rect 7020 14641 7124 14654
rect 7020 13067 7049 14641
rect 7095 13067 7124 14641
rect 7020 13054 7124 13067
rect 7180 14641 7284 14654
rect 7180 13067 7209 14641
rect 7255 13067 7284 14641
rect 7180 13054 7284 13067
rect 7340 14641 7444 14654
rect 7340 13067 7369 14641
rect 7415 13067 7444 14641
rect 7340 13054 7444 13067
rect 7500 14641 7604 14654
rect 7500 13067 7529 14641
rect 7575 13067 7604 14641
rect 7500 13054 7604 13067
rect 7660 14641 7764 14654
rect 7660 13067 7689 14641
rect 7735 13067 7764 14641
rect 7660 13054 7764 13067
rect 7820 14641 7924 14654
rect 7820 13067 7849 14641
rect 7895 13067 7924 14641
rect 7820 13054 7924 13067
rect 7980 14641 8084 14654
rect 7980 13067 8009 14641
rect 8055 13067 8084 14641
rect 7980 13054 8084 13067
rect 8140 14641 8244 14654
rect 8140 13067 8169 14641
rect 8215 13067 8244 14641
rect 8140 13054 8244 13067
rect 8300 14641 8404 14654
rect 8300 13067 8329 14641
rect 8375 13067 8404 14641
rect 8300 13054 8404 13067
rect 8460 14641 8548 14654
rect 8460 13067 8489 14641
rect 8535 13067 8548 14641
rect 8460 13054 8548 13067
<< ndiffc >>
rect 2535 13067 2581 14641
rect 2695 13067 2741 14641
rect 2855 13067 2901 14641
rect 2987 13067 3033 14641
rect 3147 13067 3193 14641
rect 3307 13067 3353 14641
rect 3467 13067 3513 14641
rect 3627 13067 3673 14641
rect 3787 13067 3833 14641
rect 3947 13067 3993 14641
rect 4107 13067 4153 14641
rect 4267 13067 4313 14641
rect 4405 13067 4451 14641
rect 4565 13067 4611 14641
rect 4725 13067 4771 14641
rect 4885 13067 4931 14641
rect 5045 13067 5091 14641
rect 5205 13067 5251 14641
rect 5365 13067 5411 14641
rect 5525 13067 5571 14641
rect 5685 13067 5731 14641
<< pdiffc >>
rect 5929 13067 5975 14641
rect 6089 13067 6135 14641
rect 6249 13067 6295 14641
rect 6409 13067 6455 14641
rect 6569 13067 6615 14641
rect 6729 13067 6775 14641
rect 6889 13067 6935 14641
rect 7049 13067 7095 14641
rect 7209 13067 7255 14641
rect 7369 13067 7415 14641
rect 7529 13067 7575 14641
rect 7689 13067 7735 14641
rect 7849 13067 7895 14641
rect 8009 13067 8055 14641
rect 8169 13067 8215 14641
rect 8329 13067 8375 14641
rect 8489 13067 8535 14641
<< psubdiff >>
rect 2559 12953 2699 12984
rect 2559 12863 2587 12953
rect 2677 12863 2699 12953
rect 2559 12836 2699 12863
<< nsubdiff >>
rect 5902 14887 6051 14915
rect 5902 14797 5928 14887
rect 6018 14797 6051 14887
rect 5902 14771 6051 14797
<< psubdiffcont >>
rect 2587 12863 2677 12953
<< nsubdiffcont >>
rect 5928 14797 6018 14887
<< polysilicon >>
rect 2610 14698 2826 14734
rect 2610 14654 2666 14698
rect 2770 14654 2826 14698
rect 3062 14698 4238 14734
rect 3062 14654 3118 14698
rect 3222 14654 3278 14698
rect 3382 14654 3438 14698
rect 3542 14654 3598 14698
rect 3702 14654 3758 14698
rect 3862 14654 3918 14698
rect 4022 14654 4078 14698
rect 4182 14654 4238 14698
rect 4480 14698 5656 14734
rect 4480 14654 4536 14698
rect 4640 14654 4696 14698
rect 4800 14654 4856 14698
rect 4960 14654 5016 14698
rect 5120 14654 5176 14698
rect 5280 14654 5336 14698
rect 5440 14654 5496 14698
rect 5600 14654 5656 14698
rect 6004 14698 8460 14734
rect 6004 14654 6060 14698
rect 6164 14654 6220 14698
rect 6324 14654 6380 14698
rect 6484 14654 6540 14698
rect 6644 14654 6700 14698
rect 6804 14654 6860 14698
rect 6964 14654 7020 14698
rect 7124 14654 7180 14698
rect 7284 14654 7340 14698
rect 7444 14654 7500 14698
rect 7604 14654 7660 14698
rect 7764 14654 7820 14698
rect 7924 14654 7980 14698
rect 8084 14654 8140 14698
rect 8244 14654 8300 14698
rect 8404 14654 8460 14698
rect 2610 13010 2666 13054
rect 2770 13010 2826 13054
rect 3062 13010 3118 13054
rect 3222 13010 3278 13054
rect 3382 13010 3438 13054
rect 3542 13010 3598 13054
rect 3702 13010 3758 13054
rect 3862 13010 3918 13054
rect 4022 13010 4078 13054
rect 4182 13010 4238 13054
rect 4480 13010 4536 13054
rect 4640 13010 4696 13054
rect 4800 13010 4856 13054
rect 4960 13010 5016 13054
rect 5120 13010 5176 13054
rect 5280 13010 5336 13054
rect 5440 13010 5496 13054
rect 5600 13010 5656 13054
rect 6004 13010 6060 13054
rect 6164 13010 6220 13054
rect 6324 13010 6380 13054
rect 6484 13010 6540 13054
rect 6644 13010 6700 13054
rect 6804 13010 6860 13054
rect 6964 13010 7020 13054
rect 7124 13010 7180 13054
rect 7284 13010 7340 13054
rect 7444 13010 7500 13054
rect 7604 13010 7660 13054
rect 7764 13010 7820 13054
rect 7924 13010 7980 13054
rect 8084 13010 8140 13054
rect 8244 13010 8300 13054
rect 8404 13010 8460 13054
<< metal1 >>
rect 2570 14887 8590 14932
rect 2570 14797 5928 14887
rect 6018 14797 8590 14887
rect 2570 14756 8590 14797
rect 2520 14641 2596 14652
rect 2520 14640 2535 14641
rect 2581 14640 2596 14641
rect 2520 14588 2532 14640
rect 2584 14588 2596 14640
rect 2520 14584 2535 14588
rect 2581 14584 2596 14588
rect 2695 14641 2741 14652
rect 2535 13056 2581 13067
rect 2680 13120 2695 13124
rect 2840 14641 2916 14652
rect 2840 14640 2855 14641
rect 2901 14640 2916 14641
rect 2840 14588 2852 14640
rect 2904 14588 2916 14640
rect 2840 14584 2855 14588
rect 2741 13120 2756 13124
rect 2680 13068 2692 13120
rect 2744 13068 2756 13120
rect 2680 13067 2695 13068
rect 2741 13067 2756 13068
rect 2680 13056 2756 13067
rect 2901 14584 2916 14588
rect 2972 14641 3048 14652
rect 2972 14640 2987 14641
rect 3033 14640 3048 14641
rect 2972 14588 2984 14640
rect 3036 14588 3048 14640
rect 2972 14584 2987 14588
rect 2855 13056 2901 13067
rect 3033 14584 3048 14588
rect 3147 14641 3193 14652
rect 2987 13056 3033 13067
rect 3132 13120 3147 13124
rect 3292 14641 3368 14652
rect 3292 14640 3307 14641
rect 3353 14640 3368 14641
rect 3292 14588 3304 14640
rect 3356 14588 3368 14640
rect 3292 14584 3307 14588
rect 3193 13120 3208 13124
rect 3132 13068 3144 13120
rect 3196 13068 3208 13120
rect 3132 13067 3147 13068
rect 3193 13067 3208 13068
rect 3132 13056 3208 13067
rect 3353 14584 3368 14588
rect 3467 14641 3513 14652
rect 3307 13056 3353 13067
rect 3452 13120 3467 13124
rect 3612 14641 3688 14652
rect 3612 14640 3627 14641
rect 3673 14640 3688 14641
rect 3612 14588 3624 14640
rect 3676 14588 3688 14640
rect 3612 14584 3627 14588
rect 3513 13120 3528 13124
rect 3452 13068 3464 13120
rect 3516 13068 3528 13120
rect 3452 13067 3467 13068
rect 3513 13067 3528 13068
rect 3452 13056 3528 13067
rect 3673 14584 3688 14588
rect 3787 14641 3833 14652
rect 3627 13056 3673 13067
rect 3772 13120 3787 13124
rect 3932 14641 4008 14652
rect 3932 14640 3947 14641
rect 3993 14640 4008 14641
rect 3932 14588 3944 14640
rect 3996 14588 4008 14640
rect 3932 14584 3947 14588
rect 3833 13120 3848 13124
rect 3772 13068 3784 13120
rect 3836 13068 3848 13120
rect 3772 13067 3787 13068
rect 3833 13067 3848 13068
rect 3772 13056 3848 13067
rect 3993 14584 4008 14588
rect 4107 14641 4153 14652
rect 3947 13056 3993 13067
rect 4092 13120 4107 13124
rect 4252 14641 4328 14652
rect 4252 14640 4267 14641
rect 4313 14640 4328 14641
rect 4252 14588 4264 14640
rect 4316 14588 4328 14640
rect 4252 14584 4267 14588
rect 4153 13120 4168 13124
rect 4092 13068 4104 13120
rect 4156 13068 4168 13120
rect 4092 13067 4107 13068
rect 4153 13067 4168 13068
rect 4092 13056 4168 13067
rect 4313 14584 4328 14588
rect 4390 14641 4466 14652
rect 4390 14640 4405 14641
rect 4451 14640 4466 14641
rect 4390 14588 4402 14640
rect 4454 14588 4466 14640
rect 4390 14584 4405 14588
rect 4267 13056 4313 13067
rect 4451 14584 4466 14588
rect 4565 14641 4611 14652
rect 4405 13056 4451 13067
rect 4550 13120 4565 13124
rect 4710 14641 4786 14652
rect 4710 14640 4725 14641
rect 4771 14640 4786 14641
rect 4710 14588 4722 14640
rect 4774 14588 4786 14640
rect 4710 14584 4725 14588
rect 4611 13120 4626 13124
rect 4550 13068 4562 13120
rect 4614 13068 4626 13120
rect 4550 13067 4565 13068
rect 4611 13067 4626 13068
rect 4550 13056 4626 13067
rect 4771 14584 4786 14588
rect 4885 14641 4931 14652
rect 4725 13056 4771 13067
rect 4870 13120 4885 13124
rect 5030 14641 5106 14652
rect 5030 14640 5045 14641
rect 5091 14640 5106 14641
rect 5030 14588 5042 14640
rect 5094 14588 5106 14640
rect 5030 14584 5045 14588
rect 4931 13120 4946 13124
rect 4870 13068 4882 13120
rect 4934 13068 4946 13120
rect 4870 13067 4885 13068
rect 4931 13067 4946 13068
rect 4870 13056 4946 13067
rect 5091 14584 5106 14588
rect 5205 14641 5251 14652
rect 5045 13056 5091 13067
rect 5190 13120 5205 13124
rect 5350 14641 5426 14652
rect 5350 14640 5365 14641
rect 5411 14640 5426 14641
rect 5350 14588 5362 14640
rect 5414 14588 5426 14640
rect 5350 14584 5365 14588
rect 5251 13120 5266 13124
rect 5190 13068 5202 13120
rect 5254 13068 5266 13120
rect 5190 13067 5205 13068
rect 5251 13067 5266 13068
rect 5190 13056 5266 13067
rect 5411 14584 5426 14588
rect 5525 14641 5571 14652
rect 5365 13056 5411 13067
rect 5510 13120 5525 13124
rect 5670 14641 5746 14652
rect 5670 14640 5685 14641
rect 5731 14640 5746 14641
rect 5670 14588 5682 14640
rect 5734 14588 5746 14640
rect 5670 14584 5685 14588
rect 5571 13120 5586 13124
rect 5510 13068 5522 13120
rect 5574 13068 5586 13120
rect 5510 13067 5525 13068
rect 5571 13067 5586 13068
rect 5510 13056 5586 13067
rect 5731 14584 5746 14588
rect 5914 14641 5990 14652
rect 5914 14640 5929 14641
rect 5975 14640 5990 14641
rect 5914 14588 5926 14640
rect 5978 14588 5990 14640
rect 5914 14584 5929 14588
rect 5685 13056 5731 13067
rect 5975 14584 5990 14588
rect 6089 14641 6135 14652
rect 5929 13056 5975 13067
rect 6074 13120 6089 13124
rect 6234 14641 6310 14652
rect 6234 14640 6249 14641
rect 6295 14640 6310 14641
rect 6234 14588 6246 14640
rect 6298 14588 6310 14640
rect 6234 14584 6249 14588
rect 6135 13120 6150 13124
rect 6074 13068 6086 13120
rect 6138 13068 6150 13120
rect 6074 13067 6089 13068
rect 6135 13067 6150 13068
rect 6074 13056 6150 13067
rect 6295 14584 6310 14588
rect 6409 14641 6455 14652
rect 6249 13056 6295 13067
rect 6394 13120 6409 13124
rect 6554 14641 6630 14652
rect 6554 14640 6569 14641
rect 6615 14640 6630 14641
rect 6554 14588 6566 14640
rect 6618 14588 6630 14640
rect 6554 14584 6569 14588
rect 6455 13120 6470 13124
rect 6394 13068 6406 13120
rect 6458 13068 6470 13120
rect 6394 13067 6409 13068
rect 6455 13067 6470 13068
rect 6394 13056 6470 13067
rect 6615 14584 6630 14588
rect 6729 14641 6775 14652
rect 6569 13056 6615 13067
rect 6714 13120 6729 13124
rect 6874 14641 6950 14652
rect 6874 14640 6889 14641
rect 6935 14640 6950 14641
rect 6874 14588 6886 14640
rect 6938 14588 6950 14640
rect 6874 14584 6889 14588
rect 6775 13120 6790 13124
rect 6714 13068 6726 13120
rect 6778 13068 6790 13120
rect 6714 13067 6729 13068
rect 6775 13067 6790 13068
rect 6714 13056 6790 13067
rect 6935 14584 6950 14588
rect 7049 14641 7095 14652
rect 6889 13056 6935 13067
rect 7034 13120 7049 13124
rect 7194 14641 7270 14652
rect 7194 14640 7209 14641
rect 7255 14640 7270 14641
rect 7194 14588 7206 14640
rect 7258 14588 7270 14640
rect 7194 14584 7209 14588
rect 7095 13120 7110 13124
rect 7034 13068 7046 13120
rect 7098 13068 7110 13120
rect 7034 13067 7049 13068
rect 7095 13067 7110 13068
rect 7034 13056 7110 13067
rect 7255 14584 7270 14588
rect 7369 14641 7415 14652
rect 7209 13056 7255 13067
rect 7354 13120 7369 13124
rect 7514 14641 7590 14652
rect 7514 14640 7529 14641
rect 7575 14640 7590 14641
rect 7514 14588 7526 14640
rect 7578 14588 7590 14640
rect 7514 14584 7529 14588
rect 7415 13120 7430 13124
rect 7354 13068 7366 13120
rect 7418 13068 7430 13120
rect 7354 13067 7369 13068
rect 7415 13067 7430 13068
rect 7354 13056 7430 13067
rect 7575 14584 7590 14588
rect 7689 14641 7735 14652
rect 7529 13056 7575 13067
rect 7674 13120 7689 13124
rect 7834 14641 7910 14652
rect 7834 14640 7849 14641
rect 7895 14640 7910 14641
rect 7834 14588 7846 14640
rect 7898 14588 7910 14640
rect 7834 14584 7849 14588
rect 7735 13120 7750 13124
rect 7674 13068 7686 13120
rect 7738 13068 7750 13120
rect 7674 13067 7689 13068
rect 7735 13067 7750 13068
rect 7674 13056 7750 13067
rect 7895 14584 7910 14588
rect 8009 14641 8055 14652
rect 7849 13056 7895 13067
rect 7994 13120 8009 13124
rect 8154 14641 8230 14652
rect 8154 14640 8169 14641
rect 8215 14640 8230 14641
rect 8154 14588 8166 14640
rect 8218 14588 8230 14640
rect 8154 14584 8169 14588
rect 8055 13120 8070 13124
rect 7994 13068 8006 13120
rect 8058 13068 8070 13120
rect 7994 13067 8009 13068
rect 8055 13067 8070 13068
rect 7994 13056 8070 13067
rect 8215 14584 8230 14588
rect 8329 14641 8375 14652
rect 8169 13056 8215 13067
rect 8314 13120 8329 13124
rect 8475 14641 8551 14652
rect 8475 14640 8489 14641
rect 8535 14640 8551 14641
rect 8475 14588 8487 14640
rect 8539 14588 8551 14640
rect 8475 14584 8489 14588
rect 8375 13120 8390 13124
rect 8314 13068 8326 13120
rect 8378 13068 8390 13120
rect 8314 13067 8329 13068
rect 8375 13067 8390 13068
rect 8314 13056 8390 13067
rect 8535 14584 8551 14588
rect 8489 13056 8535 13067
rect 2502 12953 8607 13000
rect 2502 12863 2587 12953
rect 2677 12863 8607 12953
rect 2502 12824 8607 12863
<< via1 >>
rect 2532 14588 2535 14640
rect 2535 14588 2581 14640
rect 2581 14588 2584 14640
rect 2852 14588 2855 14640
rect 2855 14588 2901 14640
rect 2901 14588 2904 14640
rect 2692 13068 2695 13120
rect 2695 13068 2741 13120
rect 2741 13068 2744 13120
rect 2984 14588 2987 14640
rect 2987 14588 3033 14640
rect 3033 14588 3036 14640
rect 3304 14588 3307 14640
rect 3307 14588 3353 14640
rect 3353 14588 3356 14640
rect 3144 13068 3147 13120
rect 3147 13068 3193 13120
rect 3193 13068 3196 13120
rect 3624 14588 3627 14640
rect 3627 14588 3673 14640
rect 3673 14588 3676 14640
rect 3464 13068 3467 13120
rect 3467 13068 3513 13120
rect 3513 13068 3516 13120
rect 3944 14588 3947 14640
rect 3947 14588 3993 14640
rect 3993 14588 3996 14640
rect 3784 13068 3787 13120
rect 3787 13068 3833 13120
rect 3833 13068 3836 13120
rect 4264 14588 4267 14640
rect 4267 14588 4313 14640
rect 4313 14588 4316 14640
rect 4104 13068 4107 13120
rect 4107 13068 4153 13120
rect 4153 13068 4156 13120
rect 4402 14588 4405 14640
rect 4405 14588 4451 14640
rect 4451 14588 4454 14640
rect 4722 14588 4725 14640
rect 4725 14588 4771 14640
rect 4771 14588 4774 14640
rect 4562 13068 4565 13120
rect 4565 13068 4611 13120
rect 4611 13068 4614 13120
rect 5042 14588 5045 14640
rect 5045 14588 5091 14640
rect 5091 14588 5094 14640
rect 4882 13068 4885 13120
rect 4885 13068 4931 13120
rect 4931 13068 4934 13120
rect 5362 14588 5365 14640
rect 5365 14588 5411 14640
rect 5411 14588 5414 14640
rect 5202 13068 5205 13120
rect 5205 13068 5251 13120
rect 5251 13068 5254 13120
rect 5682 14588 5685 14640
rect 5685 14588 5731 14640
rect 5731 14588 5734 14640
rect 5522 13068 5525 13120
rect 5525 13068 5571 13120
rect 5571 13068 5574 13120
rect 5926 14588 5929 14640
rect 5929 14588 5975 14640
rect 5975 14588 5978 14640
rect 6246 14588 6249 14640
rect 6249 14588 6295 14640
rect 6295 14588 6298 14640
rect 6086 13068 6089 13120
rect 6089 13068 6135 13120
rect 6135 13068 6138 13120
rect 6566 14588 6569 14640
rect 6569 14588 6615 14640
rect 6615 14588 6618 14640
rect 6406 13068 6409 13120
rect 6409 13068 6455 13120
rect 6455 13068 6458 13120
rect 6886 14588 6889 14640
rect 6889 14588 6935 14640
rect 6935 14588 6938 14640
rect 6726 13068 6729 13120
rect 6729 13068 6775 13120
rect 6775 13068 6778 13120
rect 7206 14588 7209 14640
rect 7209 14588 7255 14640
rect 7255 14588 7258 14640
rect 7046 13068 7049 13120
rect 7049 13068 7095 13120
rect 7095 13068 7098 13120
rect 7526 14588 7529 14640
rect 7529 14588 7575 14640
rect 7575 14588 7578 14640
rect 7366 13068 7369 13120
rect 7369 13068 7415 13120
rect 7415 13068 7418 13120
rect 7846 14588 7849 14640
rect 7849 14588 7895 14640
rect 7895 14588 7898 14640
rect 7686 13068 7689 13120
rect 7689 13068 7735 13120
rect 7735 13068 7738 13120
rect 8166 14588 8169 14640
rect 8169 14588 8215 14640
rect 8215 14588 8218 14640
rect 8006 13068 8009 13120
rect 8009 13068 8055 13120
rect 8055 13068 8058 13120
rect 8487 14588 8489 14640
rect 8489 14588 8535 14640
rect 8535 14588 8539 14640
rect 8326 13068 8329 13120
rect 8329 13068 8375 13120
rect 8375 13068 8378 13120
<< metal2 >>
rect 2520 14640 2916 14652
rect 2520 14588 2532 14640
rect 2584 14588 2852 14640
rect 2904 14588 2916 14640
rect 2520 14584 2916 14588
rect 2972 14640 4328 14652
rect 2972 14588 2984 14640
rect 3036 14588 3304 14640
rect 3356 14588 3624 14640
rect 3676 14588 3944 14640
rect 3996 14588 4264 14640
rect 4316 14588 4328 14640
rect 2972 14584 4328 14588
rect 4390 14640 5746 14652
rect 4390 14588 4402 14640
rect 4454 14588 4722 14640
rect 4774 14588 5042 14640
rect 5094 14588 5362 14640
rect 5414 14588 5682 14640
rect 5734 14588 5746 14640
rect 4390 14584 5746 14588
rect 5914 14640 8551 14652
rect 5914 14588 5926 14640
rect 5978 14588 6246 14640
rect 6298 14588 6566 14640
rect 6618 14588 6886 14640
rect 6938 14588 7206 14640
rect 7258 14588 7526 14640
rect 7578 14588 7846 14640
rect 7898 14588 8166 14640
rect 8218 14588 8487 14640
rect 8539 14588 8551 14640
rect 5914 14584 8551 14588
rect 2680 13120 8390 13124
rect 2680 13068 2692 13120
rect 2744 13068 3144 13120
rect 3196 13068 3464 13120
rect 3516 13068 3784 13120
rect 3836 13068 4104 13120
rect 4156 13068 4562 13120
rect 4614 13068 4882 13120
rect 4934 13068 5202 13120
rect 5254 13068 5522 13120
rect 5574 13068 6086 13120
rect 6138 13068 6406 13120
rect 6458 13068 6726 13120
rect 6778 13068 7046 13120
rect 7098 13068 7366 13120
rect 7418 13068 7686 13120
rect 7738 13068 8006 13120
rect 8058 13068 8326 13120
rect 8378 13068 8390 13120
rect 2680 13056 8390 13068
<< labels >>
flabel metal1 2502 12824 8607 13000 1 FreeSans 800 0 0 0 VSS
port 11 n
flabel metal2 2680 13056 8390 13124 1 FreeSans 800 0 0 0 Cbtm
port 7 n
flabel polysilicon 4480 14698 5656 14734 1 FreeSans 320 180 0 0 EN_VSS
port 9 n
flabel metal2 4390 14584 5746 14652 1 FreeSans 320 180 0 0 VREF_GND
port 2 n
flabel polysilicon 3062 14698 4238 14734 1 FreeSans 320 180 0 0 EN_VCM
port 5 n
flabel metal2 2972 14584 4328 14652 1 FreeSans 320 180 0 0 VCM
port 1 n
flabel polysilicon 2610 14698 2826 14734 1 FreeSans 320 0 0 0 EN_VIN
port 10 n
flabel metal2 2520 14584 2916 14652 5 FreeSans 320 0 0 0 VIN
port 3 s
flabel metal1 2570 14756 8590 14932 1 FreeSans 800 0 0 0 VDD
port 8 n
flabel metal2 5920 14590 8550 14650 0 FreeSans 320 0 0 0 VREF
port 4 nsew
flabel polysilicon 6004 14698 8460 14734 0 FreeSans 320 0 0 0 EN_VREF_Z
port 6 nsew
<< end >>
