magic
tech gf180mcuD
magscale 1 10
timestamp 1757658519
<< nwell >>
rect 4090 4760 4206 5213
rect 2391 4749 2502 4757
rect 3897 4749 4206 4760
rect 2101 4738 4206 4749
rect 2100 4704 4206 4738
rect 2100 4690 4119 4704
rect 2101 4680 4119 4690
rect 2101 4679 4047 4680
rect 2391 4656 2502 4679
rect 3920 4658 4047 4679
rect 5670 4653 7687 4734
rect 1998 2874 2114 2875
rect 1998 2808 2115 2874
rect 5670 2828 9682 2858
rect 9759 2828 9767 3316
rect 5584 2811 9767 2828
rect 1999 2807 2115 2808
rect 5670 2776 9682 2811
rect 9759 2807 9767 2811
rect 7559 2767 7677 2776
rect 213 2324 221 2332
rect 2000 992 2114 993
rect 1998 991 2114 992
rect 1998 921 2115 991
rect 4118 810 4119 1016
rect 7559 960 7677 1030
rect 5584 948 9767 960
rect 5671 920 9681 948
rect 7559 911 7677 920
<< pwell >>
rect 17 4103 74 4182
rect 1989 3805 2120 3807
rect 108 3784 4119 3805
rect 7550 3784 7682 3796
rect 22 3760 4204 3784
rect 5669 3762 9681 3784
rect 5584 3758 9681 3762
rect 5669 3727 9681 3758
rect 7550 3716 7682 3727
rect 65 3610 70 3678
rect 4256 3350 5531 3365
rect 4243 3304 5544 3350
rect 4256 3290 5531 3304
rect 1989 1937 1991 1963
rect 1989 1905 2120 1937
rect 22 1881 4204 1905
rect 7550 1897 7682 1925
rect 9680 1897 9681 1919
rect 5670 1882 9681 1897
rect 108 1873 4119 1881
rect 5584 1878 9681 1882
rect 1989 1861 2120 1873
rect 5670 1847 9681 1878
rect 7550 1834 7682 1847
rect 4256 1686 5531 1705
rect 4243 1640 5544 1686
rect 4256 1630 5531 1640
<< psubdiff >>
rect 3994 5594 4315 5628
rect 3994 5518 4062 5594
rect 4163 5518 4315 5594
rect 3994 5502 4315 5518
rect 5470 5575 5661 5595
rect 5470 5492 5503 5575
rect 5639 5492 5661 5575
rect 5470 5478 5661 5492
rect 1989 3760 2120 3807
rect 7550 3716 7682 3796
rect 4256 3350 5531 3365
rect 4243 3304 5544 3350
rect 4256 3290 5531 3304
rect 1989 1937 1991 1963
rect 1989 1861 2120 1937
rect 7550 1834 7682 1925
rect 4256 1686 5531 1705
rect 4243 1640 5544 1686
rect 4256 1630 5531 1640
<< nsubdiff >>
rect 2391 4741 2502 4757
rect 2391 4671 2407 4741
rect 2488 4671 2502 4741
rect 2391 4656 2502 4671
rect 1998 2874 2114 2875
rect 1998 2808 2115 2874
rect 1999 2807 2115 2808
rect 7559 2767 7677 2855
rect 2000 992 2114 993
rect 1998 991 2114 992
rect 1998 921 2115 991
rect 7559 911 7677 1030
<< psubdiffcont >>
rect 4062 5518 4163 5594
rect 5503 5492 5639 5575
<< nsubdiffcont >>
rect 2407 4671 2488 4741
<< metal1 >>
rect 250 6084 320 6099
rect 250 5997 262 6084
rect 317 5997 320 6084
rect 250 5990 320 5997
rect 251 5323 320 5990
rect 3986 5594 4317 5630
rect 3986 5518 4062 5594
rect 4163 5518 4317 5594
rect 3986 5501 4317 5518
rect 1490 5323 2474 5324
rect 251 5254 2474 5323
rect 2833 5199 2932 5213
rect 2833 5142 2845 5199
rect 2919 5142 2932 5199
rect 2833 5136 2932 5142
rect 4257 4932 4317 5501
rect 5470 5595 5530 5596
rect 5470 5575 5712 5595
rect 5470 5492 5503 5575
rect 5639 5492 5712 5575
rect 5470 5475 5712 5492
rect 5470 4910 5530 5475
rect 6420 5081 6525 5097
rect 6420 5010 6439 5081
rect 6509 5010 6525 5081
rect 10626 5069 10701 5085
rect 7539 5062 8741 5063
rect 10626 5062 10639 5069
rect 6420 5000 6525 5010
rect 7539 4999 10639 5062
rect 10626 4996 10639 4999
rect 10693 4996 10701 5069
rect 10626 4982 10701 4996
rect 2391 4749 2502 4757
rect 3897 4749 4119 4760
rect 2101 4741 4119 4749
rect 2101 4738 2407 4741
rect 2100 4690 2407 4738
rect 2101 4679 2407 4690
rect 2391 4671 2407 4679
rect 2488 4733 4119 4741
rect 2488 4679 3920 4733
rect 2488 4671 2502 4679
rect 2391 4656 2502 4671
rect 4047 4680 4119 4733
rect 5670 4720 7687 4734
rect 5670 4653 5730 4720
rect 5880 4653 7687 4720
rect 10763 4477 10854 4494
rect 10763 4397 10775 4477
rect 10840 4397 10854 4477
rect 10763 4390 10854 4397
rect 9666 4221 9773 4246
rect 9666 4144 9691 4221
rect 9759 4199 9773 4221
rect 10628 4199 10697 4210
rect 9759 4194 10697 4199
rect 9759 4144 10642 4194
rect 9666 4127 10642 4144
rect 9709 4126 10642 4127
rect 10628 4121 10642 4126
rect 10694 4121 10697 4194
rect 10628 4108 10697 4121
rect -709 3996 -630 4000
rect -711 3980 -630 3996
rect -711 3891 -697 3980
rect -641 3891 -630 3980
rect -711 2485 -630 3891
rect 1989 3805 2120 3807
rect 4084 3805 4275 3907
rect 108 3760 4275 3805
rect 4117 3640 4275 3760
rect 4214 3638 4275 3640
rect 5505 3876 5584 3905
rect 5505 3784 5687 3876
rect 7550 3784 7682 3796
rect 5505 3727 9681 3784
rect 5505 3639 5687 3727
rect 7550 3716 7682 3727
rect 5505 3638 5584 3639
rect 4256 3290 5531 3365
rect 9877 3360 9948 3372
rect 9877 3255 9885 3360
rect 9942 3255 9948 3360
rect 9877 3241 9948 3255
rect 1998 2874 2114 2875
rect 1998 2873 2115 2874
rect 108 2864 4119 2873
rect 108 2801 3718 2864
rect 3824 2801 4119 2864
rect 108 2799 4119 2801
rect 5670 2849 9682 2858
rect 5670 2790 5970 2849
rect 6108 2790 9682 2849
rect 5670 2776 9682 2790
rect 7559 2767 7677 2776
rect -711 2404 -694 2485
rect -640 2404 -630 2485
rect -711 2386 -630 2404
rect -220 2135 -140 2150
rect -220 2130 -206 2135
rect -1050 2090 -206 2130
rect -1050 1991 -1027 2090
rect -975 2057 -206 2090
rect -152 2057 -140 2135
rect -975 2040 -140 2057
rect -975 2039 -207 2040
rect -975 1991 -949 2039
rect 4214 2026 4272 2027
rect -1050 1969 -949 1991
rect 108 1873 4272 2026
rect -212 1842 -137 1867
rect 1989 1861 2120 1873
rect -1210 1836 -1130 1837
rect -212 1836 -202 1842
rect -1210 1764 -202 1836
rect -149 1764 -137 1842
rect -1210 1755 -137 1764
rect 4081 1758 4272 1873
rect 5516 1997 5584 2026
rect 5516 1897 5694 1997
rect 7550 1897 7682 1925
rect 9680 1897 9681 1919
rect 5516 1847 9681 1897
rect 5516 1760 5694 1847
rect 7550 1834 7682 1847
rect 5516 1759 5583 1760
rect -1210 1754 -151 1755
rect -1210 1402 -1130 1754
rect 4256 1630 5531 1705
rect -1210 1326 -1198 1402
rect -1137 1326 -1130 1402
rect -1210 1310 -1130 1326
rect 2000 992 2114 993
rect 1998 991 2114 992
rect 1998 985 2115 991
rect 108 919 3716 985
rect 4118 985 4119 1016
rect 3830 919 4119 985
rect 5670 948 6012 960
rect 5671 920 6012 948
rect 4118 810 4119 919
rect 7559 960 7677 1030
rect 6190 920 9681 960
rect 7559 911 7677 920
rect -1211 643 -1130 660
rect -1211 571 -1199 643
rect -1139 571 -1130 643
rect -1211 553 -1130 571
rect -1051 643 -966 660
rect -1051 567 -1040 643
rect -978 567 -966 643
rect -1209 131 -1131 553
rect -1051 287 -966 567
rect -878 646 -794 663
rect -878 570 -867 646
rect -805 570 -794 646
rect -878 290 -794 570
rect -708 648 -624 665
rect -708 572 -697 648
rect -635 572 -624 648
rect -708 292 -624 572
rect -1210 48 -1130 131
rect -1210 -24 -1198 48
rect -1144 -24 -1130 48
rect -1210 -39 -1130 -24
rect -1052 47 -965 287
rect -1052 -23 -1037 47
rect -984 -23 -965 47
rect -1052 -40 -965 -23
rect -879 50 -794 290
rect -879 -20 -864 50
rect -811 -20 -794 50
rect -879 -37 -794 -20
rect -709 52 -624 292
rect -709 -18 -694 52
rect -641 -18 -624 52
rect 4102 27 4272 146
rect 5521 140 5576 146
rect 5521 26 5682 140
rect 5564 19 5682 26
rect 9878 65 9947 3241
rect 10000 2565 10070 2579
rect 10000 2506 10006 2565
rect 10063 2506 10070 2565
rect 10000 342 10070 2506
rect 10141 2564 10212 2581
rect 10141 2562 10213 2564
rect 10141 2498 10154 2562
rect 10000 306 10011 342
rect 9999 267 10011 306
rect 10063 267 10070 342
rect 9999 250 10070 267
rect 10139 2476 10154 2498
rect 10211 2476 10213 2562
rect 10139 2474 10213 2476
rect 10139 2445 10212 2474
rect 10139 351 10209 2445
rect 10764 1680 10854 4390
rect 11589 1680 11705 1681
rect 10764 1579 11705 1680
rect 11193 1451 11302 1469
rect 11193 1350 11216 1451
rect 11293 1350 11302 1451
rect 11193 1339 11302 1350
rect 10900 1196 11102 1207
rect 10900 1130 10918 1196
rect 11028 1130 11102 1196
rect 10900 1116 11102 1130
rect 10759 1027 10914 1042
rect 10759 967 10777 1027
rect 10866 967 10914 1027
rect 10759 955 10914 967
rect 10628 864 10736 874
rect 10628 809 10645 864
rect 10724 809 10736 864
rect 10628 800 10736 809
rect 10630 709 10721 800
rect 10822 758 10914 955
rect 10822 717 10916 758
rect 10139 259 10210 351
rect 10139 190 10209 259
rect 10139 110 10149 190
rect 10202 110 10209 190
rect 10139 91 10209 110
rect -709 -35 -624 -18
rect 9878 -8 9884 65
rect 9941 -8 9947 65
rect 9878 -21 9947 -8
rect 2280 -112 2411 -111
rect 10630 -112 10720 709
rect 2279 -118 10722 -112
rect 2279 -202 2295 -118
rect 2397 -202 10722 -118
rect 2279 -210 10722 -202
rect 10630 -211 10720 -210
rect 10823 -304 10916 717
rect 10576 -305 10916 -304
rect 7326 -306 10916 -305
rect 2280 -316 10916 -306
rect 2280 -392 2299 -316
rect 2391 -392 10916 -316
rect 2280 -397 10916 -392
rect 11009 -499 11102 1116
rect 11195 1108 11300 1339
rect 2277 -509 11102 -499
rect 2277 -591 2289 -509
rect 2397 -552 11102 -509
rect 2397 -591 11100 -552
rect 2277 -596 11100 -591
rect 10862 -597 11100 -596
rect 11194 -691 11300 1108
rect 11411 501 11523 508
rect 10945 -693 11300 -691
rect 2284 -703 11300 -693
rect 2284 -781 2301 -703
rect 2399 -781 11300 -703
rect 11410 486 11523 501
rect 11410 372 11430 486
rect 11507 372 11523 486
rect 11410 359 11523 372
rect 11410 -693 11519 359
rect 11410 -719 11520 -693
rect 2284 -789 11300 -781
rect 7624 -791 11300 -789
rect 11411 -890 11520 -719
rect 2295 -893 11520 -890
rect 2295 -907 11522 -893
rect 2295 -989 2316 -907
rect 2414 -989 11522 -907
rect 2295 -1001 11522 -989
rect 2305 -1070 10245 -1069
rect 11589 -1070 11705 1579
rect 2305 -1077 11705 -1070
rect 2305 -1130 2324 -1077
rect 2421 -1130 11705 -1077
rect 2305 -1141 11705 -1130
rect 6717 -1142 11705 -1141
<< via1 >>
rect 262 5997 317 6084
rect 2845 5142 2919 5199
rect 3590 5115 3676 5182
rect 6076 5113 6162 5173
rect 6439 5010 6509 5081
rect 7292 5002 7375 5056
rect 10639 4996 10693 5069
rect 3920 4586 4047 4733
rect 5730 4620 5880 4720
rect 10775 4397 10840 4477
rect 9691 4144 9759 4221
rect 10642 4121 10694 4194
rect -697 3891 -641 3980
rect 9885 3255 9942 3360
rect 3718 2801 3824 2864
rect 5970 2790 6108 2849
rect -694 2404 -640 2485
rect -1027 1991 -975 2090
rect -206 2057 -152 2135
rect -202 1764 -149 1842
rect -1198 1326 -1137 1402
rect 3716 912 3830 1010
rect 6012 914 6190 999
rect -1199 571 -1139 643
rect -1040 567 -978 643
rect -867 570 -805 646
rect -697 572 -635 648
rect 4875 510 4991 649
rect -1198 -24 -1144 48
rect -1037 -23 -984 47
rect -864 -20 -811 50
rect -694 -18 -641 52
rect 10006 2506 10063 2565
rect 10011 267 10063 342
rect 10154 2476 10211 2562
rect 11216 1350 11293 1451
rect 10918 1130 11028 1196
rect 10777 967 10866 1027
rect 10645 809 10724 864
rect 10149 110 10202 190
rect 9884 -8 9941 65
rect 2295 -202 2397 -118
rect 2299 -392 2391 -316
rect 2289 -591 2397 -509
rect 2301 -781 2399 -703
rect 11430 372 11507 486
rect 2316 -989 2414 -907
rect 2324 -1130 2421 -1077
<< metal2 >>
rect 9951 6261 10013 6262
rect 1429 6258 2394 6261
rect 8165 6259 8423 6260
rect 3220 6258 8423 6259
rect -1386 5906 -1303 6248
rect -1385 399 -1303 5906
rect -1213 5909 -1130 6250
rect -1051 5909 -968 6250
rect -1213 5200 -1129 5909
rect -1051 5908 -966 5909
rect -1212 1595 -1129 5200
rect -1050 4720 -966 5908
rect -881 5908 -798 6250
rect -1049 2306 -967 4720
rect -881 3475 -799 5908
rect -712 4207 -629 6250
rect -551 5868 -464 6249
rect -388 6081 -299 6247
rect -389 6003 -299 6081
rect -241 6075 -151 6249
rect -80 6076 10 6248
rect -241 6069 -150 6075
rect -240 6008 -150 6069
rect -388 5871 -299 6003
rect -241 5997 -150 6008
rect -81 6069 10 6076
rect 88 6069 179 6249
rect -81 6008 9 6069
rect 89 6008 179 6069
rect -81 5998 10 6008
rect -551 5544 -466 5868
rect -551 5451 -540 5544
rect -476 5451 -466 5544
rect -551 5439 -466 5451
rect -387 5532 -302 5871
rect -241 5868 -151 5997
rect -387 5451 -377 5532
rect -314 5451 -302 5532
rect -240 5554 -153 5868
rect -80 5752 10 5998
rect 88 5945 179 6008
rect 250 6084 329 6250
rect 250 5997 262 6084
rect 317 5997 329 6084
rect 250 5983 329 5997
rect 1429 6180 8423 6258
rect 88 5874 95 5945
rect 169 5874 179 5945
rect 88 5862 179 5874
rect -80 5669 -73 5752
rect -2 5669 10 5752
rect -80 5660 10 5669
rect -240 5481 -227 5554
rect -165 5481 -153 5554
rect -240 5470 -153 5481
rect -387 5439 -302 5451
rect 1429 5345 1510 6180
rect 1955 6178 8423 6180
rect 1955 6177 8166 6178
rect -550 5264 1510 5345
rect 1567 6096 7969 6097
rect 1567 6033 8275 6096
rect -711 4185 -630 4207
rect -711 4100 -698 4185
rect -637 4100 -630 4185
rect -711 4089 -630 4100
rect -709 3980 -630 4000
rect -709 3891 -697 3980
rect -641 3891 -630 3980
rect -709 3879 -630 3891
rect -881 3400 -868 3475
rect -812 3400 -799 3475
rect -881 3388 -799 3400
rect -740 3670 -659 3681
rect -740 3600 -729 3670
rect -666 3600 -659 3670
rect -740 3321 -659 3600
rect -880 3240 -659 3321
rect -1049 2230 -1036 2306
rect -975 2230 -967 2306
rect -1049 2214 -967 2230
rect -1050 2123 -967 2130
rect -1212 1525 -1199 1595
rect -1138 1525 -1129 1595
rect -1212 1508 -1129 1525
rect -1051 2090 -967 2123
rect -1051 1991 -1027 2090
rect -975 1991 -967 2090
rect -1210 1402 -1129 1411
rect -1210 1326 -1198 1402
rect -1137 1326 -1129 1402
rect -1210 1314 -1129 1326
rect -1211 1310 -1129 1314
rect -1211 643 -1130 1310
rect -1211 571 -1199 643
rect -1139 571 -1130 643
rect -1211 554 -1130 571
rect -1051 660 -967 1991
rect -879 664 -800 3240
rect -740 3239 -659 3240
rect -711 2485 -630 2500
rect -711 2404 -694 2485
rect -640 2404 -630 2485
rect -711 2386 -630 2404
rect -710 665 -630 2386
rect -550 781 -469 5264
rect 1567 5184 1630 6033
rect 3105 6032 8275 6033
rect 1955 5968 2227 5969
rect -404 5121 1630 5184
rect 1687 5967 2671 5968
rect 3219 5967 8129 5968
rect 1687 5895 8129 5967
rect 8202 5900 8275 6032
rect 1687 5894 2671 5895
rect 1687 5893 1761 5894
rect -404 5120 1532 5121
rect -404 1204 -340 5120
rect 1687 5056 1760 5893
rect 7919 5824 7981 5825
rect 1818 5822 1963 5823
rect 3220 5822 7981 5824
rect 1818 5821 7981 5822
rect -274 4983 1760 5056
rect 1816 5764 7981 5821
rect 1816 5763 7799 5764
rect 1816 5762 3224 5763
rect 1816 5760 1963 5762
rect -274 3133 -201 4983
rect 1816 4909 1876 5760
rect -130 4849 1876 4909
rect 1936 5642 7861 5703
rect 1936 5641 3224 5642
rect -130 3909 -66 4849
rect 1936 4790 2000 5641
rect 2841 5461 4030 5462
rect 2841 5460 4875 5461
rect 2831 5459 4875 5460
rect 6525 5459 7343 5461
rect 2831 5458 7343 5459
rect 2831 5382 7389 5458
rect 2831 5379 6690 5382
rect 2831 5376 4030 5379
rect 2831 5199 2943 5376
rect 7274 5357 7389 5382
rect 2831 5142 2845 5199
rect 2919 5142 2943 5199
rect 6087 5303 6532 5304
rect 6087 5287 6840 5303
rect 6087 5238 6733 5287
rect 2831 5135 2943 5142
rect 3578 5190 4591 5191
rect 6087 5190 6176 5238
rect 6721 5207 6733 5238
rect 6822 5207 6840 5287
rect 6721 5190 6840 5207
rect 3578 5182 6176 5190
rect 3578 5115 3590 5182
rect 3676 5173 6176 5182
rect 3676 5115 6076 5173
rect 3578 5113 6076 5115
rect 6162 5113 6176 5173
rect 3578 5109 6176 5113
rect 4514 5108 6078 5109
rect 6420 5081 6525 5097
rect -10 4728 2000 4790
rect 3897 4733 4119 4760
rect -10 4461 50 4728
rect 1528 4727 1998 4728
rect 3897 4690 3920 4733
rect 3896 4586 3920 4690
rect 4047 4690 4119 4733
rect 4517 4693 4629 5022
rect 6420 5010 6439 5081
rect 6509 5010 6525 5081
rect 7274 5067 7392 5357
rect 6420 5000 6525 5010
rect 7272 5056 7397 5067
rect 7272 5002 7292 5056
rect 7375 5002 7397 5056
rect 6420 4921 6524 5000
rect 7272 4986 7397 5002
rect 6420 4920 7635 4921
rect 6420 4902 7711 4920
rect 6420 4835 7619 4902
rect 7686 4835 7711 4902
rect 6420 4820 7711 4835
rect 7800 4811 7861 5642
rect 7920 4930 7981 5764
rect 8055 5062 8129 5895
rect 8203 5191 8275 5900
rect 8349 5864 8423 6178
rect 8350 5323 8423 5864
rect 9317 5323 9390 6260
rect 8350 5250 9390 5323
rect 8203 5190 8352 5191
rect 9447 5190 9520 6257
rect 8203 5118 9520 5190
rect 9580 5062 9650 6258
rect 8055 4990 9650 5062
rect 8055 4989 9649 4990
rect 9709 4930 9770 6259
rect 7920 4869 9770 4930
rect 7800 4810 8753 4811
rect 9830 4810 9890 6260
rect 7800 4750 9890 4810
rect 9947 5080 10013 6261
rect 10088 5467 10156 6261
rect 10089 5080 10156 5467
rect 10224 5467 10292 6261
rect 10359 5770 10432 6261
rect 10359 5467 10431 5770
rect 10224 5080 10291 5467
rect 10360 5080 10430 5467
rect 10492 5080 10558 6260
rect 10626 5329 10702 6260
rect 10625 5289 10702 5329
rect 10625 5198 10634 5289
rect 10693 5198 10702 5289
rect 10625 5191 10702 5198
rect 10626 5189 10702 5191
rect 5710 4720 5900 4730
rect 5710 4700 5730 4720
rect 5580 4693 5730 4700
rect 4517 4690 5730 4693
rect 4047 4620 5730 4690
rect 5880 4620 5900 4720
rect 9947 4691 10014 5080
rect 10089 5078 10157 5080
rect 10224 5078 10292 5080
rect 10360 5078 10431 5080
rect 10492 5078 10559 5080
rect 7395 4623 10014 4691
rect 4047 4600 5900 4620
rect 4047 4598 5584 4600
rect 4047 4586 4630 4598
rect 3896 4570 4630 4586
rect 3901 4569 4630 4570
rect 0 4182 92 4211
rect 721 4206 853 4363
rect 0 4103 17 4182
rect 74 4103 92 4182
rect 0 4089 92 4103
rect 1287 4130 1370 4131
rect 3242 4130 3959 4131
rect 1287 4129 3959 4130
rect 1287 4128 4064 4129
rect 4141 4128 4209 4255
rect 1287 4059 4209 4128
rect 1287 4020 1370 4059
rect -1 4000 1370 4020
rect -274 2662 -200 3133
rect -130 3084 -60 3909
rect -1 3903 14 4000
rect 80 3940 1370 4000
rect 80 3939 877 3940
rect 80 3903 91 3939
rect -1 3880 91 3903
rect 1 3705 74 3708
rect 0 3678 74 3705
rect 0 3610 14 3678
rect 70 3672 74 3678
rect 70 3610 4211 3672
rect 0 3590 4211 3610
rect 1 3589 4211 3590
rect 67 3588 4211 3589
rect -1 3492 75 3516
rect -1 3393 9 3492
rect 65 3456 75 3492
rect 65 3393 84 3456
rect -1 3387 84 3393
rect 0 3385 84 3387
rect 4118 3263 4211 3588
rect 3880 3120 3968 3136
rect -130 3065 10 3084
rect 21 3065 22 3083
rect -130 3003 22 3065
rect 3880 3042 3893 3120
rect 3960 3042 3968 3120
rect 3880 3021 3968 3042
rect 3689 2881 3846 2885
rect 4517 2881 4629 4569
rect 7411 4347 7483 4623
rect 9769 4450 9912 4451
rect 9769 4381 9945 4450
rect 9666 4221 9773 4246
rect 5562 4132 5668 4149
rect 5562 4072 5575 4132
rect 5650 4072 5668 4132
rect 9666 4144 9691 4221
rect 9759 4144 9773 4221
rect 9666 4127 9773 4144
rect 5562 4060 5668 4072
rect 9875 3978 9945 4381
rect 9875 3931 9946 3978
rect 9877 3368 9946 3931
rect 9877 3360 9948 3368
rect 9684 3325 9772 3343
rect 9684 3246 9698 3325
rect 9759 3246 9772 3325
rect 9684 3233 9772 3246
rect 9877 3255 9885 3360
rect 9942 3255 9948 3360
rect 9877 3241 9948 3255
rect 3689 2877 4629 2881
rect 7411 2911 7480 3148
rect 9671 3110 9776 3131
rect 9671 3026 9686 3110
rect 9764 3026 9776 3110
rect 9671 3010 9776 3026
rect 7411 2910 9877 2911
rect 10090 2910 10157 5078
rect 5580 2877 6132 2878
rect 3689 2864 6132 2877
rect 3689 2801 3718 2864
rect 3824 2849 6132 2864
rect 3824 2801 5970 2849
rect 3689 2790 5970 2801
rect 6108 2790 6132 2849
rect 7411 2844 10157 2910
rect 9775 2843 10157 2844
rect 3689 2780 6132 2790
rect 10225 2780 10292 5078
rect 10361 2941 10431 5078
rect 3690 2772 6132 2780
rect 3690 2771 4629 2772
rect -274 2581 11 2662
rect 21 2581 22 2661
rect -274 2580 -200 2581
rect 0 2291 79 2325
rect 0 2224 14 2291
rect 70 2224 79 2291
rect 0 2210 79 2224
rect 4124 2151 4210 2354
rect -220 2139 329 2151
rect 496 2139 4210 2151
rect -220 2135 4210 2139
rect -220 2057 -206 2135
rect -152 2081 4210 2135
rect -152 2080 4201 2081
rect -152 2057 -139 2080
rect -220 2040 -139 2057
rect -212 1842 -137 1867
rect -212 1764 -202 1842
rect -149 1817 -137 1842
rect -149 1764 205 1817
rect -212 1755 205 1764
rect 143 1720 205 1755
rect 424 1720 2962 1721
rect 143 1658 4212 1720
rect 3855 1657 4212 1658
rect 1 1596 93 1614
rect 1 1518 16 1596
rect 77 1518 93 1596
rect 1 1505 93 1518
rect 4149 1382 4212 1657
rect 3512 1239 3603 1254
rect -404 1203 -189 1204
rect -404 1123 15 1203
rect 3512 1145 3527 1239
rect 3595 1145 3603 1239
rect 3512 1130 3603 1145
rect 3690 1010 3855 1027
rect 3690 912 3716 1010
rect 3830 1000 3855 1010
rect 4517 1007 4629 2771
rect 7413 2714 10292 2780
rect 7413 2461 7481 2714
rect 9775 2713 10292 2714
rect 10360 2935 10431 2941
rect 10000 2573 10070 2579
rect 9767 2565 10070 2573
rect 9767 2506 10006 2565
rect 10063 2506 10070 2565
rect 9767 2502 10070 2506
rect 10000 2488 10070 2502
rect 10141 2564 10212 2581
rect 10141 2562 10213 2564
rect 10141 2476 10154 2562
rect 10211 2476 10213 2562
rect 10141 2474 10213 2476
rect 10141 2445 10212 2474
rect 9702 2366 9783 2376
rect 9702 2275 9715 2366
rect 9775 2275 9783 2366
rect 9702 2263 9783 2275
rect 6091 1657 6190 1672
rect 6091 1586 6096 1657
rect 6181 1586 6190 1657
rect 6091 1554 6190 1586
rect 6034 1480 6194 1554
rect 9674 1463 9781 1479
rect 9674 1362 9686 1463
rect 9769 1362 9781 1463
rect 9674 1352 9781 1362
rect 7410 1059 7481 1291
rect 9680 1228 9788 1238
rect 9680 1145 9696 1228
rect 9781 1145 9788 1228
rect 9680 1126 9788 1145
rect 10063 1059 10161 1062
rect 10360 1059 10429 2935
rect 7410 1038 10430 1059
rect 4517 1005 5583 1007
rect 4517 1000 6208 1005
rect 3830 999 6208 1000
rect 3830 914 6012 999
rect 6190 914 6208 999
rect 7411 990 10430 1038
rect 3830 912 6208 914
rect 3690 894 6208 912
rect 4517 890 6208 894
rect -550 700 11 781
rect 3319 707 3414 722
rect -1051 643 -966 660
rect -1051 567 -1040 643
rect -978 567 -966 643
rect -1051 552 -966 567
rect -879 646 -794 664
rect -879 570 -867 646
rect -805 570 -794 646
rect -1051 551 -967 552
rect -879 549 -794 570
rect -710 648 -624 665
rect -710 572 -697 648
rect -635 572 -624 648
rect 3319 639 3330 707
rect 3404 639 3414 707
rect 3319 621 3414 639
rect -710 551 -624 572
rect -710 550 -630 551
rect -880 399 -794 402
rect -710 399 -624 404
rect -1385 330 95 399
rect 551 311 3233 312
rect 4149 311 4211 521
rect 550 250 4211 311
rect -880 210 -794 213
rect -710 210 -624 215
rect 550 210 610 250
rect 1396 249 3910 250
rect -1383 150 610 210
rect -1383 -129 -1320 150
rect -1384 -331 -1320 -129
rect -1386 -361 -1320 -331
rect -1210 48 -1129 60
rect -1210 -24 -1198 48
rect -1144 -24 -1129 48
rect -1210 -361 -1129 -24
rect -1053 47 -965 60
rect -1053 -23 -1037 47
rect -984 -23 -965 47
rect -1053 -150 -965 -23
rect -880 50 -794 63
rect -880 -20 -864 50
rect -811 -20 -794 50
rect -880 -114 -794 -20
rect -710 52 -624 65
rect -710 -18 -694 52
rect -641 -18 -624 52
rect 4517 -16 4629 890
rect 7414 880 7480 881
rect 10493 880 10559 5078
rect 10626 5069 10701 5085
rect 10626 4996 10639 5069
rect 10693 4996 10701 5069
rect 10626 4992 10701 4996
rect 10625 4713 10701 4992
rect 10779 4920 10846 4925
rect 10626 4330 10701 4713
rect 10771 4913 10846 4920
rect 10771 4829 10779 4913
rect 10841 4829 10846 4913
rect 10771 4817 10846 4829
rect 10771 4639 10845 4817
rect 10770 4494 10846 4639
rect 10763 4477 10854 4494
rect 10763 4397 10775 4477
rect 10840 4397 10854 4477
rect 10763 4390 10854 4397
rect 10768 4330 10840 4331
rect 10626 4270 10840 4330
rect 7414 814 10559 880
rect 10628 4194 10697 4210
rect 10628 4121 10642 4194
rect 10694 4121 10697 4194
rect 10628 4108 10697 4121
rect 10628 874 10696 4108
rect 10768 3460 10840 4270
rect 10768 3456 10980 3460
rect 10768 3399 10981 3456
rect 10760 3322 10830 3340
rect 10760 3238 10772 3322
rect 10828 3238 10830 3322
rect 10760 1042 10830 3238
rect 10899 3040 10981 3399
rect 10900 2510 10981 3040
rect 10900 2430 11140 2510
rect 10900 2357 10972 2369
rect 10900 2267 10905 2357
rect 10965 2267 10972 2357
rect 10900 2256 10972 2267
rect 10900 1207 10971 2256
rect 11058 2163 11140 2430
rect 11059 1610 11140 2163
rect 11059 1532 11460 1610
rect 11059 1530 11461 1532
rect 11193 1468 11302 1469
rect 11193 1451 11303 1468
rect 11193 1350 11216 1451
rect 11293 1350 11303 1451
rect 11193 1339 11303 1350
rect 11195 1338 11303 1339
rect 10900 1196 11039 1207
rect 10900 1130 10918 1196
rect 11028 1130 11039 1196
rect 10900 1116 11039 1130
rect 10760 1027 10880 1042
rect 10760 967 10777 1027
rect 10866 967 10880 1027
rect 10760 954 10880 967
rect 10628 864 10736 874
rect 4842 649 5021 673
rect 4842 510 4875 649
rect 4991 510 5021 649
rect 7414 577 7480 814
rect 10628 809 10645 864
rect 10724 809 10736 864
rect 10628 800 10736 809
rect 9763 713 10739 714
rect 9763 645 10740 713
rect 10279 525 10377 545
rect 4842 485 5021 510
rect 9672 493 9778 517
rect 9672 374 9683 493
rect 9769 374 9778 493
rect 10279 434 10295 525
rect 10365 492 10377 525
rect 10365 434 10571 492
rect 10279 410 10571 434
rect 10280 409 10571 410
rect 9672 363 9778 374
rect 10210 351 10403 352
rect 10169 350 10403 351
rect 5921 342 6382 349
rect 5921 286 6290 342
rect 6375 286 6382 342
rect 10000 342 10403 350
rect 10000 306 10011 342
rect 5921 279 6382 286
rect 9999 267 10011 306
rect 10063 267 10403 342
rect 9999 259 10403 267
rect 9999 250 10070 259
rect 10140 200 10210 201
rect 10140 190 10250 200
rect 10140 110 10149 190
rect 10202 110 10250 190
rect 10140 91 10250 110
rect 9878 65 9947 80
rect 9878 -8 9884 65
rect 9941 44 9947 65
rect 9941 -8 10100 44
rect -880 -150 -795 -114
rect -1052 -337 -965 -150
rect -879 -337 -795 -150
rect -710 -125 -624 -18
rect 9878 -31 10100 -8
rect 4080 -95 9950 -90
rect -560 -111 2292 -109
rect -560 -118 2411 -111
rect -710 -337 -623 -125
rect -560 -126 2295 -118
rect -561 -202 2295 -126
rect 2397 -202 2411 -118
rect 4080 -151 4094 -95
rect 4162 -151 9950 -95
rect 4080 -159 9950 -151
rect -561 -210 2411 -202
rect -561 -335 -474 -210
rect 3880 -232 4354 -231
rect 3880 -237 9804 -232
rect 3880 -294 3890 -237
rect 3965 -294 9804 -237
rect 3880 -301 9804 -294
rect -416 -305 2275 -304
rect -417 -306 2282 -305
rect -417 -316 2407 -306
rect -1052 -361 -964 -337
rect -1386 -1010 -1321 -361
rect -1207 -1009 -1131 -361
rect -1387 -1208 -1320 -1010
rect -1208 -1207 -1130 -1009
rect -1051 -1010 -964 -361
rect -882 -1010 -795 -337
rect -1051 -1021 -963 -1010
rect -1050 -1209 -963 -1021
rect -882 -1208 -794 -1010
rect -713 -1022 -622 -337
rect -562 -478 -473 -335
rect -712 -1209 -622 -1022
rect -564 -498 -473 -478
rect -417 -392 2299 -316
rect 2391 -392 2407 -316
rect 9582 -374 9655 -373
rect -417 -396 2407 -392
rect -564 -1022 -476 -498
rect -417 -705 -328 -396
rect 2280 -397 2407 -396
rect 3696 -381 9655 -374
rect 3696 -437 3708 -381
rect 3776 -437 9655 -381
rect 3696 -446 9655 -437
rect -420 -760 -328 -705
rect -260 -509 2411 -499
rect -260 -591 2289 -509
rect 2397 -591 2411 -509
rect -260 -596 2411 -591
rect 3512 -521 9384 -520
rect 9445 -521 9521 -520
rect 3512 -529 9521 -521
rect 3512 -587 3522 -529
rect 3595 -587 9521 -529
rect 3512 -593 9521 -587
rect -260 -707 -171 -596
rect 3320 -676 9387 -668
rect -564 -1209 -477 -1022
rect -420 -1210 -330 -760
rect -261 -1010 -171 -707
rect -104 -693 2387 -692
rect -104 -703 2410 -693
rect -104 -781 2301 -703
rect 2399 -781 2410 -703
rect 3320 -733 3332 -676
rect 3404 -733 9387 -676
rect 3320 -741 9387 -733
rect -104 -787 2410 -781
rect -102 -788 2410 -787
rect -261 -1020 -170 -1010
rect -102 -1014 19 -788
rect 2284 -789 2410 -788
rect 9311 -825 9387 -741
rect 81 -907 2429 -890
rect 81 -989 2316 -907
rect 2414 -989 2429 -907
rect 81 -1001 2429 -989
rect -102 -1020 20 -1014
rect 81 -1018 200 -1001
rect -260 -1210 -170 -1020
rect -101 -1211 20 -1020
rect 80 -1210 200 -1018
rect 2305 -1070 2431 -1069
rect 276 -1077 2431 -1070
rect 276 -1130 2324 -1077
rect 2421 -1130 2431 -1077
rect 276 -1140 2431 -1130
rect 276 -1210 395 -1140
rect 2305 -1141 2431 -1140
rect 9310 -1114 9388 -825
rect 9445 -956 9521 -593
rect 9582 -822 9655 -446
rect 9732 -512 9804 -301
rect 9732 -526 9805 -512
rect 9310 -1222 9389 -1114
rect 9446 -1130 9521 -956
rect 9581 -1083 9656 -822
rect 9447 -1219 9521 -1130
rect 9580 -1220 9656 -1083
rect 9733 -823 9805 -526
rect 9878 -823 9950 -159
rect 10025 -167 10100 -31
rect 10026 -823 10100 -167
rect 9733 -1058 9808 -823
rect 9733 -1132 9809 -1058
rect 9734 -1220 9809 -1132
rect 9878 -1221 9953 -823
rect 10026 -1220 10101 -823
rect 10175 -1221 10250 91
rect 10326 110 10403 259
rect 10484 231 10571 409
rect 10654 323 10740 645
rect 11378 640 11461 1530
rect 11378 580 11660 640
rect 11379 570 11660 580
rect 11411 492 11523 508
rect 11411 367 11420 492
rect 11514 367 11523 492
rect 11411 359 11523 367
rect 10481 226 10571 231
rect 10326 -1220 10401 110
rect 10481 -821 10570 226
rect 10480 -1220 10570 -821
rect 10653 -952 10740 323
rect 11589 300 11659 570
rect 10810 298 11659 300
rect 10654 -1220 10740 -952
rect 10809 230 11659 298
rect 10809 -1220 10896 230
rect 11590 229 11659 230
<< via2 >>
rect -540 5451 -476 5544
rect -377 5451 -314 5532
rect 95 5874 169 5945
rect -73 5669 -2 5752
rect -227 5481 -165 5554
rect -698 4100 -637 4185
rect -697 3891 -641 3980
rect -868 3400 -812 3475
rect -729 3600 -666 3670
rect -1036 2230 -975 2306
rect -1199 1525 -1138 1595
rect 6733 5207 6822 5287
rect 7619 4835 7686 4902
rect 10634 5198 10693 5289
rect 4101 4419 4165 4475
rect 17 4103 74 4182
rect 14 3903 80 4000
rect 14 3610 70 3678
rect 9 3393 65 3492
rect 3893 3042 3960 3120
rect 5575 4072 5650 4132
rect 5737 3364 5816 3420
rect 9698 3246 9759 3325
rect 9686 3026 9764 3110
rect 3707 2538 3776 2596
rect 14 2224 70 2291
rect 16 1518 77 1596
rect 3527 1145 3595 1239
rect 10154 2476 10211 2562
rect 9715 2275 9775 2366
rect 5912 2192 5987 2248
rect 6096 1586 6181 1657
rect 9686 1362 9769 1463
rect 9696 1145 9781 1228
rect 3330 639 3404 707
rect 10779 4829 10841 4913
rect 10772 3238 10828 3322
rect 10905 2267 10965 2357
rect 11216 1350 11293 1451
rect 4875 510 4991 649
rect 9683 374 9769 493
rect 10295 434 10365 525
rect 6290 286 6375 342
rect 4094 -151 4162 -95
rect 3890 -294 3965 -237
rect 3708 -437 3776 -381
rect 3522 -587 3595 -529
rect 3332 -733 3404 -676
rect 11420 486 11514 492
rect 11420 372 11430 486
rect 11430 372 11507 486
rect 11507 372 11514 486
rect 11420 367 11514 372
<< metal3 >>
rect 89 5954 1532 5957
rect 89 5952 3965 5954
rect 89 5951 6112 5952
rect 89 5945 6384 5951
rect 89 5874 95 5945
rect 169 5874 6384 5945
rect 89 5860 6384 5874
rect 89 5859 1532 5860
rect 3897 5854 6384 5860
rect 5820 5853 6384 5854
rect -79 5758 1532 5762
rect -79 5757 3964 5758
rect -79 5752 6190 5757
rect -79 5669 -73 5752
rect -2 5700 6190 5752
rect -2 5669 6191 5700
rect -79 5664 6191 5669
rect -79 5663 1532 5664
rect 3897 5659 6191 5664
rect 3897 5658 5987 5659
rect -551 5544 -467 5559
rect -551 5451 -540 5544
rect -476 5451 -467 5544
rect -551 5439 -467 5451
rect -387 5532 -302 5591
rect -387 5451 -377 5532
rect -314 5451 -302 5532
rect -239 5557 1532 5567
rect 3897 5557 5995 5562
rect -239 5554 5995 5557
rect -239 5481 -227 5554
rect -165 5481 5995 5554
rect -239 5473 5995 5481
rect -239 5472 1532 5473
rect 3897 5467 5995 5473
rect -550 5193 -468 5439
rect -387 5377 -302 5451
rect -387 5368 1532 5377
rect 3897 5371 5729 5372
rect 3897 5368 5825 5371
rect -387 5284 5825 5368
rect -387 5283 1532 5284
rect 3897 5278 5825 5284
rect -550 5187 1532 5193
rect 3897 5187 4900 5188
rect -550 5186 5558 5187
rect -550 5104 5651 5186
rect 1523 5103 5651 5104
rect 3897 5099 5651 5103
rect 5562 5077 5651 5099
rect 5730 5077 5824 5278
rect 5899 5077 5994 5467
rect 6092 5077 6191 5659
rect 6284 5077 6383 5853
rect 6721 5301 6840 5303
rect 6721 5289 10702 5301
rect 6721 5287 10634 5289
rect 6721 5207 6733 5287
rect 6822 5207 10634 5287
rect 6721 5198 10634 5207
rect 10693 5198 10702 5289
rect 6721 5190 10702 5198
rect 10624 5189 10702 5190
rect 4842 4518 5021 5020
rect 5562 4695 5652 5077
rect 5730 5075 5825 5077
rect 5899 5075 5995 5077
rect 6092 5075 6192 5077
rect 6284 5075 6384 5077
rect 5731 4866 5825 5075
rect 5731 4699 5824 4866
rect 5900 4699 5995 5075
rect 6093 4908 6192 5075
rect 6093 4699 6191 4908
rect 6285 4699 6384 5075
rect 10779 4920 10846 4925
rect 7593 4913 10846 4920
rect 7593 4902 10779 4913
rect 7593 4835 7619 4902
rect 7686 4835 10779 4902
rect 7593 4829 10779 4835
rect 10841 4829 10846 4913
rect 7593 4820 10846 4829
rect 10771 4817 10846 4820
rect 5730 4695 5824 4699
rect 5899 4695 5995 4699
rect 6092 4695 6191 4699
rect 6284 4695 6384 4699
rect 5562 4680 5651 4695
rect 4080 4475 4170 4490
rect 4080 4419 4101 4475
rect 4165 4419 4170 4475
rect 0 4198 93 4211
rect -621 4197 93 4198
rect -712 4185 93 4197
rect -712 4100 -698 4185
rect -637 4182 93 4185
rect -637 4103 17 4182
rect 74 4103 93 4182
rect -637 4100 93 4103
rect -712 4090 93 4100
rect -712 4089 -166 4090
rect -1 4000 91 4020
rect -709 3980 14 4000
rect -709 3891 -697 3980
rect -641 3903 14 3980
rect 80 3903 91 4000
rect -641 3891 91 3903
rect -709 3880 91 3891
rect -709 3879 43 3880
rect 4080 3760 4170 4419
rect 1 3705 74 3708
rect 0 3681 74 3705
rect -740 3678 74 3681
rect -740 3670 14 3678
rect -740 3600 -729 3670
rect -666 3610 14 3670
rect 70 3610 74 3678
rect -666 3600 74 3610
rect -740 3590 74 3600
rect 1 3589 74 3590
rect -1 3496 75 3516
rect -886 3492 75 3496
rect -886 3475 9 3492
rect -886 3400 -868 3475
rect -812 3400 9 3475
rect -886 3393 9 3400
rect 65 3393 75 3492
rect -886 3388 75 3393
rect -886 3387 22 3388
rect 3880 3120 3968 3137
rect 3880 3042 3893 3120
rect 3960 3042 3968 3120
rect 3698 2596 3787 2604
rect 3698 2538 3707 2596
rect 3776 2538 3787 2596
rect -1050 2321 -478 2322
rect 0 2321 79 2325
rect -1050 2306 79 2321
rect -1050 2230 -1036 2306
rect -975 2291 79 2306
rect -975 2230 14 2291
rect -1050 2224 14 2230
rect 70 2224 79 2291
rect -1050 2213 79 2224
rect -787 2212 79 2213
rect 0 2210 79 2212
rect 3698 1905 3787 2538
rect 3696 1874 3787 1905
rect 3880 1905 3968 3042
rect 4080 1905 4169 3760
rect -1212 1596 93 1614
rect -1212 1595 16 1596
rect -1212 1525 -1199 1595
rect -1138 1525 16 1595
rect -1212 1518 16 1525
rect 77 1518 93 1596
rect -1212 1507 93 1518
rect 1 1505 93 1507
rect 3512 1239 3603 1254
rect 3512 1145 3527 1239
rect 3595 1145 3603 1239
rect 3319 707 3414 722
rect 3319 639 3330 707
rect 3404 639 3414 707
rect 3319 -146 3414 639
rect 3319 -635 3413 -146
rect 3512 -529 3603 1145
rect 3696 -381 3786 1874
rect 3880 -204 3970 1905
rect 4080 -75 4170 1905
rect 4840 649 5021 4518
rect 5563 4149 5651 4680
rect 5562 4132 5668 4149
rect 5562 4072 5575 4132
rect 5650 4072 5668 4132
rect 5562 4060 5668 4072
rect 5730 3420 5823 4695
rect 5730 3364 5737 3420
rect 5816 3364 5823 3420
rect 5730 3355 5823 3364
rect 5899 2248 5994 4695
rect 5899 2192 5912 2248
rect 5987 2192 5994 2248
rect 5899 2181 5994 2192
rect 6092 1657 6190 4695
rect 6092 1586 6096 1657
rect 6181 1586 6190 1657
rect 6092 1574 6190 1586
rect 6284 4494 6383 4695
rect 4840 510 4875 649
rect 4991 510 5021 649
rect 4840 485 5021 510
rect 4840 -17 5019 485
rect 6284 342 6382 4494
rect 9684 3327 9772 3343
rect 10760 3327 10830 3340
rect 9684 3325 10830 3327
rect 9684 3246 9698 3325
rect 9759 3322 10830 3325
rect 9759 3246 10772 3322
rect 9684 3238 10772 3246
rect 10828 3238 10830 3322
rect 9684 3233 10830 3238
rect 10760 3223 10830 3233
rect 9671 3110 10280 3131
rect 9671 3026 9686 3110
rect 9764 3026 10280 3110
rect 9671 3012 10280 3026
rect 9671 3010 9776 3012
rect 10160 2584 10279 3012
rect 10137 2562 10280 2584
rect 10137 2476 10154 2562
rect 10211 2476 10280 2562
rect 10137 2442 10280 2476
rect 9702 2366 9783 2376
rect 9702 2275 9715 2366
rect 9775 2364 9783 2366
rect 10900 2364 10972 2369
rect 9775 2357 10972 2364
rect 9775 2275 10905 2357
rect 9702 2267 10905 2275
rect 10965 2267 10972 2357
rect 9702 2263 10972 2267
rect 9719 2261 10972 2263
rect 10900 2256 10972 2261
rect 9674 1463 9781 1479
rect 9674 1362 9686 1463
rect 9769 1461 9781 1463
rect 11193 1461 11302 1469
rect 9769 1451 11302 1461
rect 9769 1362 11216 1451
rect 9674 1352 11216 1362
rect 9779 1350 11216 1352
rect 11293 1350 11302 1451
rect 11193 1339 11302 1350
rect 11199 1338 11302 1339
rect 9679 1228 10374 1241
rect 9679 1145 9696 1228
rect 9781 1145 10374 1228
rect 9679 1127 10374 1145
rect 10283 757 10373 1127
rect 10283 746 10374 757
rect 10279 567 10377 746
rect 10279 529 10378 567
rect 10280 525 10378 529
rect 9674 493 9780 517
rect 9674 385 9683 493
rect 6284 286 6290 342
rect 6375 286 6382 342
rect 6284 280 6382 286
rect 9671 374 9683 385
rect 9769 374 9780 493
rect 10280 434 10295 525
rect 10365 434 10378 525
rect 10280 409 10378 434
rect 11409 492 11538 515
rect 9671 350 9780 374
rect 11409 367 11420 492
rect 11514 367 11538 492
rect 11409 350 11538 367
rect 9671 255 11538 350
rect 9671 254 11537 255
rect 4079 -95 4170 -75
rect 4079 -151 4094 -95
rect 4162 -151 4170 -95
rect 4079 -160 4170 -151
rect 3880 -237 3971 -204
rect 3880 -294 3890 -237
rect 3965 -294 3971 -237
rect 3880 -301 3971 -294
rect 3696 -437 3708 -381
rect 3776 -437 3786 -381
rect 3696 -446 3786 -437
rect 3512 -587 3522 -529
rect 3595 -587 3603 -529
rect 3512 -593 3603 -587
rect 3320 -676 3412 -635
rect 3320 -733 3332 -676
rect 3404 -733 3412 -676
rect 3320 -741 3412 -733
use and_or  and_or_0
timestamp 1757388344
transform 1 0 112 0 1 90
box -112 -90 4101 866
use and_or  and_or_1
timestamp 1757388344
transform 1 0 112 0 -1 1814
box -112 -90 4101 866
use and_or  and_or_2
timestamp 1757388344
transform 1 0 112 0 1 1970
box -112 -90 4101 866
use and_or  and_or_3
timestamp 1757388344
transform 1 0 112 0 -1 3696
box -112 -90 4101 866
use and_or  and_or_4
timestamp 1757388344
transform 1 0 112 0 1 3850
box -112 -90 4101 866
use and_or  and_or_5
timestamp 1757388344
transform 1 0 5674 0 1 3820
box -112 -90 4101 866
use and_or  and_or_6
timestamp 1757388344
transform 1 0 5674 0 1 1942
box -112 -90 4101 866
use and_or  and_or_7
timestamp 1757388344
transform 1 0 5673 0 -1 3664
box -112 -90 4101 866
use and_or  and_or_8
timestamp 1757388344
transform 1 0 5674 0 -1 1786
box -112 -90 4101 866
use and_or  and_or_9
timestamp 1757388344
transform 1 0 5675 0 1 84
box -112 -90 4101 866
use decap_12  decap_12_0
timestamp 1757415140
transform 1 0 4279 0 1 59
box -60 -60 1288 1612
use decap_12  decap_12_1
timestamp 1757415140
transform 1 0 4279 0 1 1720
box -60 -60 1288 1612
use decap_12  decap_12_2
timestamp 1757415140
transform 1 0 4280 0 1 3380
box -60 -60 1288 1612
use gf180mcu_fd_sc_mcu7t5v0__and2_4  gf180mcu_fd_sc_mcu7t5v0__and2_4_0 ~/conda-gf180mcu-env/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 2100 0 -1 5566
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__or2_4  gf180mcu_fd_sc_mcu7t5v0__or2_4_0 ~/conda-gf180mcu-env/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 5670 0 -1 5535
box -86 -86 2102 870
<< labels >>
flabel metal2 9313 -1218 9382 -1114 0 FreeSans 160 0 0 0 EN_VREF_Z_O[0]
port 46 nsew
flabel metal2 9450 -1213 9519 -1109 0 FreeSans 160 0 0 0 EN_VREF_Z_O[1]
port 45 nsew
flabel metal2 9583 -1215 9652 -1111 0 FreeSans 160 0 0 0 EN_VREF_Z_O[2]
port 44 nsew
flabel metal2 9737 -1216 9806 -1112 0 FreeSans 160 0 0 0 EN_VREF_Z_O[3]
port 43 nsew
flabel metal2 9881 -1215 9950 -1111 0 FreeSans 160 0 0 0 EN_VREF_Z_O[4]
port 42 nsew
flabel metal2 10030 -1216 10099 -1112 0 FreeSans 160 0 0 0 EN_VREF_Z_O[5]
port 41 nsew
flabel metal2 10180 -1216 10249 -1112 0 FreeSans 160 0 0 0 EN_VREF_Z_O[6]
port 40 nsew
flabel metal2 10329 -1216 10398 -1112 0 FreeSans 160 0 0 0 EN_VREF_Z_O[7]
port 39 nsew
flabel metal2 10485 -1216 10564 -1108 0 FreeSans 160 0 0 0 EN_VREF_Z_O[8]
port 38 nsew
flabel metal2 10658 -1214 10737 -1106 0 FreeSans 160 0 0 0 EN_VREF_Z_O[9]
port 37 nsew
flabel metal2 10813 -1216 10892 -1108 0 FreeSans 160 0 0 0 EN_VREF_Z_O[10]
port 36 nsew
flabel metal2 9321 6176 9383 6252 0 FreeSans 160 0 0 0 EN_VSS_O[0]
port 35 nsew
flabel metal2 9454 6177 9516 6253 0 FreeSans 160 0 0 0 EN_VSS_O[1]
port 34 nsew
flabel metal2 9582 6177 9644 6253 0 FreeSans 160 0 0 0 EN_VSS_O[2]
port 33 nsew
flabel metal2 9713 6171 9769 6252 0 FreeSans 160 0 0 0 EN_VSS_O[3]
port 32 nsew
flabel metal2 9832 6176 9888 6257 0 FreeSans 160 0 0 0 EN_VSS_O[4]
port 31 nsew
flabel metal2 9951 6176 10012 6260 0 FreeSans 160 0 0 0 EN_VSS_O[5]
port 30 nsew
flabel metal2 10090 6175 10153 6259 0 FreeSans 160 0 0 0 EN_VSS_O[6]
port 29 nsew
flabel metal2 10226 6174 10289 6258 0 FreeSans 160 0 0 0 EN_VSS_O[7]
port 28 nsew
flabel metal2 10363 6168 10426 6255 0 FreeSans 160 0 0 0 EN_VSS_O[8]
port 27 nsew
flabel metal2 10494 6169 10557 6256 0 FreeSans 160 0 0 0 EN_VSS_O[9]
port 26 nsew
flabel metal2 10628 6160 10701 6256 0 FreeSans 160 0 0 0 EN_VSS_O[10]
port 25 nsew
flabel metal3 4854 6 5011 4993 0 FreeSans 320 0 0 0 VSS
port 24 nsew
flabel metal2 4528 94 4623 5002 0 FreeSans 320 0 0 0 VDD
port 23 nsew
flabel metal2 -1385 -1205 -1322 -1100 0 FreeSans 160 0 0 0 EN_VREF_Z_I[0]
port 22 nsew
flabel metal2 -1206 -1205 -1132 -1101 0 FreeSans 160 0 0 0 EN_VREF_Z_I[1]
port 21 nsew
flabel metal2 -1047 -1205 -965 -1101 0 FreeSans 160 0 0 0 EN_VREF_Z_I[2]
port 20 nsew
flabel metal2 -880 -1206 -796 -1104 0 FreeSans 160 0 0 0 EN_VREF_Z_I[3]
port 19 nsew
flabel metal2 -709 -1206 -625 -1104 0 FreeSans 160 0 0 0 EN_VREF_Z_I[4]
port 18 nsew
flabel metal2 -562 -1207 -478 -1105 0 FreeSans 160 0 0 0 EN_VREF_Z_I[5]
port 17 nsew
flabel metal2 -417 -1207 -333 -1105 0 FreeSans 160 0 0 0 EN_VREF_Z_I[6]
port 16 nsew
flabel metal2 -258 -1208 -171 -1107 0 FreeSans 160 0 0 0 EN_VREF_Z_I[7]
port 15 nsew
flabel metal2 -98 -1209 16 -1078 0 FreeSans 160 0 0 0 EN_VREF_Z_I[8]
port 14 nsew
flabel metal2 81 -1209 199 -1077 0 FreeSans 160 0 0 0 EN_VREF_Z_I[9]
port 13 nsew
flabel metal2 276 -1210 394 -1078 0 FreeSans 160 0 0 0 EN_VREF_Z_I[10]
port 12 nsew
flabel metal2 -1385 6149 -1304 6246 0 FreeSans 160 0 0 0 EN_VSS_I[0]
port 11 nsew
flabel metal2 -1212 6150 -1131 6249 0 FreeSans 160 0 0 0 EN_VSS_I[1]
port 10 nsew
flabel metal2 -1050 6151 -969 6250 0 FreeSans 160 0 0 0 EN_VSS_I[2]
port 9 nsew
flabel metal2 -880 6150 -799 6249 0 FreeSans 160 0 0 0 EN_VSS_I[3]
port 8 nsew
flabel metal2 -712 6149 -629 6249 0 FreeSans 160 0 0 0 EN_VSS_I[4]
port 7 nsew
flabel metal2 -550 6138 -465 6245 0 FreeSans 160 0 0 0 EN_VSS_I[5]
port 6 nsew
flabel metal2 -388 6137 -299 6245 0 FreeSans 160 0 0 0 EN_VSS_I[6]
port 5 nsew
flabel metal2 -240 6136 -152 6249 0 FreeSans 160 0 0 0 EN_VSS_I[7]
port 4 nsew
flabel metal2 -80 6146 10 6248 0 FreeSans 160 0 0 0 EN_VSS_I[8]
port 3 nsew
flabel metal2 89 6147 179 6249 0 FreeSans 160 0 0 0 EN_VSS_I[9]
port 2 nsew
flabel metal2 250 6161 329 6250 0 FreeSans 160 0 0 0 EN_VSS_I[10]
port 1 nsew
<< end >>
