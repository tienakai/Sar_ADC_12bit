magic
tech gf180mcuD
magscale 1 10
timestamp 1757727097
<< nwell >>
rect -778 -1798 778 1798
<< pmos >>
rect -604 68 -544 1668
rect -440 68 -380 1668
rect -276 68 -216 1668
rect -112 68 -52 1668
rect 52 68 112 1668
rect 216 68 276 1668
rect 380 68 440 1668
rect 544 68 604 1668
rect -604 -1668 -544 -68
rect -440 -1668 -380 -68
rect -276 -1668 -216 -68
rect -112 -1668 -52 -68
rect 52 -1668 112 -68
rect 216 -1668 276 -68
rect 380 -1668 440 -68
rect 544 -1668 604 -68
<< pdiff >>
rect -692 1655 -604 1668
rect -692 81 -679 1655
rect -633 81 -604 1655
rect -692 68 -604 81
rect -544 1655 -440 1668
rect -544 81 -515 1655
rect -469 81 -440 1655
rect -544 68 -440 81
rect -380 1655 -276 1668
rect -380 81 -351 1655
rect -305 81 -276 1655
rect -380 68 -276 81
rect -216 1655 -112 1668
rect -216 81 -187 1655
rect -141 81 -112 1655
rect -216 68 -112 81
rect -52 1655 52 1668
rect -52 81 -23 1655
rect 23 81 52 1655
rect -52 68 52 81
rect 112 1655 216 1668
rect 112 81 141 1655
rect 187 81 216 1655
rect 112 68 216 81
rect 276 1655 380 1668
rect 276 81 305 1655
rect 351 81 380 1655
rect 276 68 380 81
rect 440 1655 544 1668
rect 440 81 469 1655
rect 515 81 544 1655
rect 440 68 544 81
rect 604 1655 692 1668
rect 604 81 633 1655
rect 679 81 692 1655
rect 604 68 692 81
rect -692 -81 -604 -68
rect -692 -1655 -679 -81
rect -633 -1655 -604 -81
rect -692 -1668 -604 -1655
rect -544 -81 -440 -68
rect -544 -1655 -515 -81
rect -469 -1655 -440 -81
rect -544 -1668 -440 -1655
rect -380 -81 -276 -68
rect -380 -1655 -351 -81
rect -305 -1655 -276 -81
rect -380 -1668 -276 -1655
rect -216 -81 -112 -68
rect -216 -1655 -187 -81
rect -141 -1655 -112 -81
rect -216 -1668 -112 -1655
rect -52 -81 52 -68
rect -52 -1655 -23 -81
rect 23 -1655 52 -81
rect -52 -1668 52 -1655
rect 112 -81 216 -68
rect 112 -1655 141 -81
rect 187 -1655 216 -81
rect 112 -1668 216 -1655
rect 276 -81 380 -68
rect 276 -1655 305 -81
rect 351 -1655 380 -81
rect 276 -1668 380 -1655
rect 440 -81 544 -68
rect 440 -1655 469 -81
rect 515 -1655 544 -81
rect 440 -1668 544 -1655
rect 604 -81 692 -68
rect 604 -1655 633 -81
rect 679 -1655 692 -81
rect 604 -1668 692 -1655
<< pdiffc >>
rect -679 81 -633 1655
rect -515 81 -469 1655
rect -351 81 -305 1655
rect -187 81 -141 1655
rect -23 81 23 1655
rect 141 81 187 1655
rect 305 81 351 1655
rect 469 81 515 1655
rect 633 81 679 1655
rect -679 -1655 -633 -81
rect -515 -1655 -469 -81
rect -351 -1655 -305 -81
rect -187 -1655 -141 -81
rect -23 -1655 23 -81
rect 141 -1655 187 -81
rect 305 -1655 351 -81
rect 469 -1655 515 -81
rect 633 -1655 679 -81
<< polysilicon >>
rect -604 1668 -544 1712
rect -440 1668 -380 1712
rect -276 1668 -216 1712
rect -112 1668 -52 1712
rect 52 1668 112 1712
rect 216 1668 276 1712
rect 380 1668 440 1712
rect 544 1668 604 1712
rect -604 24 -544 68
rect -440 24 -380 68
rect -276 24 -216 68
rect -112 24 -52 68
rect 52 24 112 68
rect 216 24 276 68
rect 380 24 440 68
rect 544 24 604 68
rect -604 -68 -544 -24
rect -440 -68 -380 -24
rect -276 -68 -216 -24
rect -112 -68 -52 -24
rect 52 -68 112 -24
rect 216 -68 276 -24
rect 380 -68 440 -24
rect 544 -68 604 -24
rect -604 -1712 -544 -1668
rect -440 -1712 -380 -1668
rect -276 -1712 -216 -1668
rect -112 -1712 -52 -1668
rect 52 -1712 112 -1668
rect 216 -1712 276 -1668
rect 380 -1712 440 -1668
rect 544 -1712 604 -1668
<< metal1 >>
rect -679 1655 -633 1666
rect -679 70 -633 81
rect -515 1655 -469 1666
rect -515 70 -469 81
rect -351 1655 -305 1666
rect -351 70 -305 81
rect -187 1655 -141 1666
rect -187 70 -141 81
rect -23 1655 23 1666
rect -23 70 23 81
rect 141 1655 187 1666
rect 141 70 187 81
rect 305 1655 351 1666
rect 305 70 351 81
rect 469 1655 515 1666
rect 469 70 515 81
rect 633 1655 679 1666
rect 633 70 679 81
rect -679 -81 -633 -70
rect -679 -1666 -633 -1655
rect -515 -81 -469 -70
rect -515 -1666 -469 -1655
rect -351 -81 -305 -70
rect -351 -1666 -305 -1655
rect -187 -81 -141 -70
rect -187 -1666 -141 -1655
rect -23 -81 23 -70
rect -23 -1666 23 -1655
rect 141 -81 187 -70
rect 141 -1666 187 -1655
rect 305 -81 351 -70
rect 305 -1666 351 -1655
rect 469 -81 515 -70
rect 469 -1666 515 -1655
rect 633 -81 679 -70
rect 633 -1666 679 -1655
<< properties >>
string gencell pfet_03v3
string library gf180mcu
string parameters w 8 l 0.3 m 2 nf 8 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {pfet_03v3 pfet_06v0}
<< end >>
