magic
tech gf180mcuD
magscale 1 10
timestamp 1757727097
<< nwell >>
rect -450 -3534 450 3534
<< pmos >>
rect -276 1804 -216 3404
rect -112 1804 -52 3404
rect 52 1804 112 3404
rect 216 1804 276 3404
rect -276 68 -216 1668
rect -112 68 -52 1668
rect 52 68 112 1668
rect 216 68 276 1668
rect -276 -1668 -216 -68
rect -112 -1668 -52 -68
rect 52 -1668 112 -68
rect 216 -1668 276 -68
rect -276 -3404 -216 -1804
rect -112 -3404 -52 -1804
rect 52 -3404 112 -1804
rect 216 -3404 276 -1804
<< pdiff >>
rect -364 3391 -276 3404
rect -364 1817 -351 3391
rect -305 1817 -276 3391
rect -364 1804 -276 1817
rect -216 3391 -112 3404
rect -216 1817 -187 3391
rect -141 1817 -112 3391
rect -216 1804 -112 1817
rect -52 3391 52 3404
rect -52 1817 -23 3391
rect 23 1817 52 3391
rect -52 1804 52 1817
rect 112 3391 216 3404
rect 112 1817 141 3391
rect 187 1817 216 3391
rect 112 1804 216 1817
rect 276 3391 364 3404
rect 276 1817 305 3391
rect 351 1817 364 3391
rect 276 1804 364 1817
rect -364 1655 -276 1668
rect -364 81 -351 1655
rect -305 81 -276 1655
rect -364 68 -276 81
rect -216 1655 -112 1668
rect -216 81 -187 1655
rect -141 81 -112 1655
rect -216 68 -112 81
rect -52 1655 52 1668
rect -52 81 -23 1655
rect 23 81 52 1655
rect -52 68 52 81
rect 112 1655 216 1668
rect 112 81 141 1655
rect 187 81 216 1655
rect 112 68 216 81
rect 276 1655 364 1668
rect 276 81 305 1655
rect 351 81 364 1655
rect 276 68 364 81
rect -364 -81 -276 -68
rect -364 -1655 -351 -81
rect -305 -1655 -276 -81
rect -364 -1668 -276 -1655
rect -216 -81 -112 -68
rect -216 -1655 -187 -81
rect -141 -1655 -112 -81
rect -216 -1668 -112 -1655
rect -52 -81 52 -68
rect -52 -1655 -23 -81
rect 23 -1655 52 -81
rect -52 -1668 52 -1655
rect 112 -81 216 -68
rect 112 -1655 141 -81
rect 187 -1655 216 -81
rect 112 -1668 216 -1655
rect 276 -81 364 -68
rect 276 -1655 305 -81
rect 351 -1655 364 -81
rect 276 -1668 364 -1655
rect -364 -1817 -276 -1804
rect -364 -3391 -351 -1817
rect -305 -3391 -276 -1817
rect -364 -3404 -276 -3391
rect -216 -1817 -112 -1804
rect -216 -3391 -187 -1817
rect -141 -3391 -112 -1817
rect -216 -3404 -112 -3391
rect -52 -1817 52 -1804
rect -52 -3391 -23 -1817
rect 23 -3391 52 -1817
rect -52 -3404 52 -3391
rect 112 -1817 216 -1804
rect 112 -3391 141 -1817
rect 187 -3391 216 -1817
rect 112 -3404 216 -3391
rect 276 -1817 364 -1804
rect 276 -3391 305 -1817
rect 351 -3391 364 -1817
rect 276 -3404 364 -3391
<< pdiffc >>
rect -351 1817 -305 3391
rect -187 1817 -141 3391
rect -23 1817 23 3391
rect 141 1817 187 3391
rect 305 1817 351 3391
rect -351 81 -305 1655
rect -187 81 -141 1655
rect -23 81 23 1655
rect 141 81 187 1655
rect 305 81 351 1655
rect -351 -1655 -305 -81
rect -187 -1655 -141 -81
rect -23 -1655 23 -81
rect 141 -1655 187 -81
rect 305 -1655 351 -81
rect -351 -3391 -305 -1817
rect -187 -3391 -141 -1817
rect -23 -3391 23 -1817
rect 141 -3391 187 -1817
rect 305 -3391 351 -1817
<< polysilicon >>
rect -276 3404 -216 3448
rect -112 3404 -52 3448
rect 52 3404 112 3448
rect 216 3404 276 3448
rect -276 1760 -216 1804
rect -112 1760 -52 1804
rect 52 1760 112 1804
rect 216 1760 276 1804
rect -276 1668 -216 1712
rect -112 1668 -52 1712
rect 52 1668 112 1712
rect 216 1668 276 1712
rect -276 24 -216 68
rect -112 24 -52 68
rect 52 24 112 68
rect 216 24 276 68
rect -276 -68 -216 -24
rect -112 -68 -52 -24
rect 52 -68 112 -24
rect 216 -68 276 -24
rect -276 -1712 -216 -1668
rect -112 -1712 -52 -1668
rect 52 -1712 112 -1668
rect 216 -1712 276 -1668
rect -276 -1804 -216 -1760
rect -112 -1804 -52 -1760
rect 52 -1804 112 -1760
rect 216 -1804 276 -1760
rect -276 -3448 -216 -3404
rect -112 -3448 -52 -3404
rect 52 -3448 112 -3404
rect 216 -3448 276 -3404
<< metal1 >>
rect -351 3391 -305 3402
rect -351 1806 -305 1817
rect -187 3391 -141 3402
rect -187 1806 -141 1817
rect -23 3391 23 3402
rect -23 1806 23 1817
rect 141 3391 187 3402
rect 141 1806 187 1817
rect 305 3391 351 3402
rect 305 1806 351 1817
rect -351 1655 -305 1666
rect -351 70 -305 81
rect -187 1655 -141 1666
rect -187 70 -141 81
rect -23 1655 23 1666
rect -23 70 23 81
rect 141 1655 187 1666
rect 141 70 187 81
rect 305 1655 351 1666
rect 305 70 351 81
rect -351 -81 -305 -70
rect -351 -1666 -305 -1655
rect -187 -81 -141 -70
rect -187 -1666 -141 -1655
rect -23 -81 23 -70
rect -23 -1666 23 -1655
rect 141 -81 187 -70
rect 141 -1666 187 -1655
rect 305 -81 351 -70
rect 305 -1666 351 -1655
rect -351 -1817 -305 -1806
rect -351 -3402 -305 -3391
rect -187 -1817 -141 -1806
rect -187 -3402 -141 -3391
rect -23 -1817 23 -1806
rect -23 -3402 23 -3391
rect 141 -1817 187 -1806
rect 141 -3402 187 -3391
rect 305 -1817 351 -1806
rect 305 -3402 351 -3391
<< properties >>
string gencell pfet_03v3
string library gf180mcu
string parameters w 8 l 0.3 m 4 nf 4 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {pfet_03v3 pfet_06v0}
<< end >>
