magic
tech gf180mcuD
magscale 1 10
timestamp 1757727097
<< nwell >>
rect -334 -2650 3601 2164
<< pmos >>
rect 1916 130 1976 1730
rect 2080 130 2140 1730
rect 2244 130 2304 1730
rect 2408 130 2468 1730
rect 2572 130 2632 1730
rect 2736 130 2796 1730
rect 2900 130 2960 1730
rect 3064 130 3124 1730
rect 175 -2123 235 -523
rect 339 -2123 399 -523
rect 503 -2123 563 -523
rect 667 -2123 727 -523
rect 831 -2123 891 -523
rect 995 -2123 1055 -523
rect 1159 -2123 1219 -523
rect 1323 -2123 1383 -523
rect 1917 -2123 1977 -523
rect 2081 -2123 2141 -523
rect 2245 -2123 2305 -523
rect 2409 -2123 2469 -523
rect 2573 -2123 2633 -523
rect 2737 -2123 2797 -523
rect 2901 -2123 2961 -523
rect 3065 -2123 3125 -523
<< pdiff >>
rect 95 132 167 1728
rect 263 132 335 1728
rect 427 132 499 1728
rect 591 132 663 1728
rect 754 132 826 1728
rect 919 132 991 1728
rect 1083 132 1155 1728
rect 1246 132 1318 1728
rect 1388 132 1460 1728
rect 1828 1717 1916 1730
rect 1828 143 1841 1717
rect 1887 143 1916 1717
rect 1828 130 1916 143
rect 1976 1717 2080 1730
rect 1976 143 2005 1717
rect 2051 143 2080 1717
rect 1976 130 2080 143
rect 2140 1717 2244 1730
rect 2140 143 2169 1717
rect 2215 143 2244 1717
rect 2140 130 2244 143
rect 2304 1717 2408 1730
rect 2304 143 2333 1717
rect 2379 143 2408 1717
rect 2304 130 2408 143
rect 2468 1717 2572 1730
rect 2468 143 2497 1717
rect 2543 143 2572 1717
rect 2468 130 2572 143
rect 2632 1717 2736 1730
rect 2632 143 2661 1717
rect 2707 143 2736 1717
rect 2632 130 2736 143
rect 2796 1717 2900 1730
rect 2796 143 2825 1717
rect 2871 143 2900 1717
rect 2796 130 2900 143
rect 2960 1717 3064 1730
rect 2960 143 2989 1717
rect 3035 143 3064 1717
rect 2960 130 3064 143
rect 3124 1717 3212 1730
rect 3124 143 3153 1717
rect 3199 143 3212 1717
rect 3124 130 3212 143
rect 87 -536 175 -523
rect 87 -2110 100 -536
rect 146 -2110 175 -536
rect 87 -2123 175 -2110
rect 235 -536 339 -523
rect 235 -2110 264 -536
rect 310 -2110 339 -536
rect 235 -2123 339 -2110
rect 399 -536 503 -523
rect 399 -2110 428 -536
rect 474 -2110 503 -536
rect 399 -2123 503 -2110
rect 563 -536 667 -523
rect 563 -2110 592 -536
rect 638 -2110 667 -536
rect 563 -2123 667 -2110
rect 727 -536 831 -523
rect 727 -2110 756 -536
rect 802 -2110 831 -536
rect 727 -2123 831 -2110
rect 891 -536 995 -523
rect 891 -2110 920 -536
rect 966 -2110 995 -536
rect 891 -2123 995 -2110
rect 1055 -536 1159 -523
rect 1055 -2110 1084 -536
rect 1130 -2110 1159 -536
rect 1055 -2123 1159 -2110
rect 1219 -536 1323 -523
rect 1219 -2110 1248 -536
rect 1294 -2110 1323 -536
rect 1219 -2123 1323 -2110
rect 1383 -536 1471 -523
rect 1383 -2110 1412 -536
rect 1458 -2110 1471 -536
rect 1383 -2123 1471 -2110
rect 1829 -536 1917 -523
rect 1829 -2110 1842 -536
rect 1888 -2110 1917 -536
rect 1829 -2123 1917 -2110
rect 1977 -536 2081 -523
rect 1977 -2110 2006 -536
rect 2052 -2110 2081 -536
rect 1977 -2123 2081 -2110
rect 2141 -536 2245 -523
rect 2141 -2110 2170 -536
rect 2216 -2110 2245 -536
rect 2141 -2123 2245 -2110
rect 2305 -536 2409 -523
rect 2305 -2110 2334 -536
rect 2380 -2110 2409 -536
rect 2305 -2123 2409 -2110
rect 2469 -536 2573 -523
rect 2469 -2110 2498 -536
rect 2544 -2110 2573 -536
rect 2469 -2123 2573 -2110
rect 2633 -536 2737 -523
rect 2633 -2110 2662 -536
rect 2708 -2110 2737 -536
rect 2633 -2123 2737 -2110
rect 2797 -536 2901 -523
rect 2797 -2110 2826 -536
rect 2872 -2110 2901 -536
rect 2797 -2123 2901 -2110
rect 2961 -536 3065 -523
rect 2961 -2110 2990 -536
rect 3036 -2110 3065 -536
rect 2961 -2123 3065 -2110
rect 3125 -536 3213 -523
rect 3125 -2110 3154 -536
rect 3200 -2110 3213 -536
rect 3125 -2123 3213 -2110
<< pdiffc >>
rect 1841 143 1887 1717
rect 2005 143 2051 1717
rect 2169 143 2215 1717
rect 2333 143 2379 1717
rect 2497 143 2543 1717
rect 2661 143 2707 1717
rect 2825 143 2871 1717
rect 2989 143 3035 1717
rect 3153 143 3199 1717
rect 100 -2110 146 -536
rect 264 -2110 310 -536
rect 428 -2110 474 -536
rect 592 -2110 638 -536
rect 756 -2110 802 -536
rect 920 -2110 966 -536
rect 1084 -2110 1130 -536
rect 1248 -2110 1294 -536
rect 1412 -2110 1458 -536
rect 1842 -2110 1888 -536
rect 2006 -2110 2052 -536
rect 2170 -2110 2216 -536
rect 2334 -2110 2380 -536
rect 2498 -2110 2544 -536
rect 2662 -2110 2708 -536
rect 2826 -2110 2872 -536
rect 2990 -2110 3036 -536
rect 3154 -2110 3200 -536
<< nsubdiff >>
rect -174 1991 3381 2059
rect -175 1970 3381 1991
rect -175 1894 -80 1970
rect -174 1859 -82 1894
rect -174 -2271 -159 1859
rect -99 -2271 -82 1859
rect 1550 1813 1640 1970
rect 3292 1899 3381 1970
rect 1550 4 1566 1813
rect 1627 4 1640 1813
rect 3292 1813 3382 1899
rect 1550 -28 1640 4
rect 1550 -60 1642 -28
rect 3292 4 3308 1813
rect 3369 4 3382 1813
rect 3292 -38 3382 4
rect 3292 -60 3384 -38
rect 1551 -360 1642 -60
rect 1551 -440 1641 -360
rect 3293 -370 3384 -60
rect -174 -2294 -82 -2271
rect -174 -2380 -79 -2294
rect 1551 -2249 1567 -440
rect 1628 -2249 1641 -440
rect 3293 -440 3383 -370
rect 1551 -2294 1641 -2249
rect -175 -2382 63 -2380
rect 1548 -2382 1643 -2294
rect 3293 -2249 3309 -440
rect 3370 -2249 3383 -440
rect 3293 -2297 3383 -2249
rect 3289 -2382 3384 -2297
rect -175 -2394 3384 -2382
rect -175 -2471 3380 -2394
<< nsubdiffcont >>
rect -159 -2271 -99 1859
rect 1566 4 1627 1813
rect 3308 4 3369 1813
rect 1567 -2249 1628 -440
rect 3309 -2249 3370 -440
<< polysilicon >>
rect 160 1865 251 1880
rect 160 1816 177 1865
rect 236 1816 251 1865
rect 160 1800 251 1816
rect 485 1864 576 1880
rect 485 1813 500 1864
rect 561 1813 576 1864
rect 485 1800 576 1813
rect 815 1865 906 1879
rect 815 1814 830 1865
rect 891 1814 906 1865
rect 174 1770 235 1800
rect 502 1770 563 1800
rect 815 1799 906 1814
rect 1144 1864 1235 1879
rect 1144 1813 1160 1864
rect 1221 1813 1235 1864
rect 1144 1799 1235 1813
rect 830 1769 890 1799
rect 1158 1769 1218 1799
rect 337 20 398 92
rect 665 20 726 90
rect 994 25 1054 91
rect 993 20 1054 25
rect 1322 24 1382 91
rect 1322 20 1383 24
rect 320 1 412 20
rect 320 -47 335 1
rect 395 -47 412 1
rect 320 -60 412 -47
rect 650 1 742 20
rect 650 -47 666 1
rect 726 -47 742 1
rect 650 -60 742 -47
rect 978 1 1070 20
rect 978 -47 995 1
rect 1055 -47 1070 1
rect 978 -60 1070 -47
rect 1305 3 1397 20
rect 1305 -45 1321 3
rect 1381 -45 1397 3
rect 1305 -60 1397 -45
rect 1902 1865 1993 1880
rect 1902 1816 1919 1865
rect 1978 1816 1993 1865
rect 1902 1800 1993 1816
rect 2227 1864 2318 1880
rect 2227 1813 2242 1864
rect 2303 1813 2318 1864
rect 2227 1800 2318 1813
rect 2557 1865 2648 1879
rect 2557 1814 2572 1865
rect 2633 1814 2648 1865
rect 1916 1770 1977 1800
rect 1916 1730 1976 1770
rect 2080 1730 2140 1774
rect 2244 1770 2305 1800
rect 2557 1799 2648 1814
rect 2886 1864 2977 1879
rect 2886 1813 2902 1864
rect 2963 1813 2977 1864
rect 2886 1799 2977 1813
rect 2244 1730 2304 1770
rect 2408 1730 2468 1774
rect 2572 1730 2632 1799
rect 2736 1730 2796 1774
rect 2900 1730 2960 1799
rect 3064 1730 3124 1774
rect 1916 86 1976 130
rect 2080 92 2140 130
rect 2079 20 2140 92
rect 2244 86 2304 130
rect 2408 90 2468 130
rect 2407 20 2468 90
rect 2572 86 2632 130
rect 2736 25 2796 130
rect 2900 86 2960 130
rect 2735 20 2796 25
rect 3064 24 3124 130
rect 3064 20 3125 24
rect 2062 1 2154 20
rect 2062 -47 2077 1
rect 2137 -47 2154 1
rect 2062 -60 2154 -47
rect 2392 1 2484 20
rect 2392 -47 2408 1
rect 2468 -47 2484 1
rect 2392 -60 2484 -47
rect 2720 1 2812 20
rect 2720 -47 2737 1
rect 2797 -47 2812 1
rect 2720 -60 2812 -47
rect 3047 3 3139 20
rect 3047 -45 3063 3
rect 3123 -45 3139 3
rect 3047 -60 3139 -45
rect 161 -388 252 -373
rect 161 -437 178 -388
rect 237 -437 252 -388
rect 161 -453 252 -437
rect 486 -389 577 -373
rect 486 -440 501 -389
rect 562 -440 577 -389
rect 486 -453 577 -440
rect 816 -388 907 -374
rect 816 -439 831 -388
rect 892 -439 907 -388
rect 175 -483 236 -453
rect 175 -523 235 -483
rect 339 -523 399 -479
rect 503 -483 564 -453
rect 816 -454 907 -439
rect 1145 -389 1236 -374
rect 1145 -440 1161 -389
rect 1222 -440 1236 -389
rect 1145 -454 1236 -440
rect 503 -523 563 -483
rect 667 -523 727 -479
rect 831 -523 891 -454
rect 995 -523 1055 -479
rect 1159 -523 1219 -454
rect 1323 -523 1383 -479
rect 175 -2167 235 -2123
rect 339 -2161 399 -2123
rect 338 -2233 399 -2161
rect 503 -2167 563 -2123
rect 667 -2163 727 -2123
rect 666 -2233 727 -2163
rect 831 -2167 891 -2123
rect 995 -2228 1055 -2123
rect 1159 -2167 1219 -2123
rect 994 -2233 1055 -2228
rect 1323 -2229 1383 -2123
rect 1323 -2233 1384 -2229
rect 321 -2252 413 -2233
rect 321 -2300 336 -2252
rect 396 -2300 413 -2252
rect 321 -2313 413 -2300
rect 651 -2252 743 -2233
rect 651 -2300 667 -2252
rect 727 -2300 743 -2252
rect 651 -2313 743 -2300
rect 979 -2252 1071 -2233
rect 979 -2300 996 -2252
rect 1056 -2300 1071 -2252
rect 979 -2313 1071 -2300
rect 1306 -2250 1398 -2233
rect 1306 -2298 1322 -2250
rect 1382 -2298 1398 -2250
rect 1903 -388 1994 -373
rect 1903 -437 1920 -388
rect 1979 -437 1994 -388
rect 1903 -453 1994 -437
rect 2228 -389 2319 -373
rect 2228 -440 2243 -389
rect 2304 -440 2319 -389
rect 2228 -453 2319 -440
rect 2558 -388 2649 -374
rect 2558 -439 2573 -388
rect 2634 -439 2649 -388
rect 1917 -483 1978 -453
rect 1917 -523 1977 -483
rect 2081 -523 2141 -479
rect 2245 -483 2306 -453
rect 2558 -454 2649 -439
rect 2887 -389 2978 -374
rect 2887 -440 2903 -389
rect 2964 -440 2978 -389
rect 2887 -454 2978 -440
rect 2245 -523 2305 -483
rect 2409 -523 2469 -479
rect 2573 -523 2633 -454
rect 2737 -523 2797 -479
rect 2901 -523 2961 -454
rect 3065 -523 3125 -479
rect 1917 -2167 1977 -2123
rect 2081 -2161 2141 -2123
rect 2080 -2233 2141 -2161
rect 2245 -2167 2305 -2123
rect 2409 -2163 2469 -2123
rect 2408 -2233 2469 -2163
rect 2573 -2167 2633 -2123
rect 2737 -2228 2797 -2123
rect 2901 -2167 2961 -2123
rect 2736 -2233 2797 -2228
rect 3065 -2229 3125 -2123
rect 3065 -2233 3126 -2229
rect 2063 -2252 2155 -2233
rect 1306 -2313 1398 -2298
rect 2063 -2300 2078 -2252
rect 2138 -2300 2155 -2252
rect 2063 -2313 2155 -2300
rect 2393 -2252 2485 -2233
rect 2393 -2300 2409 -2252
rect 2469 -2300 2485 -2252
rect 2393 -2313 2485 -2300
rect 2721 -2252 2813 -2233
rect 2721 -2300 2738 -2252
rect 2798 -2300 2813 -2252
rect 2721 -2313 2813 -2300
rect 3048 -2250 3140 -2233
rect 3048 -2298 3064 -2250
rect 3124 -2298 3140 -2250
rect 3048 -2313 3140 -2298
<< polycontact >>
rect 177 1816 236 1865
rect 500 1813 561 1864
rect 830 1814 891 1865
rect 1160 1813 1221 1864
rect 335 -47 395 1
rect 666 -47 726 1
rect 995 -47 1055 1
rect 1321 -45 1381 3
rect 1919 1816 1978 1865
rect 2242 1813 2303 1864
rect 2572 1814 2633 1865
rect 2902 1813 2963 1864
rect 2077 -47 2137 1
rect 2408 -47 2468 1
rect 2737 -47 2797 1
rect 3063 -45 3123 3
rect 178 -437 237 -388
rect 501 -440 562 -389
rect 831 -439 892 -388
rect 1161 -440 1222 -389
rect 336 -2300 396 -2252
rect 667 -2300 727 -2252
rect 996 -2300 1056 -2252
rect 1322 -2298 1382 -2250
rect 1920 -437 1979 -388
rect 2243 -440 2304 -389
rect 2573 -439 2634 -388
rect 2903 -440 2964 -389
rect 2078 -2300 2138 -2252
rect 2409 -2300 2469 -2252
rect 2738 -2300 2798 -2252
rect 3064 -2298 3124 -2250
<< metal1 >>
rect -174 1991 3381 2059
rect -175 1970 3381 1991
rect -175 1894 -80 1970
rect -174 1859 -82 1894
rect -174 -2271 -159 1859
rect -99 -2271 -82 1859
rect -22 1879 635 1881
rect -22 1865 1235 1879
rect -22 1816 177 1865
rect 236 1864 830 1865
rect 236 1816 500 1864
rect -22 393 45 1816
rect 160 1813 500 1816
rect 561 1814 830 1864
rect 891 1864 1235 1865
rect 891 1814 1160 1864
rect 561 1813 1160 1814
rect 1221 1813 1235 1864
rect 160 1810 1235 1813
rect 160 1800 251 1810
rect 485 1800 576 1810
rect 815 1799 906 1810
rect 1144 1799 1235 1810
rect 1550 1813 1640 1970
rect 3292 1899 3381 1970
rect 95 1713 167 1728
rect -22 8 46 393
rect 95 150 103 1713
rect 155 150 167 1713
rect 95 132 167 150
rect 263 1714 335 1728
rect 263 150 267 1714
rect 319 150 335 1714
rect 263 132 335 150
rect 427 1714 499 1728
rect 427 150 434 1714
rect 486 150 499 1714
rect 427 132 499 150
rect 591 1714 663 1728
rect 591 150 601 1714
rect 653 150 663 1714
rect 591 132 663 150
rect 754 1714 826 1728
rect 754 150 763 1714
rect 815 150 826 1714
rect 754 132 826 150
rect 919 1714 991 1728
rect 919 150 930 1714
rect 982 150 991 1714
rect 919 132 991 150
rect 1083 1714 1155 1728
rect 1083 150 1095 1714
rect 1147 150 1155 1714
rect 1083 132 1155 150
rect 1246 1714 1318 1728
rect 1246 150 1257 1714
rect 1309 150 1318 1714
rect 1246 132 1318 150
rect 1388 1713 1460 1728
rect 1388 149 1398 1713
rect 1450 149 1460 1713
rect 1388 132 1460 149
rect 320 10 412 20
rect 650 10 742 20
rect 978 10 1070 20
rect 1305 10 1397 20
rect 320 8 1397 10
rect -22 1 1320 8
rect 1383 6 1397 8
rect -22 -47 335 1
rect 395 -47 666 1
rect 726 -47 995 1
rect 1055 -47 1320 1
rect -22 -51 1320 -47
rect 1383 -51 1398 6
rect -22 -60 1398 -51
rect 1550 4 1566 1813
rect 1627 4 1640 1813
rect 1550 -28 1640 4
rect 1720 1879 2377 1881
rect 1720 1865 2977 1879
rect 1720 1816 1919 1865
rect 1978 1864 2572 1865
rect 1978 1816 2242 1864
rect 1720 393 1787 1816
rect 1902 1813 2242 1816
rect 2303 1814 2572 1864
rect 2633 1864 2977 1865
rect 2633 1814 2902 1864
rect 2303 1813 2902 1814
rect 2963 1813 2977 1864
rect 1902 1810 2977 1813
rect 1902 1800 1993 1810
rect 2227 1800 2318 1810
rect 2557 1799 2648 1810
rect 2886 1799 2977 1810
rect 3292 1813 3382 1899
rect 1837 1717 1909 1728
rect 1720 8 1788 393
rect 1837 143 1841 1717
rect 1887 1713 1909 1717
rect 1897 150 1909 1713
rect 1887 143 1909 150
rect 1837 132 1909 143
rect 2005 1717 2077 1728
rect 2051 1714 2077 1717
rect 2061 150 2077 1714
rect 2051 143 2077 150
rect 2005 132 2077 143
rect 2169 1717 2241 1728
rect 2215 1714 2241 1717
rect 2228 150 2241 1714
rect 2215 143 2241 150
rect 2169 132 2241 143
rect 2333 1717 2405 1728
rect 2379 1714 2405 1717
rect 2395 150 2405 1714
rect 2379 143 2405 150
rect 2333 132 2405 143
rect 2496 1717 2568 1728
rect 2496 143 2497 1717
rect 2543 1714 2568 1717
rect 2557 150 2568 1714
rect 2543 143 2568 150
rect 2496 132 2568 143
rect 2661 1717 2733 1728
rect 2707 1714 2733 1717
rect 2724 150 2733 1714
rect 2707 143 2733 150
rect 2661 132 2733 143
rect 2825 1717 2897 1728
rect 2871 1714 2897 1717
rect 2889 150 2897 1714
rect 2871 143 2897 150
rect 2825 132 2897 143
rect 2988 1717 3060 1728
rect 2988 143 2989 1717
rect 3035 1714 3060 1717
rect 3051 150 3060 1714
rect 3035 143 3060 150
rect 2988 132 3060 143
rect 3130 1717 3202 1728
rect 3130 1713 3153 1717
rect 3130 149 3140 1713
rect 3130 143 3153 149
rect 3199 143 3202 1717
rect 3130 132 3202 143
rect 2062 10 2154 20
rect 2392 10 2484 20
rect 2720 10 2812 20
rect 3047 10 3139 20
rect 2062 8 3139 10
rect 1720 1 2078 8
rect 2142 6 3139 8
rect 2142 3 3140 6
rect 2142 1 3063 3
rect 1550 -60 1642 -28
rect 1720 -47 2077 1
rect 2142 -47 2408 1
rect 2468 -47 2737 1
rect 2797 -45 3063 1
rect 3123 -45 3140 3
rect 2797 -47 3140 -45
rect 1720 -48 2078 -47
rect 2142 -48 3140 -47
rect 1720 -60 3140 -48
rect 3292 4 3308 1813
rect 3369 4 3382 1813
rect 3292 -38 3382 4
rect 3292 -60 3384 -38
rect 1551 -360 1642 -60
rect -174 -2294 -82 -2271
rect -21 -374 636 -372
rect -21 -383 1236 -374
rect -21 -388 1159 -383
rect -21 -437 178 -388
rect 237 -389 831 -388
rect 237 -437 501 -389
rect -21 -1860 46 -437
rect 161 -440 501 -437
rect 562 -439 831 -389
rect 892 -439 1159 -388
rect 562 -440 1159 -439
rect 161 -443 1159 -440
rect 161 -453 252 -443
rect 486 -453 577 -443
rect 816 -454 907 -443
rect 1145 -444 1159 -443
rect 1222 -444 1236 -383
rect 1145 -454 1236 -444
rect 1551 -440 1641 -360
rect 3293 -370 3384 -60
rect 96 -536 168 -525
rect -21 -2245 47 -1860
rect 96 -2110 100 -536
rect 146 -540 168 -536
rect 156 -2103 168 -540
rect 146 -2110 168 -2103
rect 96 -2121 168 -2110
rect 264 -536 336 -525
rect 310 -539 336 -536
rect 320 -2103 336 -539
rect 310 -2110 336 -2103
rect 264 -2121 336 -2110
rect 428 -536 500 -525
rect 474 -539 500 -536
rect 487 -2103 500 -539
rect 474 -2110 500 -2103
rect 428 -2121 500 -2110
rect 592 -536 664 -525
rect 638 -539 664 -536
rect 654 -2103 664 -539
rect 638 -2110 664 -2103
rect 592 -2121 664 -2110
rect 755 -536 827 -525
rect 755 -2110 756 -536
rect 802 -539 827 -536
rect 816 -2103 827 -539
rect 802 -2110 827 -2103
rect 755 -2121 827 -2110
rect 920 -536 992 -525
rect 966 -539 992 -536
rect 983 -2103 992 -539
rect 966 -2110 992 -2103
rect 920 -2121 992 -2110
rect 1084 -536 1156 -525
rect 1130 -539 1156 -536
rect 1148 -2103 1156 -539
rect 1130 -2110 1156 -2103
rect 1084 -2121 1156 -2110
rect 1247 -536 1319 -525
rect 1247 -2110 1248 -536
rect 1294 -539 1319 -536
rect 1310 -2103 1319 -539
rect 1294 -2110 1319 -2103
rect 1247 -2121 1319 -2110
rect 1389 -536 1461 -525
rect 1389 -540 1412 -536
rect 1389 -2104 1399 -540
rect 1389 -2110 1412 -2104
rect 1458 -2110 1461 -536
rect 1389 -2121 1461 -2110
rect 321 -2243 413 -2233
rect 651 -2243 743 -2233
rect 979 -2243 1071 -2233
rect 1306 -2243 1398 -2233
rect 321 -2245 1398 -2243
rect -21 -2247 1398 -2245
rect -21 -2250 1399 -2247
rect -21 -2252 1322 -2250
rect -174 -2380 -79 -2294
rect -21 -2300 336 -2252
rect 396 -2300 667 -2252
rect 727 -2300 996 -2252
rect 1056 -2298 1322 -2252
rect 1382 -2298 1399 -2250
rect 1551 -2249 1567 -440
rect 1628 -2249 1641 -440
rect 1551 -2294 1641 -2249
rect 1721 -374 2378 -372
rect 1721 -380 2978 -374
rect 1721 -437 1917 -380
rect 1980 -388 2978 -380
rect 1980 -389 2573 -388
rect 1721 -1860 1788 -437
rect 1903 -439 1917 -437
rect 1980 -439 2243 -389
rect 1903 -440 2243 -439
rect 2304 -439 2573 -389
rect 2634 -389 2978 -388
rect 2634 -439 2903 -389
rect 2304 -440 2903 -439
rect 2964 -440 2978 -389
rect 1903 -443 2978 -440
rect 1903 -453 1994 -443
rect 2228 -453 2319 -443
rect 2558 -454 2649 -443
rect 2887 -454 2978 -443
rect 3293 -440 3383 -370
rect 1838 -536 1910 -525
rect 1721 -2245 1789 -1860
rect 1838 -2110 1842 -536
rect 1888 -540 1910 -536
rect 1898 -2103 1910 -540
rect 1888 -2110 1910 -2103
rect 1838 -2121 1910 -2110
rect 2006 -536 2078 -525
rect 2052 -539 2078 -536
rect 2062 -2103 2078 -539
rect 2052 -2110 2078 -2103
rect 2006 -2121 2078 -2110
rect 2170 -536 2242 -525
rect 2216 -539 2242 -536
rect 2229 -2103 2242 -539
rect 2216 -2110 2242 -2103
rect 2170 -2121 2242 -2110
rect 2334 -536 2406 -525
rect 2380 -539 2406 -536
rect 2396 -2103 2406 -539
rect 2380 -2110 2406 -2103
rect 2334 -2121 2406 -2110
rect 2497 -536 2569 -525
rect 2497 -2110 2498 -536
rect 2544 -539 2569 -536
rect 2558 -2103 2569 -539
rect 2544 -2110 2569 -2103
rect 2497 -2121 2569 -2110
rect 2662 -536 2734 -525
rect 2708 -539 2734 -536
rect 2725 -2103 2734 -539
rect 2708 -2110 2734 -2103
rect 2662 -2121 2734 -2110
rect 2826 -536 2898 -525
rect 2872 -539 2898 -536
rect 2890 -2103 2898 -539
rect 2872 -2110 2898 -2103
rect 2826 -2121 2898 -2110
rect 2989 -536 3061 -525
rect 2989 -2110 2990 -536
rect 3036 -539 3061 -536
rect 3052 -2103 3061 -539
rect 3036 -2110 3061 -2103
rect 2989 -2121 3061 -2110
rect 3131 -536 3203 -525
rect 3131 -540 3154 -536
rect 3131 -2104 3141 -540
rect 3131 -2110 3154 -2104
rect 3200 -2110 3203 -536
rect 3131 -2121 3203 -2110
rect 2063 -2243 2155 -2233
rect 2393 -2243 2485 -2233
rect 2721 -2243 2813 -2233
rect 3048 -2243 3140 -2233
rect 2063 -2245 3140 -2243
rect 1721 -2247 3140 -2245
rect 1721 -2250 3141 -2247
rect 1721 -2252 3064 -2250
rect 1056 -2300 1399 -2298
rect -21 -2313 1399 -2300
rect -175 -2382 63 -2380
rect 1548 -2382 1643 -2294
rect 1721 -2300 2078 -2252
rect 2138 -2300 2409 -2252
rect 2469 -2300 2738 -2252
rect 2798 -2298 3064 -2252
rect 3124 -2298 3141 -2250
rect 3293 -2249 3309 -440
rect 3370 -2249 3383 -440
rect 3293 -2297 3383 -2249
rect 2798 -2300 3141 -2298
rect 1721 -2313 3141 -2300
rect 3289 -2382 3384 -2297
rect -175 -2394 3384 -2382
rect -175 -2471 3380 -2394
<< via1 >>
rect 103 150 155 1713
rect 267 150 319 1714
rect 434 150 486 1714
rect 601 150 653 1714
rect 763 150 815 1714
rect 930 150 982 1714
rect 1095 150 1147 1714
rect 1257 150 1309 1714
rect 1398 149 1450 1713
rect 1320 3 1383 8
rect 1320 -45 1321 3
rect 1321 -45 1381 3
rect 1381 -45 1383 3
rect 1320 -51 1383 -45
rect 1845 150 1887 1713
rect 1887 150 1897 1713
rect 2009 150 2051 1714
rect 2051 150 2061 1714
rect 2176 150 2215 1714
rect 2215 150 2228 1714
rect 2343 150 2379 1714
rect 2379 150 2395 1714
rect 2505 150 2543 1714
rect 2543 150 2557 1714
rect 2672 150 2707 1714
rect 2707 150 2724 1714
rect 2837 150 2871 1714
rect 2871 150 2889 1714
rect 2999 150 3035 1714
rect 3035 150 3051 1714
rect 3140 149 3153 1713
rect 3153 149 3192 1713
rect 2078 1 2142 8
rect 2078 -47 2137 1
rect 2137 -47 2142 1
rect 2078 -48 2142 -47
rect 1159 -389 1222 -383
rect 1159 -440 1161 -389
rect 1161 -440 1222 -389
rect 1159 -444 1222 -440
rect 104 -2103 146 -540
rect 146 -2103 156 -540
rect 268 -2103 310 -539
rect 310 -2103 320 -539
rect 435 -2103 474 -539
rect 474 -2103 487 -539
rect 602 -2103 638 -539
rect 638 -2103 654 -539
rect 764 -2103 802 -539
rect 802 -2103 816 -539
rect 931 -2103 966 -539
rect 966 -2103 983 -539
rect 1096 -2103 1130 -539
rect 1130 -2103 1148 -539
rect 1258 -2103 1294 -539
rect 1294 -2103 1310 -539
rect 1399 -2104 1412 -540
rect 1412 -2104 1451 -540
rect 1917 -388 1980 -380
rect 1917 -437 1920 -388
rect 1920 -437 1979 -388
rect 1979 -437 1980 -388
rect 1917 -439 1980 -437
rect 1846 -2103 1888 -540
rect 1888 -2103 1898 -540
rect 2010 -2103 2052 -539
rect 2052 -2103 2062 -539
rect 2177 -2103 2216 -539
rect 2216 -2103 2229 -539
rect 2344 -2103 2380 -539
rect 2380 -2103 2396 -539
rect 2506 -2103 2544 -539
rect 2544 -2103 2558 -539
rect 2673 -2103 2708 -539
rect 2708 -2103 2725 -539
rect 2838 -2103 2872 -539
rect 2872 -2103 2890 -539
rect 3000 -2103 3036 -539
rect 3036 -2103 3052 -539
rect 3141 -2104 3154 -540
rect 3154 -2104 3193 -540
<< metal2 >>
rect 95 1713 167 1728
rect 95 150 103 1713
rect 155 150 167 1713
rect 95 132 167 150
rect 263 1714 335 1728
rect 263 150 267 1714
rect 319 150 335 1714
rect 263 132 335 150
rect 427 1714 499 1728
rect 427 150 434 1714
rect 486 150 499 1714
rect 427 132 499 150
rect 591 1714 663 1728
rect 591 150 601 1714
rect 653 150 663 1714
rect 591 132 663 150
rect 754 1714 826 1728
rect 754 150 763 1714
rect 815 150 826 1714
rect 754 132 826 150
rect 919 1714 991 1728
rect 919 150 930 1714
rect 982 150 991 1714
rect 919 132 991 150
rect 1083 1714 1155 1728
rect 1083 150 1095 1714
rect 1147 150 1155 1714
rect 1083 132 1155 150
rect 1246 1714 1318 1728
rect 1246 150 1257 1714
rect 1309 150 1318 1714
rect 1246 132 1318 150
rect 1388 1713 1460 1728
rect 1388 149 1398 1713
rect 1450 149 1460 1713
rect 1388 132 1460 149
rect 1837 1713 1909 1728
rect 1837 150 1845 1713
rect 1897 150 1909 1713
rect 1837 132 1909 150
rect 2005 1714 2077 1728
rect 2005 150 2009 1714
rect 2061 150 2077 1714
rect 2005 132 2077 150
rect 2169 1714 2241 1728
rect 2169 150 2176 1714
rect 2228 150 2241 1714
rect 2169 132 2241 150
rect 2333 1714 2405 1728
rect 2333 150 2343 1714
rect 2395 150 2405 1714
rect 2333 132 2405 150
rect 2496 1714 2568 1728
rect 2496 150 2505 1714
rect 2557 150 2568 1714
rect 2496 132 2568 150
rect 2661 1714 2733 1728
rect 2661 150 2672 1714
rect 2724 150 2733 1714
rect 2661 132 2733 150
rect 2825 1714 2897 1728
rect 2825 150 2837 1714
rect 2889 150 2897 1714
rect 2825 132 2897 150
rect 2988 1714 3060 1728
rect 2988 150 2999 1714
rect 3051 150 3060 1714
rect 2988 132 3060 150
rect 3130 1713 3202 1728
rect 3130 149 3140 1713
rect 3192 149 3202 1713
rect 3130 132 3202 149
rect 1305 8 1398 20
rect 1305 -51 1320 8
rect 1383 -51 1398 8
rect 2061 8 2152 20
rect 2061 -19 2078 8
rect 1305 -60 1398 -51
rect 2060 -48 2078 -19
rect 2142 -19 2152 8
rect 2142 -48 2154 -19
rect 2060 -101 2154 -48
rect 1490 -105 2154 -101
rect 1489 -169 2154 -105
rect 1489 -170 2152 -169
rect 1489 -374 1558 -170
rect 1147 -383 1558 -374
rect 1147 -444 1159 -383
rect 1222 -443 1558 -383
rect 1903 -380 1996 -373
rect 1903 -439 1917 -380
rect 1980 -439 1996 -380
rect 1222 -444 1236 -443
rect 1147 -452 1236 -444
rect 1903 -453 1996 -439
rect 96 -540 168 -525
rect 96 -2103 104 -540
rect 156 -2103 168 -540
rect 96 -2121 168 -2103
rect 264 -539 336 -525
rect 264 -2103 268 -539
rect 320 -2103 336 -539
rect 264 -2121 336 -2103
rect 428 -539 500 -525
rect 428 -2103 435 -539
rect 487 -2103 500 -539
rect 428 -2121 500 -2103
rect 592 -539 664 -525
rect 592 -2103 602 -539
rect 654 -2103 664 -539
rect 592 -2121 664 -2103
rect 755 -539 827 -525
rect 755 -2103 764 -539
rect 816 -2103 827 -539
rect 755 -2121 827 -2103
rect 920 -539 992 -525
rect 920 -2103 931 -539
rect 983 -2103 992 -539
rect 920 -2121 992 -2103
rect 1084 -539 1156 -525
rect 1084 -2103 1096 -539
rect 1148 -2103 1156 -539
rect 1084 -2121 1156 -2103
rect 1247 -539 1319 -525
rect 1247 -2103 1258 -539
rect 1310 -2103 1319 -539
rect 1247 -2121 1319 -2103
rect 1389 -540 1461 -525
rect 1389 -2104 1399 -540
rect 1451 -2104 1461 -540
rect 1389 -2121 1461 -2104
rect 1838 -540 1910 -525
rect 1838 -2103 1846 -540
rect 1898 -2103 1910 -540
rect 1838 -2121 1910 -2103
rect 2006 -539 2078 -525
rect 2006 -2103 2010 -539
rect 2062 -2103 2078 -539
rect 2006 -2121 2078 -2103
rect 2170 -539 2242 -525
rect 2170 -2103 2177 -539
rect 2229 -2103 2242 -539
rect 2170 -2121 2242 -2103
rect 2334 -539 2406 -525
rect 2334 -2103 2344 -539
rect 2396 -2103 2406 -539
rect 2334 -2121 2406 -2103
rect 2497 -539 2569 -525
rect 2497 -2103 2506 -539
rect 2558 -2103 2569 -539
rect 2497 -2121 2569 -2103
rect 2662 -539 2734 -525
rect 2662 -2103 2673 -539
rect 2725 -2103 2734 -539
rect 2662 -2121 2734 -2103
rect 2826 -539 2898 -525
rect 2826 -2103 2838 -539
rect 2890 -2103 2898 -539
rect 2826 -2121 2898 -2103
rect 2989 -539 3061 -525
rect 2989 -2103 3000 -539
rect 3052 -2103 3061 -539
rect 2989 -2121 3061 -2103
rect 3131 -540 3203 -525
rect 3131 -2104 3141 -540
rect 3193 -2104 3203 -540
rect 3131 -2121 3203 -2104
<< via2 >>
rect 1320 -51 1383 8
rect 1917 -439 1980 -380
<< metal3 >>
rect 1305 8 1398 20
rect 1305 -51 1320 8
rect 1383 -51 1398 8
rect 1305 -60 1398 -51
rect 1314 -149 1392 -60
rect 1314 -229 1992 -149
rect 1910 -373 1991 -229
rect 1903 -380 1996 -373
rect 1903 -439 1917 -380
rect 1980 -439 1996 -380
rect 1903 -453 1996 -439
use pfet_03v3_CSJ2S3  pfet_03v3_CSJ2S3_0
timestamp 1757727097
transform 1 0 778 0 1 930
box -778 -930 778 930
use pfet_03v3_CSJ2S3  pfet_03v3_CSJ2S3_1
timestamp 1757727097
transform 1 0 2520 0 1 930
box -778 -930 778 930
use pfet_03v3_CSJ2S3  pfet_03v3_CSJ2S3_2
timestamp 1757727097
transform 1 0 2521 0 1 -1323
box -778 -930 778 930
use pfet_03v3_CSJ2S3  pfet_03v3_CSJ2S3_3
timestamp 1757727097
transform 1 0 779 0 1 -1323
box -778 -930 778 930
<< end >>
