magic
tech gf180mcuD
magscale 1 10
timestamp 1757241197
<< nwell >>
rect 2686 1955 3254 2198
rect 2684 -115 3255 1955
<< pwell >>
rect 3288 1954 3765 2198
rect 3284 1946 3765 1954
rect 3284 792 3760 1946
rect 3284 741 4128 792
rect 3284 95 4125 741
rect 3285 -114 4124 95
<< nmos >>
rect 3432 215 3488 1815
rect 3592 215 3648 1815
rect 3924 215 3980 615
<< pmos >>
rect 2858 225 2914 1825
rect 3018 225 3074 1825
<< ndiff >>
rect 3344 1802 3432 1815
rect 3344 228 3357 1802
rect 3403 228 3432 1802
rect 3344 215 3432 228
rect 3488 1802 3592 1815
rect 3488 228 3517 1802
rect 3563 228 3592 1802
rect 3488 215 3592 228
rect 3648 1802 3736 1815
rect 3648 228 3677 1802
rect 3723 228 3736 1802
rect 3648 215 3736 228
rect 3834 596 3924 615
rect 3834 240 3849 596
rect 3895 240 3924 596
rect 3834 215 3924 240
rect 3980 596 4077 615
rect 3980 240 4013 596
rect 4059 240 4077 596
rect 3980 215 4077 240
rect 4010 214 4077 215
<< pdiff >>
rect 2770 1812 2858 1825
rect 2770 238 2783 1812
rect 2829 238 2858 1812
rect 2770 225 2858 238
rect 2914 1812 3018 1825
rect 2914 238 2943 1812
rect 2989 238 3018 1812
rect 2914 225 3018 238
rect 3074 1812 3162 1825
rect 3074 238 3103 1812
rect 3149 238 3162 1812
rect 3074 225 3162 238
<< ndiffc >>
rect 3357 228 3403 1802
rect 3517 228 3563 1802
rect 3677 228 3723 1802
rect 3849 240 3895 596
rect 4013 240 4059 596
<< pdiffc >>
rect 2783 238 2829 1812
rect 2943 238 2989 1812
rect 3103 238 3149 1812
<< psubdiff >>
rect 3344 43 4114 85
rect 3344 -51 3443 43
rect 4058 -51 4114 43
rect 3344 -74 4114 -51
<< nsubdiff >>
rect 2744 2147 3205 2170
rect 2744 2030 2788 2147
rect 3183 2030 3205 2147
rect 2744 2007 3205 2030
<< psubdiffcont >>
rect 3443 -51 4058 43
<< nsubdiffcont >>
rect 2788 2030 3183 2147
<< polysilicon >>
rect 2858 1864 3076 1920
rect 2858 1825 2914 1864
rect 3018 1825 3074 1864
rect 3401 1856 3490 1947
rect 3593 1859 3682 1945
rect 3432 1815 3488 1856
rect 3592 1854 3682 1859
rect 3592 1815 3648 1854
rect 2858 181 2914 225
rect 3018 181 3074 225
rect 3901 652 3993 743
rect 3924 615 3980 652
rect 3432 171 3488 215
rect 3592 171 3648 215
rect 3924 169 3980 215
<< metal1 >>
rect 2744 2147 3205 2170
rect 2744 2030 2788 2147
rect 3183 2030 3205 2147
rect 2744 2007 3205 2030
rect 2783 1812 2829 1823
rect 2943 1812 2989 1823
rect 2829 1765 2835 1780
rect 2829 1697 2835 1711
rect 2783 227 2829 238
rect 3103 1812 3149 1823
rect 3357 1802 3403 1813
rect 3149 1769 3155 1782
rect 2989 335 2998 350
rect 2996 281 2998 335
rect 2989 269 2998 281
rect 2943 227 2989 238
rect 3149 1699 3155 1715
rect 3103 227 3149 238
rect 3517 1802 3563 1813
rect 3512 340 3517 352
rect 3677 1802 3723 1813
rect 3563 340 3571 352
rect 3512 286 3516 340
rect 3569 286 3571 340
rect 3512 271 3517 286
rect 3357 217 3403 228
rect 3563 271 3571 286
rect 3517 217 3563 228
rect 3677 217 3723 228
rect 3838 596 3908 609
rect 3838 340 3849 596
rect 3895 340 3908 596
rect 3838 286 3845 340
rect 3898 286 3908 340
rect 3838 240 3849 286
rect 3895 240 3908 286
rect 3838 222 3908 240
rect 4002 596 4072 609
rect 4002 240 4013 596
rect 4059 240 4072 596
rect 4002 222 4072 240
rect 3344 43 4114 85
rect 3344 -51 3443 43
rect 4058 -51 4114 43
rect 3344 -74 4114 -51
<< via1 >>
rect 2783 1711 2829 1765
rect 2829 1711 2835 1765
rect 3103 1715 3149 1769
rect 3149 1715 3155 1769
rect 2943 281 2989 335
rect 2989 281 2996 335
rect 3516 286 3517 340
rect 3517 286 3563 340
rect 3563 286 3569 340
rect 3845 286 3849 340
rect 3849 286 3895 340
rect 3895 286 3898 340
<< metal2 >>
rect 2779 1769 3165 1783
rect 2779 1765 3103 1769
rect 2779 1711 2783 1765
rect 2835 1715 3103 1765
rect 3155 1715 3165 1769
rect 2835 1711 3165 1715
rect 2779 1698 3165 1711
rect 2779 1697 2835 1698
rect 2937 340 3907 348
rect 2937 335 3516 340
rect 2937 281 2943 335
rect 2996 286 3516 335
rect 3569 286 3845 340
rect 3898 286 3907 340
rect 2996 281 3907 286
rect 2937 269 3907 281
<< labels >>
flabel metal1 3358 372 3397 609 0 FreeSans 160 0 0 0 VCM
port 1 nsew
flabel metal1 4008 275 4069 558 0 FreeSans 160 0 0 0 VIN
port 3 nsew
flabel metal2 2851 1702 3079 1766 0 FreeSans 160 0 0 0 VREF
port 4 nsew
flabel polysilicon 3402 1860 3488 1940 0 FreeSans 160 0 0 0 EN_VCM
port 5 nsew
flabel polysilicon 2870 1868 3072 1915 0 FreeSans 160 0 0 0 EN_VREF_Z
port 6 nsew
flabel metal2 3055 276 3438 339 0 FreeSans 160 0 0 0 Cbtm
port 7 nsew
flabel metal1 2770 2031 3194 2152 0 FreeSans 320 0 0 0 VDD
port 8 nsew
flabel polysilicon 3597 1860 3680 1938 0 FreeSans 160 0 0 0 EN_VSS
port 9 nsew
flabel polysilicon 3906 656 3989 734 0 FreeSans 160 0 0 0 EN_VIN
port 10 nsew
flabel metal1 3409 -57 4088 56 0 FreeSans 320 0 0 0 VSS
port 11 nsew
flabel metal1 3679 381 3719 1770 0 FreeSans 160 0 0 0 VREF_GND
port 2 nsew
<< end >>
