magic
tech gf180mcuD
magscale 1 5
timestamp 1757840551
use ppolyf_u_1k_MM5P8U  ppolyf_u_1k_MM5P8U_0
timestamp 1757840551
transform 1 0 838 0 1 1299
box -868 -1329 868 1329
<< end >>
