magic
tech gf180mcuD
magscale 1 10
timestamp 1757414101
<< nwell >>
rect -212 -216 212 216
<< pwell >>
rect -236 216 236 240
rect -236 -216 -212 216
rect 212 -216 236 216
rect -236 -240 236 -216
<< nsubdiff >>
rect -188 87 -100 100
rect -188 -87 -175 87
rect -129 -87 -100 87
rect -188 -100 -100 -87
rect 100 87 188 100
rect 100 -87 129 87
rect 175 -87 188 87
rect 100 -100 188 -87
<< nsubdiffcont >>
rect -175 -87 -129 87
rect 129 -87 175 87
<< nvaractor >>
rect -100 -100 100 100
<< polysilicon >>
rect -100 179 100 192
rect -100 133 -87 179
rect 87 133 100 179
rect -100 100 100 133
rect -100 -133 100 -100
rect -100 -179 -87 -133
rect 87 -179 100 -133
rect -100 -192 100 -179
<< polycontact >>
rect -87 133 87 179
rect -87 -179 87 -133
<< metal1 >>
rect -98 133 -87 179
rect 87 133 98 179
rect -175 87 -129 98
rect -175 -98 -129 -87
rect 129 87 175 98
rect 129 -98 175 -87
rect -98 -179 -87 -133
rect 87 -179 98 -133
<< properties >>
string gencell nmoscap_3p3
string library gf180mcu
string parameters w 1.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {nmoscap_3p3 nmoscap_6p0}
<< end >>
