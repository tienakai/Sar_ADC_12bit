magic
tech gf180mcuD
magscale 1 10
timestamp 1757750971
<< nwell >>
rect -111 -170 4560 1880
<< nsubdiff >>
rect 4429 1784 4530 1850
rect 4429 1626 4454 1784
rect 4430 40 4454 1626
rect 4510 40 4530 1784
rect 4430 -105 4530 40
<< nsubdiffcont >>
rect 4454 40 4510 1784
<< metal1 >>
rect 65 1705 156 1815
rect 408 1705 499 1816
rect 81 1704 156 1705
rect 750 1704 841 1815
rect 1092 1705 1183 1816
rect 1434 1705 1525 1816
rect 1776 1705 1867 1816
rect 2118 1704 2209 1815
rect 2460 1705 2551 1816
rect 2802 1705 2893 1816
rect 3144 1704 3235 1815
rect 3486 1705 3577 1816
rect 3828 1705 3919 1816
rect 4170 1704 4261 1815
rect 4429 1784 4530 1850
rect 4429 1626 4454 1784
rect 4430 40 4454 1626
rect 4510 40 4530 1784
rect 66 -73 157 38
rect 408 -72 499 39
rect 750 -72 841 39
rect 1092 -71 1183 40
rect 1434 -72 1525 39
rect 1776 -71 1867 40
rect 2118 -72 2209 39
rect 2460 -71 2551 40
rect 2802 -71 2893 40
rect 3143 -72 3234 39
rect 3486 -72 3577 39
rect 3827 -72 3918 39
rect 4171 -72 4262 39
rect 4430 -105 4530 40
use pfet_03v3_3WZPEW  pfet_03v3_3WZPEW_0
timestamp 1757750971
transform 1 0 2166 0 1 872
box -2276 -978 2276 978
<< end >>
