magic
tech gf180mcuD
magscale 1 10
timestamp 1757728578
<< pwell >>
rect 100 507 180 591
rect 258 510 339 591
rect 418 510 499 591
rect 579 510 660 591
rect 83 453 95 454
rect 81 442 95 453
rect 42 384 95 442
rect 81 372 95 384
rect 661 372 730 454
<< ndiff >>
rect 83 453 95 454
rect 81 442 95 453
rect 42 384 95 442
rect 81 372 95 384
rect 661 372 730 454
<< polysilicon >>
rect 100 570 180 591
rect 100 521 120 570
rect 167 521 180 570
rect 100 507 180 521
rect 258 575 339 591
rect 258 526 278 575
rect 326 526 339 575
rect 258 510 339 526
rect 418 576 499 591
rect 418 527 435 576
rect 483 527 499 576
rect 418 510 499 527
rect 579 575 660 591
rect 579 526 598 575
rect 646 526 660 575
rect 579 510 660 526
<< polycontact >>
rect 120 521 167 570
rect 278 526 326 575
rect 435 527 483 576
rect 598 526 646 575
<< metal1 >>
rect 100 576 660 591
rect 100 575 435 576
rect 100 570 278 575
rect 100 521 120 570
rect 167 531 278 570
rect 167 521 180 531
rect 100 510 180 521
rect 258 526 278 531
rect 326 531 435 575
rect 326 526 339 531
rect 258 510 339 526
rect 418 527 435 531
rect 483 575 660 576
rect 483 531 598 575
rect 483 527 499 531
rect 418 510 499 527
rect 579 526 598 531
rect 646 526 660 575
rect 579 510 660 526
rect 723 454 724 455
rect 83 453 95 454
rect 81 447 95 453
rect 37 442 95 447
rect 37 384 42 442
rect 37 379 95 384
rect 81 372 95 379
rect 345 444 420 454
rect 345 384 357 444
rect 411 384 420 444
rect 345 372 420 384
rect 661 443 730 454
rect 661 384 672 443
rect 724 384 730 443
rect 661 372 730 384
<< via1 >>
rect 42 384 95 442
rect 357 384 411 444
rect 672 384 724 443
<< metal2 >>
rect 661 454 730 456
rect 29 444 730 454
rect 29 442 357 444
rect 29 384 42 442
rect 95 384 357 442
rect 411 443 730 444
rect 411 384 672 443
rect 724 384 730 443
rect 29 372 730 384
use nfet_03v3_N2UC85  nfet_03v3_N2UC85_0
timestamp 1757728578
transform 1 0 380 0 1 268
box -380 -268 380 268
<< end >>
