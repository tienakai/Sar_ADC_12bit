magic
tech gf180mcuD
magscale 1 10
timestamp 1757866589
<< metal1 >>
rect 36919 46464 42925 46478
rect 36919 46449 42787 46464
rect 36919 46360 36933 46449
rect 37131 46360 42787 46449
rect 36919 46358 42787 46360
rect 42915 46358 42925 46464
rect 36919 46342 42925 46358
rect 39691 39747 42675 39767
rect 39691 39742 42536 39747
rect 39691 39652 39731 39742
rect 39884 39654 42536 39742
rect 42670 39654 42675 39747
rect 39884 39652 42675 39654
rect 39691 39641 42675 39652
rect 39691 39640 42605 39641
rect 39700 39639 39901 39640
rect 39690 38880 42425 38893
rect 39690 38870 42285 38880
rect 39690 38791 39722 38870
rect 39865 38791 42285 38870
rect 39690 38786 42285 38791
rect 42410 38786 42425 38880
rect 39690 38773 42425 38786
rect 42272 38770 42425 38773
rect 39687 38659 42168 38678
rect 39687 38574 39723 38659
rect 39855 38574 42043 38659
rect 39687 38566 42043 38574
rect 42149 38566 42168 38659
rect 39687 38553 42168 38566
rect 39687 38549 42156 38553
rect 24528 37664 24650 37676
rect 24528 37579 24550 37664
rect 24637 37579 24650 37664
rect 23343 37449 23465 37465
rect 23343 37371 23357 37449
rect 23441 37371 23465 37449
rect 23343 36035 23465 37371
rect 23564 37438 23683 37448
rect 23564 37370 23579 37438
rect 23668 37370 23683 37438
rect 23564 36340 23683 37370
rect 24528 36722 24650 37579
rect 24802 37664 24913 37667
rect 24802 37647 24915 37664
rect 24802 37568 24815 37647
rect 24898 37568 24915 37647
rect 24802 37538 24915 37568
rect 24528 36637 24545 36722
rect 24632 36637 24650 36722
rect 24803 36811 24915 37538
rect 24803 36728 24819 36811
rect 24903 36728 24915 36811
rect 24803 36717 24915 36728
rect 25058 37655 25171 37676
rect 25058 37576 25070 37655
rect 25161 37576 25171 37655
rect 25058 36818 25171 37576
rect 39888 37529 42461 37534
rect 39700 37514 42461 37529
rect 39700 37513 42346 37514
rect 39700 37406 39712 37513
rect 39888 37418 42346 37513
rect 42447 37418 42461 37514
rect 39888 37406 42461 37418
rect 39700 37394 42461 37406
rect 25058 36732 25081 36818
rect 25157 36732 25171 36818
rect 25058 36710 25171 36732
rect 24528 36614 24650 36637
rect 23343 35933 23359 36035
rect 23446 35933 23465 36035
rect 23343 35919 23465 35933
rect 23558 36316 23683 36340
rect 23558 36050 23682 36316
rect 23558 36049 24391 36050
rect 23558 36038 24446 36049
rect 23558 35937 24333 36038
rect 24432 35937 24446 36038
rect 23558 35921 24446 35937
rect 27556 35579 29933 35585
rect 27556 35575 41104 35579
rect 27556 35507 27569 35575
rect 27674 35574 41104 35575
rect 27674 35516 40967 35574
rect 41091 35516 41104 35574
rect 27674 35507 41104 35516
rect 27556 35503 41104 35507
rect 27556 35502 41102 35503
rect 27556 35495 29933 35502
rect 27561 35372 30122 35378
rect 27561 35358 41319 35372
rect 27561 35288 27578 35358
rect 27663 35347 41319 35358
rect 27663 35288 41199 35347
rect 41294 35288 41319 35347
rect 27561 35275 41319 35288
rect 30000 35273 41319 35275
rect 27569 35171 30357 35175
rect 41378 35171 41522 35174
rect 27569 35162 41522 35171
rect 27569 35098 27580 35162
rect 27667 35102 41404 35162
rect 41502 35102 41522 35162
rect 27667 35098 41522 35102
rect 27569 35082 41522 35098
rect 27569 35081 30357 35082
rect 41378 35081 41522 35082
rect 27567 34996 30598 34998
rect 41490 34996 41747 34998
rect 27567 34985 41747 34996
rect 27567 34911 27586 34985
rect 27661 34974 41747 34985
rect 27661 34914 41627 34974
rect 41716 34914 41747 34974
rect 27661 34911 41747 34914
rect 27567 34900 41747 34911
rect 27567 34899 41504 34900
rect 30589 34898 41504 34899
rect 41493 34816 42003 34818
rect 30816 34806 42003 34816
rect 27558 34801 42003 34806
rect 27558 34795 41887 34801
rect 27558 34719 27583 34795
rect 27661 34727 41887 34795
rect 41988 34727 42003 34801
rect 27661 34719 42003 34727
rect 27558 34708 42003 34719
rect 27558 34707 41510 34708
rect 30816 34706 41510 34707
rect 41597 34617 42224 34620
rect 31025 34613 42224 34617
rect 27540 34600 42224 34613
rect 27540 34597 42093 34600
rect 27540 34529 27555 34597
rect 27651 34533 42093 34597
rect 42197 34533 42224 34600
rect 27651 34529 42224 34533
rect 27540 34520 42224 34529
rect 27540 34519 41665 34520
rect 27540 34515 31034 34519
<< via1 >>
rect 36933 46360 37131 46449
rect 42787 46358 42915 46464
rect 39731 39652 39884 39742
rect 42536 39654 42670 39747
rect 39722 38791 39865 38870
rect 42285 38786 42410 38880
rect 39723 38574 39855 38659
rect 42043 38566 42149 38659
rect 24550 37579 24637 37664
rect 23357 37371 23441 37449
rect 23579 37370 23668 37438
rect 24815 37568 24898 37647
rect 24545 36637 24632 36722
rect 24819 36728 24903 36811
rect 25070 37576 25161 37655
rect 39712 37406 39888 37513
rect 42346 37418 42447 37514
rect 25081 36732 25157 36818
rect 23359 35933 23446 36035
rect 24333 35937 24432 36038
rect 27569 35507 27674 35575
rect 40967 35516 41091 35574
rect 27578 35288 27663 35358
rect 41199 35288 41294 35347
rect 27580 35098 27667 35162
rect 41404 35102 41502 35162
rect 27586 34911 27661 34985
rect 41627 34914 41716 34974
rect 27583 34719 27661 34795
rect 41887 34727 41988 34801
rect 27555 34529 27651 34597
rect 42093 34533 42197 34600
<< metal2 >>
rect 32860 75838 32964 75843
rect 30588 75814 32964 75838
rect 30588 75732 30617 75814
rect 31137 75732 32964 75814
rect 30588 75719 32964 75732
rect 30580 74702 32761 74724
rect 30580 74613 30623 74702
rect 31157 74613 32761 74702
rect 30580 74597 32761 74613
rect 32401 73593 32517 73595
rect 30584 73581 32517 73593
rect 30584 73500 30621 73581
rect 31171 73500 32517 73581
rect 30584 73474 32517 73500
rect 32252 72471 32329 72473
rect 30595 72462 32329 72471
rect 30595 72383 30628 72462
rect 31170 72418 32329 72462
rect 31170 72383 32331 72418
rect 30595 72365 32331 72383
rect 32252 71872 32331 72365
rect 30591 71338 32178 71356
rect 30591 71259 30617 71338
rect 31166 71259 32178 71338
rect 30591 71243 32178 71259
rect 32082 71013 32177 71243
rect 31926 70234 32006 70236
rect 30591 70213 32006 70234
rect 30591 70136 30676 70213
rect 31145 70136 32006 70213
rect 30591 70121 32006 70136
rect 30589 69109 31724 69114
rect 30589 69093 31833 69109
rect 30589 69019 30624 69093
rect 31155 69019 31833 69093
rect 30589 69004 31833 69019
rect 30589 69001 31189 69004
rect 31393 68004 31664 68005
rect 30588 67980 31664 68004
rect 30588 67894 30638 67980
rect 31156 67894 31664 67980
rect 30588 67883 31664 67894
rect 31393 67881 31664 67883
rect 31401 66874 31487 66875
rect 30733 66850 31487 66874
rect 30733 66776 30806 66850
rect 31147 66776 31487 66850
rect 30733 66761 31487 66776
rect 31054 65755 31187 65756
rect 31009 65740 31187 65755
rect 31009 65664 31039 65740
rect 31172 65664 31187 65740
rect 31009 65642 31187 65664
rect 31009 64901 31097 65642
rect 31401 65135 31487 66761
rect 31398 65090 31487 65135
rect 31009 64900 31293 64901
rect 31009 64811 31334 64900
rect 31014 64620 31168 64636
rect 31014 64535 31030 64620
rect 31149 64535 31168 64620
rect 31014 60555 31168 64535
rect 31257 60701 31334 64811
rect 31398 63241 31483 65090
rect 31398 60842 31484 63241
rect 31571 60995 31664 67881
rect 31756 61154 31833 69004
rect 31926 61314 32006 70121
rect 32083 61502 32173 71013
rect 32252 61730 32333 71872
rect 32401 71695 32517 73474
rect 32401 61934 32518 71695
rect 32623 70871 32761 74597
rect 32623 62163 32773 70871
rect 32860 63294 32964 75719
rect 32860 62341 32965 63294
rect 32860 62340 42822 62341
rect 32860 62235 43128 62340
rect 32860 62233 42822 62235
rect 32622 62162 41482 62163
rect 32622 62160 41595 62162
rect 32622 62013 42907 62160
rect 32623 62012 42907 62013
rect 32623 62011 32773 62012
rect 32400 61817 42644 61934
rect 32401 61816 32518 61817
rect 42186 61811 42644 61817
rect 32252 61726 41575 61730
rect 32252 61724 42174 61726
rect 32252 61588 42438 61724
rect 32252 61586 32423 61588
rect 42303 61585 42438 61588
rect 32083 61501 41789 61502
rect 32083 61411 42218 61501
rect 41522 61410 42218 61411
rect 41292 61314 41903 61315
rect 31926 61234 42022 61314
rect 31926 61233 32006 61234
rect 41292 61231 42022 61234
rect 31755 61153 41756 61154
rect 31755 61077 41837 61153
rect 31756 61076 31833 61077
rect 31571 60994 41335 60995
rect 31571 60902 41703 60994
rect 31571 60901 41310 60902
rect 31397 60841 41239 60842
rect 31397 60763 41552 60841
rect 31398 60757 31484 60763
rect 35506 60702 41317 60703
rect 35506 60701 41409 60702
rect 31257 60624 41409 60701
rect 35506 60623 41409 60624
rect 41122 60565 41236 60567
rect 31445 60555 41238 60565
rect 14432 60497 14576 60502
rect 14432 60359 20761 60497
rect 31014 60408 41238 60555
rect 31014 60400 40583 60408
rect 31014 60396 31168 60400
rect 14432 57877 14576 60359
rect 38108 59817 38219 59847
rect 38108 59699 38138 59817
rect 38108 59673 38219 59699
rect 12388 57736 14576 57877
rect 12388 56840 12512 57736
rect 12368 56678 12523 56689
rect 12368 56577 12384 56678
rect 12507 56577 12523 56678
rect 12368 56560 12523 56577
rect 12504 56055 12656 56180
rect 41122 55637 41236 60408
rect 40577 55102 40708 55108
rect 41122 55102 41244 55637
rect 40572 54980 41244 55102
rect 41328 55556 41408 60623
rect 40577 51753 40728 54980
rect 41328 54921 41411 55556
rect 40846 54838 41412 54921
rect 40849 52230 40970 54838
rect 41328 54837 41411 54838
rect 41470 54766 41552 60763
rect 41610 55217 41702 60902
rect 41062 54748 41552 54766
rect 41060 54682 41552 54748
rect 40849 52052 40973 52230
rect 36916 46449 37158 46478
rect 36916 46360 36933 46449
rect 37131 46360 37158 46449
rect 36916 46300 37158 46360
rect 23347 39699 25867 39818
rect 39700 39742 39901 39756
rect 23350 39255 23469 39699
rect 39700 39652 39731 39742
rect 39884 39652 39901 39742
rect 39700 39639 39901 39652
rect 23347 37884 23469 39255
rect 23562 39274 23618 39275
rect 23562 39271 25072 39274
rect 23562 39155 25845 39271
rect 23562 39143 23684 39155
rect 25024 39154 25845 39155
rect 23347 37449 23466 37884
rect 23564 37450 23684 39143
rect 39690 38870 39894 38893
rect 39690 38791 39722 38870
rect 39865 38791 39894 38870
rect 39690 38773 39894 38791
rect 24798 38745 25860 38746
rect 24526 38624 25860 38745
rect 39690 38659 39888 38675
rect 24526 38623 25588 38624
rect 24527 37664 24649 38623
rect 39690 38574 39723 38659
rect 39855 38574 39888 38659
rect 39690 38553 39888 38574
rect 40577 38287 40727 51753
rect 40850 44846 40973 52052
rect 40850 44791 40975 44846
rect 40576 38234 40727 38287
rect 24803 38209 24908 38210
rect 24803 38208 25132 38209
rect 24803 38133 25871 38208
rect 24527 37579 24550 37664
rect 24637 37579 24649 37664
rect 24527 37564 24649 37579
rect 24802 38091 25871 38133
rect 24802 38089 25132 38091
rect 24802 37647 24908 38089
rect 24802 37568 24815 37647
rect 24898 37617 24908 37647
rect 25054 37655 25873 37667
rect 24898 37568 24907 37617
rect 24802 37540 24907 37568
rect 25054 37576 25070 37655
rect 25161 37576 25873 37655
rect 25054 37554 25873 37576
rect 23347 37371 23357 37449
rect 23441 37371 23466 37449
rect 23347 37362 23466 37371
rect 23563 37438 23684 37450
rect 23563 37370 23579 37438
rect 23668 37436 23684 37438
rect 39700 37513 39919 37529
rect 23668 37370 23683 37436
rect 39700 37406 39712 37513
rect 39888 37406 39919 37513
rect 39700 37394 39919 37406
rect 23563 37354 23683 37370
rect 40576 37306 40720 38234
rect 40852 37529 40975 44791
rect 41060 37717 41150 54682
rect 41470 54681 41552 54682
rect 41609 55176 41702 55217
rect 41609 54594 41700 55176
rect 41759 54851 41837 61077
rect 41759 54828 41847 54851
rect 41225 54503 41700 54594
rect 41225 52174 41316 54503
rect 41760 54445 41847 54828
rect 41905 54608 42022 61231
rect 42088 54608 42218 61410
rect 41424 54357 41847 54445
rect 41225 44251 41318 52174
rect 41225 38247 41319 44251
rect 41225 37877 41320 38247
rect 41425 38064 41513 54357
rect 41760 54355 41847 54357
rect 41906 54265 42011 54608
rect 41597 54160 42011 54265
rect 42087 54394 42218 54608
rect 41597 38230 41700 54160
rect 42087 54105 42217 54394
rect 42082 54104 42217 54105
rect 42073 54103 42217 54104
rect 41774 53959 42217 54103
rect 41774 38475 41918 53959
rect 42303 53898 42440 61585
rect 42023 53896 42440 53898
rect 42022 53760 42440 53896
rect 42022 39537 42160 53760
rect 42303 53756 42440 53760
rect 42501 53906 42644 61811
rect 42501 53700 42645 53906
rect 42752 53760 42907 62012
rect 42752 53745 42912 53760
rect 42273 53699 42645 53700
rect 42272 53556 42645 53699
rect 42272 42519 42427 53556
rect 42753 53457 42912 53745
rect 42517 53298 42914 53457
rect 42022 38733 42172 39537
rect 42272 38880 42428 42519
rect 42517 39747 42676 53298
rect 42753 53297 42912 53298
rect 42999 53232 43128 62235
rect 42765 53073 43128 53232
rect 42766 48024 42925 53073
rect 42766 48006 42926 48024
rect 42767 46504 42926 48006
rect 42767 46464 42925 46504
rect 42767 46358 42787 46464
rect 42915 46358 42925 46464
rect 42767 46342 42925 46358
rect 42517 39654 42536 39747
rect 42670 39654 42676 39747
rect 42517 39641 42676 39654
rect 42272 38786 42285 38880
rect 42410 38786 42428 38880
rect 42272 38770 42428 38786
rect 42024 38659 42172 38733
rect 42024 38566 42043 38659
rect 42149 38566 42172 38659
rect 42024 38553 42172 38566
rect 41774 38474 42322 38475
rect 41774 38331 42466 38474
rect 41597 38228 42079 38230
rect 41597 38136 42215 38228
rect 42323 38198 42466 38331
rect 41600 38135 42215 38136
rect 41424 38006 41995 38064
rect 41424 37967 41996 38006
rect 41225 37876 41596 37877
rect 41225 37782 41752 37876
rect 41225 37780 41320 37782
rect 41060 37627 41524 37717
rect 40852 37407 41318 37529
rect 40576 37304 40948 37306
rect 40576 37185 41099 37304
rect 40576 37182 40720 37185
rect 25305 36924 25427 36925
rect 24798 36811 24915 36822
rect 24529 36736 24652 36740
rect 24528 36722 24652 36736
rect 24528 36637 24545 36722
rect 24632 36637 24652 36722
rect 24528 36615 24652 36637
rect 23337 36049 23945 36050
rect 23337 36047 24164 36049
rect 23337 36035 24174 36047
rect 23337 35933 23359 36035
rect 23446 35933 24174 36035
rect 23337 35923 24174 35933
rect 23337 35920 23945 35923
rect 24084 34613 24174 35923
rect 24315 36038 24446 36049
rect 24315 35937 24333 36038
rect 24432 35937 24446 36038
rect 24315 34807 24446 35937
rect 24529 34998 24652 36615
rect 24798 36728 24819 36811
rect 24903 36728 24915 36811
rect 24798 35174 24915 36728
rect 25058 36818 25171 36830
rect 25058 36732 25081 36818
rect 25157 36732 25171 36818
rect 25058 36056 25171 36732
rect 25305 36804 29089 36924
rect 25052 35378 25172 36056
rect 25305 35584 25427 36804
rect 25305 35575 27682 35584
rect 25305 35507 27569 35575
rect 27674 35507 27682 35575
rect 25305 35494 27682 35507
rect 40957 35579 41099 37185
rect 41172 36711 41318 37407
rect 41387 36711 41523 37627
rect 41173 36709 41318 36711
rect 40957 35574 41104 35579
rect 40957 35516 40967 35574
rect 41091 35516 41104 35574
rect 40957 35503 41104 35516
rect 25052 35358 27678 35378
rect 25052 35288 27578 35358
rect 27663 35288 27678 35358
rect 25052 35275 27678 35288
rect 41173 35347 41319 36709
rect 41173 35288 41199 35347
rect 41294 35288 41319 35347
rect 25052 35273 25172 35275
rect 41173 35270 41319 35288
rect 24798 35162 27677 35174
rect 24798 35098 27580 35162
rect 27667 35098 27677 35162
rect 24798 35082 27677 35098
rect 24889 35080 27677 35082
rect 41378 35162 41523 36711
rect 41378 35102 41404 35162
rect 41502 35102 41523 35162
rect 41602 35106 41752 37782
rect 41378 35081 41523 35102
rect 24529 34985 27672 34998
rect 24529 34911 27586 34985
rect 27661 34911 27672 34985
rect 24529 34899 27672 34911
rect 41601 34974 41753 35106
rect 41601 34914 41627 34974
rect 41716 34914 41753 34974
rect 41601 34902 41753 34914
rect 41853 34913 41996 37967
rect 42079 35360 42215 38135
rect 42325 37579 42462 38198
rect 42325 37514 42461 37579
rect 42325 37418 42346 37514
rect 42447 37418 42461 37514
rect 42325 37399 42461 37418
rect 42079 34979 42218 35360
rect 41605 34900 41747 34902
rect 24315 34795 27672 34807
rect 24315 34719 27583 34795
rect 27661 34719 27672 34795
rect 24315 34708 27672 34719
rect 41853 34801 42003 34913
rect 41853 34727 41887 34801
rect 41988 34727 42003 34801
rect 41853 34709 42003 34727
rect 24084 34597 27665 34613
rect 24084 34529 27555 34597
rect 27651 34529 27665 34597
rect 24084 34515 27665 34529
rect 42078 34600 42222 34979
rect 42078 34533 42093 34600
rect 42197 34533 42222 34600
rect 42078 34522 42222 34533
rect 24084 34513 24174 34515
<< via2 >>
rect 30617 75732 31137 75814
rect 30623 74613 31157 74702
rect 30621 73500 31171 73581
rect 30628 72383 31170 72462
rect 30617 71259 31166 71338
rect 30676 70136 31145 70213
rect 30624 69019 31155 69093
rect 30638 67894 31156 67980
rect 30806 66776 31147 66850
rect 31039 65664 31172 65740
rect 31030 64535 31149 64620
rect 38138 59699 38227 59817
rect 23300 57689 23364 57750
rect 12384 56577 12507 56678
rect 39731 39652 39884 39742
rect 39722 38791 39865 38870
rect 39723 38574 39855 38659
rect 39712 37406 39888 37513
<< metal3 >>
rect 38108 59817 38248 59847
rect 38108 59699 38138 59817
rect 38227 59699 38248 59817
rect 38108 59673 38248 59699
rect 23287 57750 23376 57760
rect 23287 57689 23300 57750
rect 23364 57689 23376 57750
rect 23287 57680 23376 57689
rect 29842 57144 29994 57145
rect 36810 57144 36990 57805
rect 29842 57041 36990 57144
rect 29940 57040 36990 57041
rect 36810 57034 36990 57040
rect 29842 56839 36444 56945
rect 12367 56678 12524 56691
rect 12367 56577 12384 56678
rect 12507 56577 12524 56678
rect 36288 56582 36442 56839
rect 12367 56561 12524 56577
rect 6017 54601 6142 55976
rect 10996 55657 11096 55979
rect 21386 55829 21464 55887
rect 10996 55656 12247 55657
rect 10996 55564 12504 55656
rect 10652 55391 12467 55476
rect 10656 54601 10795 55391
rect 5997 54468 10795 54601
rect 10656 54466 10795 54468
rect 14965 42584 15574 42597
rect 14965 42488 15459 42584
rect 15560 42488 15574 42584
rect 14965 42476 15574 42488
rect 25307 42582 25917 42599
rect 25307 42495 25327 42582
rect 25412 42495 25917 42582
rect 25307 42481 25917 42495
rect 39700 39742 39901 39756
rect 39700 39652 39731 39742
rect 39884 39652 39901 39742
rect 39700 39639 39901 39652
rect 39690 38870 39894 38893
rect 39690 38791 39722 38870
rect 39865 38791 39894 38870
rect 39690 38773 39894 38791
rect 39690 38659 39888 38675
rect 39690 38574 39723 38659
rect 39855 38574 39888 38659
rect 39690 38553 39888 38574
rect 39700 37513 39919 37529
rect 39700 37406 39712 37513
rect 39888 37406 39919 37513
rect 39700 37394 39919 37406
<< via3 >>
rect 38138 59699 38227 59817
rect 22539 57692 22612 57752
rect 23300 57689 23364 57750
rect 12384 56577 12507 56678
rect 15459 42488 15560 42584
rect 25327 42495 25412 42582
rect 39731 39652 39884 39742
rect 39722 38791 39865 38870
rect 39723 38574 39855 38659
rect 39712 37406 39888 37513
<< metal4 >>
rect 14526 59846 14695 59853
rect 38108 59846 38248 59847
rect 14132 59817 38248 59846
rect 14132 59699 38138 59817
rect 38227 59699 38248 59817
rect 14132 59674 38248 59699
rect 14526 56732 14695 59674
rect 38108 59673 38248 59674
rect 20983 57752 22656 57781
rect 20983 57692 22539 57752
rect 22612 57692 22656 57752
rect 20983 57652 22656 57692
rect 23256 57750 23390 57779
rect 23256 57689 23300 57750
rect 23364 57689 23390 57750
rect 12398 56730 14698 56732
rect 12367 56678 14698 56730
rect 12367 56577 12384 56678
rect 12507 56577 14698 56678
rect 12367 56563 14698 56577
rect 12367 56561 14667 56563
rect 18385 55825 18530 55829
rect 20990 55825 21118 57652
rect 18379 55685 21118 55825
rect 18379 55681 21028 55685
rect 18385 53996 18530 55681
rect 23256 55490 23390 57689
rect 22299 55404 23390 55490
rect 22299 55397 23356 55404
rect 18386 47806 18527 53996
rect 15450 42593 15573 42596
rect 15450 42584 15574 42593
rect 15450 42488 15459 42584
rect 15560 42488 15574 42584
rect 15450 33797 15574 42488
rect 18386 33797 18528 47806
rect 15450 33650 18528 33797
rect 22300 33754 22445 55397
rect 25307 42589 25426 42598
rect 25305 42582 25426 42589
rect 25305 42495 25327 42582
rect 25412 42495 25426 42582
rect 25305 42481 25426 42495
rect 25305 33754 25425 42481
rect 39467 39742 39901 39758
rect 39467 39652 39731 39742
rect 39884 39652 39901 39742
rect 39467 39639 39901 39652
rect 39478 38870 39895 38895
rect 39478 38791 39722 38870
rect 39865 38791 39895 38870
rect 39478 38773 39895 38791
rect 39477 38659 39888 38675
rect 39477 38574 39723 38659
rect 39855 38574 39888 38659
rect 39477 38552 39888 38574
rect 39553 37513 39916 37529
rect 39553 37406 39712 37513
rect 39888 37406 39916 37513
rect 39553 37394 39916 37406
rect 15450 33649 18386 33650
rect 15450 33462 15574 33649
rect 22300 33614 25426 33754
rect 22300 33606 22445 33614
rect 15450 33445 15575 33462
rect 15450 33441 15576 33445
rect 15450 33360 15460 33441
rect 15564 33360 15576 33441
rect 15450 33345 15576 33360
rect 25305 33440 25425 33614
rect 25305 33371 25324 33440
rect 25403 33371 25425 33440
rect 25305 33357 25425 33371
<< via4 >>
rect 15460 33360 15564 33441
rect 25324 33371 25403 33440
<< metal5 >>
rect 15450 33441 15576 33445
rect 15450 33360 15460 33441
rect 15564 33360 15576 33441
rect 15450 33345 15576 33360
rect 25305 33440 25419 33455
rect 25305 33371 25324 33440
rect 25403 33371 25419 33440
rect 25305 33358 25419 33371
use comparator_latched  comparator_latched_0 ~/gf180xd/SAR_ADC_12BIT/layout/comparator
timestamp 1757859342
transform 1 0 6621 0 1 57051
box -2740 -2535 5894 909
use offset_calibration  offset_calibration_0 ~/gf180xd/SAR_ADC_12BIT/layout/offset_calibration
timestamp 1757859342
transform 1 0 30701 0 1 54668
box 0 -144 10208 5371
use premfilier  premfilier_0 ~/gf180xd/SAR_ADC_12BIT/layout/premfilier
timestamp 1757859342
transform -1 0 29516 0 1 58029
box -443 -3480 17080 2350
use state_machine  state_machine_0 ~/gf180xd/SAR_ADC_12BIT/layout/state_machine
timestamp 1757859342
transform 1 0 6794 0 1 62954
box 0 0 24394 27978
use SW_CDAC  SW_CDAC_0
timestamp 1757749174
transform 1 0 675 0 1 364
box -675 -364 20385 52175
use SW_CDAC  SW_CDAC_1
timestamp 1757749174
transform -1 0 40203 0 1 364
box -675 -364 20385 52175
<< labels >>
flabel metal4 15477 33660 15615 33788 0 FreeSans 320 0 0 0 VDAC_P
flabel metal4 25172 33628 25394 33738 0 FreeSans 320 0 0 0 VDAC_N
<< end >>
