magic
tech gf180mcuD
magscale 1 10
timestamp 1757749174
<< metal1 >>
rect 15349 46309 20385 46338
rect 15349 46149 15365 46309
rect 15550 46149 20385 46309
rect 15349 46129 20385 46149
rect -675 36659 -402 36660
rect -675 36622 -351 36659
rect -675 36496 -644 36622
rect -451 36496 -351 36622
rect -675 36470 -351 36496
rect -624 36469 -351 36470
<< via1 >>
rect 15365 46149 15550 46309
rect -644 36496 -451 36622
<< metal2 >>
rect 15110 47237 17570 47238
rect 13914 47169 17570 47237
rect 14941 46309 15580 46334
rect 14941 46302 15365 46309
rect 14938 46149 15365 46302
rect 15550 46149 15580 46309
rect 14938 46133 15580 46149
rect 14938 46076 15146 46133
rect 14144 45925 15148 46076
rect 17454 36737 17570 47169
rect 15134 36735 17570 36737
rect -675 36622 -402 36660
rect -675 36496 -644 36622
rect -451 36496 -402 36622
rect 14310 36621 17570 36735
rect -675 36470 -402 36496
rect -672 35819 -448 36470
rect -671 32475 -448 35819
rect -670 24422 -448 32475
rect -669 16386 -449 24422
rect 15730 17744 16221 17752
rect 15730 17688 16147 17744
rect 16203 17688 16221 17744
rect 15730 17681 16221 17688
rect 15728 17248 16695 17257
rect 15728 17192 16622 17248
rect 16678 17192 16695 17248
rect 15728 17186 16695 17192
rect 15729 16737 16909 16743
rect 15729 16681 16837 16737
rect 16893 16681 16909 16737
rect 15729 16672 16909 16681
rect -669 14131 -448 16386
rect 15726 16235 17143 16240
rect 15726 16179 17065 16235
rect 17121 16179 17143 16235
rect 15726 16169 17143 16179
rect 15726 15742 16450 15749
rect 15726 15686 16372 15742
rect 16428 15686 16450 15742
rect 15726 15678 16450 15686
rect 15726 15244 15979 15252
rect 15726 15188 15902 15244
rect 15958 15188 15979 15244
rect 15726 15181 15979 15188
rect -668 10251 -448 14131
rect 15728 13734 17398 13742
rect 15728 13678 17320 13734
rect 17376 13678 17398 13734
rect 15728 13671 17398 13678
rect 15705 12747 17655 12754
rect 15705 12691 17577 12747
rect 17633 12691 17655 12747
rect 15705 12683 17655 12691
rect 15726 11238 17876 11244
rect 15726 11182 17801 11238
rect 17857 11182 17876 11238
rect 15726 11173 17876 11182
rect -671 5971 -448 10251
rect 15712 8759 18150 8767
rect 15712 8703 18069 8759
rect 18125 8703 18150 8759
rect 15712 8696 18150 8703
rect -671 -144 -451 5971
rect 15727 5768 18395 5775
rect 15727 5712 18317 5768
rect 18373 5712 18395 5768
rect 15727 5704 18395 5712
rect -674 -145 9741 -144
rect -674 -364 20385 -145
<< via2 >>
rect 16147 17688 16203 17744
rect 16622 17192 16678 17248
rect 16837 16681 16893 16737
rect 17065 16179 17121 16235
rect 16372 15686 16428 15742
rect 15902 15188 15958 15244
rect 15651 14178 15707 14234
rect 17320 13678 17376 13734
rect 17577 12691 17633 12747
rect 17801 11182 17857 11238
rect 18069 8703 18125 8759
rect 18317 5712 18373 5768
<< metal3 >>
rect 14352 43263 18395 43391
rect 14338 43053 18150 43181
rect 14348 42800 17876 42931
rect 14344 42555 17655 42681
rect 14342 42304 17398 42430
rect 14726 35125 17143 35217
rect 14717 34910 16909 35016
rect 14718 34722 16695 34818
rect 14713 34537 16450 34634
rect 14707 34345 16221 34444
rect 14702 34151 15979 34249
rect 14700 33957 15729 34055
rect 15631 14234 15729 33957
rect 15881 15244 15979 34151
rect 16123 17744 16221 34345
rect 16123 17688 16147 17744
rect 16203 17688 16221 17744
rect 16123 17681 16221 17688
rect 16352 15742 16450 34537
rect 16597 17248 16695 34722
rect 16597 17192 16622 17248
rect 16678 17192 16695 17248
rect 16597 17186 16695 17192
rect 16811 16737 16909 34910
rect 16811 16681 16837 16737
rect 16893 16681 16909 16737
rect 16811 16672 16909 16681
rect 17045 16235 17143 35125
rect 17045 16179 17065 16235
rect 17121 16179 17143 16235
rect 17045 16169 17143 16179
rect 16352 15686 16372 15742
rect 16428 15686 16450 15742
rect 16352 15678 16450 15686
rect 15881 15188 15902 15244
rect 15958 15188 15979 15244
rect 15881 15181 15979 15188
rect 15631 14178 15651 14234
rect 15707 14178 15729 14234
rect 15631 14172 15729 14178
rect 17300 13734 17398 42304
rect 17300 13678 17320 13734
rect 17376 13678 17398 13734
rect 17300 13671 17398 13678
rect 17557 12747 17655 42555
rect 17557 12691 17577 12747
rect 17633 12691 17655 12747
rect 17557 12683 17655 12691
rect 17778 11238 17876 42800
rect 17778 11182 17801 11238
rect 17857 11182 17876 11238
rect 17778 11173 17876 11182
rect 18052 8759 18150 43053
rect 18052 8703 18069 8759
rect 18125 8703 18150 8759
rect 18052 8696 18150 8703
rect 18297 5768 18395 43263
rect 18297 5712 18317 5768
rect 18373 5712 18395 5768
rect 18297 5704 18395 5712
use bootstrap_layout  bootstrap_layout_0 ~/gf180xd/SAR_ADC_12BIT/layout/bootstraped
timestamp 1757654639
transform 1 0 -439 0 1 41503
box 1597 5140 17738 10672
use CADC_12bit  CADC_12bit_0 ~/gf180xd/SAR_ADC_12BIT/layout/CDAC
timestamp 1757690107
transform 1 0 9 0 1 32462
box 0 -32447 15721 661
use switches_full  switches_full_1 ~/gf180xd/SAR_ADC_12BIT/layout/swiyches
timestamp 1757728064
transform 1 0 244 0 1 35274
box -649 -1317 16970 11150
<< end >>
