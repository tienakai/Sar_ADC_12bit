magic
tech gf180mcuD
magscale 1 10
timestamp 1757325446
<< pwell >>
rect 399 2518 3156 2595
rect 399 2360 3158 2518
rect 399 2274 3156 2360
rect 400 2190 3156 2274
rect 398 523 3156 2190
rect 398 498 3157 523
rect 400 458 3157 498
rect 400 388 3158 458
rect 399 249 3158 388
<< psubdiff >>
rect 401 415 3156 456
rect 401 353 531 415
rect 1382 410 3156 415
rect 1382 353 2079 410
rect 401 348 2079 353
rect 2930 348 3156 410
rect 401 319 3156 348
<< psubdiffcont >>
rect 531 353 1382 415
rect 2079 348 2930 410
<< polysilicon >>
rect 588 2210 3044 2246
<< metal1 >>
rect 498 2152 574 2164
rect 498 2100 510 2152
rect 562 2100 574 2152
rect 498 2096 574 2100
rect 818 2152 894 2164
rect 818 2100 830 2152
rect 882 2100 894 2152
rect 818 2096 894 2100
rect 1138 2152 1214 2164
rect 1138 2100 1150 2152
rect 1202 2100 1214 2152
rect 1138 2096 1214 2100
rect 1458 2152 1534 2164
rect 1458 2100 1470 2152
rect 1522 2100 1534 2152
rect 1458 2096 1534 2100
rect 1778 2152 1854 2164
rect 1778 2100 1790 2152
rect 1842 2100 1854 2152
rect 1778 2096 1854 2100
rect 2098 2152 2174 2164
rect 2098 2100 2110 2152
rect 2162 2100 2174 2152
rect 2098 2096 2174 2100
rect 2418 2152 2494 2164
rect 2418 2100 2430 2152
rect 2482 2100 2494 2152
rect 2418 2096 2494 2100
rect 2738 2152 2814 2164
rect 2738 2100 2750 2152
rect 2802 2100 2814 2152
rect 2738 2096 2814 2100
rect 3058 2152 3134 2164
rect 3058 2100 3070 2152
rect 3122 2100 3134 2152
rect 3058 2096 3134 2100
rect 658 632 734 636
rect 658 580 670 632
rect 722 580 734 632
rect 658 568 734 580
rect 978 632 1054 636
rect 978 580 990 632
rect 1042 580 1054 632
rect 978 568 1054 580
rect 1298 632 1374 636
rect 1298 580 1310 632
rect 1362 580 1374 632
rect 1298 568 1374 580
rect 1618 632 1694 636
rect 1618 580 1630 632
rect 1682 580 1694 632
rect 1618 568 1694 580
rect 1938 632 2014 636
rect 1938 580 1950 632
rect 2002 580 2014 632
rect 1938 568 2014 580
rect 2258 632 2334 636
rect 2258 580 2270 632
rect 2322 580 2334 632
rect 2258 568 2334 580
rect 2578 632 2654 636
rect 2578 580 2590 632
rect 2642 580 2654 632
rect 2578 568 2654 580
rect 2898 632 2974 636
rect 2898 580 2910 632
rect 2962 580 2974 632
rect 2898 568 2974 580
rect 411 415 3151 449
rect 411 353 531 415
rect 1382 410 3151 415
rect 1382 353 2079 410
rect 411 348 2079 353
rect 2930 348 3151 410
rect 411 328 3151 348
<< via1 >>
rect 510 2100 562 2152
rect 830 2100 882 2152
rect 1150 2100 1202 2152
rect 1470 2100 1522 2152
rect 1790 2100 1842 2152
rect 2110 2100 2162 2152
rect 2430 2100 2482 2152
rect 2750 2100 2802 2152
rect 3070 2100 3122 2152
rect 670 580 722 632
rect 990 580 1042 632
rect 1310 580 1362 632
rect 1630 580 1682 632
rect 1950 580 2002 632
rect 2270 580 2322 632
rect 2590 580 2642 632
rect 2910 580 2962 632
<< metal2 >>
rect 498 2152 3134 2164
rect 498 2100 510 2152
rect 562 2100 830 2152
rect 882 2100 1150 2152
rect 1202 2100 1470 2152
rect 1522 2100 1790 2152
rect 1842 2100 2110 2152
rect 2162 2100 2430 2152
rect 2482 2100 2750 2152
rect 2802 2100 3070 2152
rect 3122 2100 3134 2152
rect 498 2096 3134 2100
rect 658 632 2974 636
rect 658 580 670 632
rect 722 580 990 632
rect 1042 580 1310 632
rect 1362 580 1630 632
rect 1682 580 1950 632
rect 2002 580 2270 632
rect 2322 580 2590 632
rect 2642 580 2910 632
rect 2962 580 2974 632
rect 658 568 2974 580
use nfet_03v3_NRY3LQ  nfet_03v3_NRY3LQ_0
timestamp 1757220328
transform 1 0 1896 0 1 1366
box -140 -868 140 868
use nfet_03v3_NRY3LQ  nfet_03v3_NRY3LQ_1
timestamp 1757220328
transform 1 0 2056 0 1 1366
box -140 -868 140 868
use nfet_03v3_NRY3LQ  nfet_03v3_NRY3LQ_2
timestamp 1757220328
transform 1 0 2216 0 1 1366
box -140 -868 140 868
use nfet_03v3_NRY3LQ  nfet_03v3_NRY3LQ_3
timestamp 1757220328
transform 1 0 2376 0 1 1366
box -140 -868 140 868
use nfet_03v3_NRY3LQ  nfet_03v3_NRY3LQ_4
timestamp 1757220328
transform 1 0 2536 0 1 1366
box -140 -868 140 868
use nfet_03v3_NRY3LQ  nfet_03v3_NRY3LQ_5
timestamp 1757220328
transform 1 0 1096 0 1 1366
box -140 -868 140 868
use nfet_03v3_NRY3LQ  nfet_03v3_NRY3LQ_6
timestamp 1757220328
transform 1 0 2856 0 1 1366
box -140 -868 140 868
use nfet_03v3_NRY3LQ  nfet_03v3_NRY3LQ_7
timestamp 1757220328
transform 1 0 2696 0 1 1366
box -140 -868 140 868
use nfet_03v3_NRY3LQ  nfet_03v3_NRY3LQ_8
timestamp 1757220328
transform 1 0 1256 0 1 1366
box -140 -868 140 868
use nfet_03v3_NRY3LQ  nfet_03v3_NRY3LQ_9
timestamp 1757220328
transform 1 0 1416 0 1 1366
box -140 -868 140 868
use nfet_03v3_NRY3LQ  nfet_03v3_NRY3LQ_10
timestamp 1757220328
transform 1 0 1576 0 1 1366
box -140 -868 140 868
use nfet_03v3_NRY3LQ  nfet_03v3_NRY3LQ_11
timestamp 1757220328
transform 1 0 1736 0 1 1366
box -140 -868 140 868
use nfet_03v3_NRY3LQ  nfet_03v3_NRY3LQ_12
timestamp 1757220328
transform 1 0 936 0 1 1366
box -140 -868 140 868
use nfet_03v3_NRY3LQ  nfet_03v3_NRY3LQ_13
timestamp 1757220328
transform 1 0 776 0 1 1366
box -140 -868 140 868
use nfet_03v3_NRY3LQ  nfet_03v3_NRY3LQ_14
timestamp 1757220328
transform 1 0 616 0 1 1366
box -140 -868 140 868
use nfet_03v3_NRY3LQ  nfet_03v3_NRY3LQ_15
timestamp 1757220328
transform 1 0 3016 0 1 1366
box -140 -868 140 868
<< labels >>
flabel metal2 658 568 2974 636 1 FreeSans 800 0 0 0 Cbtm
port 3 n
flabel polysilicon 588 2210 3044 2246 1 FreeSans 800 0 0 0 EN_VCM
port 2 n
flabel metal1 1290 329 2391 445 0 FreeSans 480 0 0 0 VSS
port 4 nsew
flabel metal2 498 2096 3134 2164 1 FreeSans 800 0 0 0 VCM
port 1 n
<< end >>
