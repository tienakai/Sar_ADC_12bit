magic
tech gf180mcuD
magscale 1 10
timestamp 1757859342
<< nwell >>
rect -204 2272 -32 2273
rect -204 2161 4744 2272
rect 8570 2180 9160 2270
rect -204 2016 4859 2161
rect 8316 2074 8576 2166
rect -204 1961 4744 2016
rect -204 141 45 1961
rect 261 1920 4333 1961
rect 100 1829 156 1840
rect 100 270 170 1829
rect 4527 1509 4583 1961
rect 8600 1417 9160 2180
rect 8541 1410 9160 1417
rect 6717 1140 6764 1210
rect 8303 800 8447 801
rect 8303 711 8491 800
rect 1312 676 1386 698
rect 1999 676 2069 691
rect 2675 676 2758 697
rect 3366 676 3441 696
rect 8541 676 8602 1410
rect 1312 620 3662 676
rect 1312 606 1386 620
rect 1661 602 1727 608
rect 1999 606 2069 620
rect 2675 589 2758 620
rect 3366 601 3441 620
rect 3904 586 4615 649
rect 5244 548 5629 638
rect 8260 478 8340 515
rect 100 245 156 270
rect 263 141 4335 156
rect 4538 141 4639 152
rect -204 -104 4735 141
rect -204 -194 419 -104
rect 1646 -116 2667 -104
rect 1620 -493 1821 -434
rect 4834 -555 4932 -59
rect 8259 -617 8340 478
rect 6830 -680 7963 -617
rect 8259 -669 8341 -617
rect 8260 -682 8341 -669
rect 8410 -769 8491 521
rect 8410 -850 8492 -769
rect 12250 -1779 12449 -1778
rect 12250 -2884 14523 -1779
rect 12250 -2888 14519 -2884
rect 13368 -2891 14519 -2888
rect 13368 -2893 14334 -2891
<< pwell >>
rect 10608 1467 12156 1600
rect 8664 1291 9385 1305
rect -279 -1946 460 -866
rect 2462 -1937 4393 -846
rect 8664 -1270 9597 1291
rect 11566 -739 11749 -579
rect 14154 -979 14459 -912
rect 9679 -1080 9684 -1024
rect 8664 -1679 9534 -1270
rect 3570 -1946 3670 -1937
rect -279 -2490 4397 -1946
rect -290 -2563 4397 -2490
rect 8661 -2185 9534 -1679
rect 10490 -1915 12012 -1880
rect 8661 -2511 10287 -2185
rect 10490 -2196 12013 -1915
rect -290 -2900 4390 -2563
rect -290 -3247 4400 -2900
rect 8643 -2935 10287 -2511
rect 10492 -2691 12013 -2196
rect 10492 -2747 11848 -2691
rect 11852 -2707 12013 -2691
rect 11851 -2747 12013 -2707
rect 8643 -2936 9427 -2935
rect 9477 -2939 10064 -2935
rect 10126 -2936 10210 -2935
rect 10492 -2974 12013 -2747
rect 14567 -2382 16520 -1943
rect 16587 -2382 16808 -1943
rect 14567 -3130 16808 -2382
rect -290 -3280 4390 -3247
<< ndiff >>
rect 2724 -1610 2726 -1210
rect 3884 -1400 3960 -1287
rect 9753 -2556 9831 -2456
rect 15805 -2658 15864 -2387
rect 15805 -2722 15868 -2658
rect 15805 -2758 15864 -2722
<< pdiff >>
rect 100 1829 156 1840
rect 100 270 170 1829
rect 100 245 156 270
rect 12489 -2533 12541 -2449
rect 12811 -2515 12863 -2463
rect 12855 -2528 12864 -2523
<< psubdiff >>
rect 8684 1287 8789 1289
rect 9262 1287 9369 1288
rect 8684 1273 9369 1287
rect 8684 1213 8804 1273
rect 9249 1213 9369 1273
rect 8684 1198 9369 1213
rect 8684 745 8789 1198
rect 9262 1128 9369 1198
rect 9262 746 9280 1128
rect 8678 637 8789 745
rect 9260 708 9280 746
rect 9355 746 9369 1128
rect 9355 708 9371 746
rect 9260 637 9371 708
rect 8678 619 9371 637
rect 8678 540 8799 619
rect 9247 540 9371 619
rect 8678 520 9371 540
rect 8680 341 8789 520
rect 2543 -904 4336 -867
rect 2543 -976 2864 -904
rect 4171 -976 4336 -904
rect 2543 -1003 4336 -976
rect -197 -1067 415 -1042
rect -197 -1217 -63 -1067
rect 307 -1217 415 -1067
rect -197 -1249 415 -1217
rect 2543 -1773 2668 -1003
rect 4197 -1771 4330 -1003
rect 2543 -1774 2670 -1773
rect 2543 -1775 2681 -1774
rect 4175 -1775 4330 -1771
rect 2543 -1813 4330 -1775
rect 2543 -1885 2798 -1813
rect 4105 -1885 4330 -1813
rect 2543 -1906 4330 -1885
rect 2593 -1908 4330 -1906
rect 8680 -1527 8699 341
rect 8773 -1527 8789 341
rect 9261 341 9370 520
rect 9261 -1522 9279 341
rect 8680 -1611 8789 -1527
rect 9259 -1527 9279 -1522
rect 9353 -1527 9370 341
rect 9259 -1534 9370 -1527
rect 9259 -1610 9368 -1534
rect 9236 -1611 9370 -1610
rect 8680 -1630 9370 -1611
rect 8680 -1696 8784 -1630
rect 9254 -1696 9370 -1630
rect 8680 -1710 9370 -1696
rect 8680 -2501 8808 -1710
rect 9236 -1711 9370 -1710
rect 9261 -1948 9370 -1870
rect 11892 -1926 11985 -1924
rect 10563 -1928 10955 -1927
rect 11820 -1928 11985 -1926
rect 10563 -1946 11985 -1928
rect 9261 -2046 9368 -1948
rect 10563 -1975 10775 -1946
rect 10562 -2000 10775 -1975
rect 11847 -2000 11985 -1946
rect 10562 -2015 11985 -2000
rect 9268 -2235 9368 -2046
rect 10560 -2020 11985 -2015
rect 10560 -2021 11827 -2020
rect 10560 -2077 10660 -2021
rect 9268 -2249 10211 -2235
rect 9268 -2301 9531 -2249
rect 10119 -2301 10211 -2249
rect 9268 -2316 10211 -2301
rect 8680 -2920 8811 -2501
rect 9268 -2839 9468 -2316
rect 9268 -2840 10060 -2839
rect 10126 -2840 10210 -2316
rect 9268 -2854 10210 -2840
rect 10562 -2839 10658 -2077
rect 11890 -2839 11985 -2020
rect 10562 -2846 11985 -2839
rect 9268 -2878 9533 -2854
rect 9384 -2902 9533 -2878
rect 10038 -2902 10210 -2854
rect 9384 -2919 10210 -2902
rect 9384 -2920 9521 -2919
rect 10058 -2935 10210 -2919
rect 10126 -2936 10210 -2935
rect 10560 -2858 11985 -2846
rect 14627 -2085 16520 -2057
rect 14627 -2140 14914 -2085
rect 15486 -2088 16520 -2085
rect 15486 -2140 15641 -2088
rect 14627 -2143 15641 -2140
rect 16213 -2143 16520 -2088
rect 14627 -2178 16520 -2143
rect 16587 -2156 16737 -2057
rect 16587 -2178 16738 -2156
rect 10560 -2912 10764 -2858
rect 11836 -2912 11985 -2858
rect 14628 -2256 14740 -2178
rect 14628 -2828 14663 -2256
rect 14718 -2828 14740 -2256
rect 10560 -2939 11985 -2912
rect 11816 -2940 11985 -2939
rect 14628 -2962 14740 -2828
rect 15598 -2253 15712 -2178
rect 15598 -2825 15625 -2253
rect 15680 -2825 15712 -2253
rect 16618 -2197 16738 -2178
rect 15598 -2957 15712 -2825
rect 16618 -2769 16645 -2197
rect 16700 -2769 16738 -2197
rect 16618 -2957 16738 -2769
rect 15598 -2962 16738 -2957
rect 14628 -2978 16738 -2962
rect 14628 -2985 16039 -2978
rect 14628 -3040 14843 -2985
rect 15415 -3033 16039 -2985
rect 16611 -3033 16738 -2978
rect 15415 -3040 16738 -3033
rect 14628 -3069 16738 -3040
rect 14816 -3074 16738 -3069
rect 15700 -3075 16738 -3074
rect 15700 -3077 16619 -3075
<< nsubdiff >>
rect -41 2160 4859 2161
rect -114 2071 4859 2160
rect 8316 2074 8576 2166
rect -114 2070 36 2071
rect -114 2005 -12 2070
rect 4538 2016 4859 2071
rect -114 218 -97 2005
rect -30 218 -12 2005
rect -114 85 -12 218
rect -114 65 -11 85
rect -112 30 -11 65
rect 4538 30 4639 152
rect -112 6 4639 30
rect -112 -61 4637 6
rect 1646 -116 2667 -61
rect 12280 -1823 14390 -1809
rect 12280 -1907 13043 -1823
rect 13641 -1907 14390 -1823
rect 12280 -1931 14390 -1907
rect 12281 -2032 12400 -1931
rect 12281 -2630 12297 -2032
rect 12381 -2630 12400 -2032
rect 13249 -2009 13368 -1931
rect 14279 -1961 14390 -1931
rect 14279 -1966 14391 -1961
rect 13249 -2103 13371 -2009
rect 12281 -2750 12400 -2630
rect 13249 -2701 13269 -2103
rect 13353 -2701 13371 -2103
rect 13249 -2749 13371 -2701
rect 14280 -2115 14391 -1966
rect 14280 -2713 14294 -2115
rect 14378 -2713 14391 -2115
rect 14280 -2749 14391 -2713
rect 13249 -2750 14391 -2749
rect 12281 -2763 14391 -2750
rect 12281 -2847 13008 -2763
rect 13606 -2847 14391 -2763
rect 12281 -2858 14391 -2847
rect 12400 -2860 14391 -2858
rect 13248 -2861 13370 -2860
rect 14249 -2861 14313 -2860
<< psubdiffcont >>
rect 8804 1213 9249 1273
rect 9280 708 9355 1128
rect 8799 540 9247 619
rect 2864 -976 4171 -904
rect -63 -1217 307 -1067
rect 2798 -1885 4105 -1813
rect 8699 -1527 8773 341
rect 9279 -1527 9353 341
rect 8784 -1696 9254 -1630
rect 10775 -2000 11847 -1946
rect 9531 -2301 10119 -2249
rect 9533 -2902 10038 -2854
rect 14914 -2140 15486 -2085
rect 15641 -2143 16213 -2088
rect 10764 -2912 11836 -2858
rect 14663 -2828 14718 -2256
rect 15625 -2825 15680 -2253
rect 16645 -2769 16700 -2197
rect 14843 -3040 15415 -2985
rect 16039 -3033 16611 -2978
<< nsubdiffcont >>
rect -97 218 -30 2005
rect 13043 -1907 13641 -1823
rect 12297 -2630 12381 -2032
rect 13269 -2701 13353 -2103
rect 14294 -2713 14378 -2115
rect 13008 -2847 13606 -2763
<< polysilicon >>
rect 2791 -1164 2889 -1081
<< metal1 >>
rect -200 2271 9156 2272
rect -202 2270 9156 2271
rect -202 2251 9157 2270
rect -202 2179 -53 2251
rect 8838 2179 9157 2251
rect -202 2178 9157 2179
rect -202 -43 -186 2178
rect -133 2160 9157 2178
rect 9437 2268 14757 2270
rect 9437 2255 14812 2268
rect 9437 2188 9517 2255
rect 14608 2188 14812 2255
rect 9437 2161 14812 2188
rect -133 2071 4859 2160
rect 8316 2074 8576 2160
rect 14709 2105 14812 2161
rect -133 2070 36 2071
rect -133 2005 -12 2070
rect 4538 2016 4859 2071
rect -133 218 -97 2005
rect -30 218 -12 2005
rect 261 1971 4377 1986
rect 261 1920 4293 1971
rect 4282 1911 4293 1920
rect 4368 1911 4377 1971
rect 4282 1876 4377 1911
rect 8739 1874 8790 1951
rect 8739 1862 8796 1874
rect 8903 1865 8953 1950
rect 100 1817 170 1829
rect 100 283 111 1817
rect 163 283 170 1817
rect 100 270 170 283
rect 289 1810 359 1829
rect 289 286 297 1810
rect 355 286 359 1810
rect 289 270 359 286
rect 437 1811 507 1829
rect 437 287 442 1811
rect 500 287 507 1811
rect 437 270 507 287
rect 635 1810 705 1829
rect 635 286 642 1810
rect 700 286 705 1810
rect 635 270 705 286
rect 775 1810 845 1829
rect 775 286 783 1810
rect 841 286 845 1810
rect 775 270 845 286
rect 974 1809 1044 1829
rect 974 285 980 1809
rect 1038 285 1044 1809
rect 974 270 1044 285
rect 1118 1808 1188 1829
rect 1118 284 1124 1808
rect 1182 284 1188 1808
rect 1118 270 1188 284
rect 1315 1808 1385 1829
rect 1315 284 1323 1808
rect 1381 284 1385 1808
rect 1315 270 1385 284
rect 1460 1809 1530 1829
rect 1460 285 1467 1809
rect 1525 285 1530 1809
rect 1460 270 1530 285
rect 1659 1810 1729 1829
rect 1659 286 1667 1810
rect 1725 286 1729 1810
rect 1659 270 1729 286
rect 1800 1810 1870 1829
rect 1800 286 1806 1810
rect 1864 286 1870 1810
rect 1800 270 1870 286
rect 2000 1808 2070 1829
rect 2000 284 2008 1808
rect 2066 284 2070 1808
rect 2000 270 2070 284
rect 2144 1808 2214 1829
rect 2144 284 2153 1808
rect 2211 284 2214 1808
rect 2144 270 2214 284
rect 2343 1809 2413 1829
rect 2343 285 2351 1809
rect 2409 285 2413 1809
rect 2343 270 2413 285
rect 2485 1810 2555 1829
rect 2485 286 2490 1810
rect 2548 286 2555 1810
rect 2485 270 2555 286
rect 2686 1810 2756 1828
rect 2686 286 2691 1810
rect 2749 286 2756 1810
rect 2686 269 2756 286
rect 2832 1807 2902 1829
rect 2832 283 2838 1807
rect 2896 283 2902 1807
rect 2832 270 2902 283
rect 3030 1806 3100 1829
rect 3030 282 3036 1806
rect 3094 282 3100 1806
rect 3030 270 3100 282
rect 3171 1806 3241 1828
rect 3171 282 3179 1806
rect 3237 282 3241 1806
rect 3171 269 3241 282
rect 3372 1807 3442 1828
rect 3372 283 3379 1807
rect 3437 283 3442 1807
rect 3372 269 3442 283
rect 3511 1810 3581 1829
rect 3511 286 3519 1810
rect 3577 286 3581 1810
rect 3511 270 3581 286
rect 3712 1811 3782 1829
rect 3712 287 3719 1811
rect 3777 287 3782 1811
rect 3712 270 3782 287
rect 3853 1812 3923 1829
rect 3853 288 3858 1812
rect 3916 288 3923 1812
rect 3853 270 3923 288
rect 4055 1811 4125 1829
rect 4055 287 4062 1811
rect 4120 287 4125 1811
rect 4055 270 4125 287
rect 4195 1811 4265 1829
rect 4195 287 4201 1811
rect 4259 287 4265 1811
rect 4195 270 4265 287
rect 4395 1809 4465 1829
rect 4395 285 4404 1809
rect 4462 285 4465 1809
rect 8739 1806 8741 1862
rect 8793 1806 8796 1862
rect 8952 1810 8953 1865
rect 8739 1793 8796 1806
rect 8739 1773 8790 1793
rect 8903 1770 8953 1810
rect 9678 1941 9748 1966
rect 9678 1790 9691 1941
rect 9743 1790 9748 1941
rect 9678 1768 9748 1790
rect 14429 1950 14498 1965
rect 14429 1788 14440 1950
rect 14497 1788 14498 1950
rect 14429 1768 14498 1788
rect 8787 1689 8891 1701
rect 8787 1626 8800 1689
rect 8883 1626 8891 1689
rect 8787 1616 8891 1626
rect 9679 1657 9748 1685
rect 9679 1515 9683 1657
rect 9739 1515 9748 1657
rect 9679 1488 9748 1515
rect 14428 1667 14497 1685
rect 14428 1505 14438 1667
rect 14495 1505 14497 1667
rect 14428 1488 14497 1505
rect 9679 1375 9748 1405
rect 8684 1287 8789 1289
rect 9262 1287 9369 1288
rect 8684 1273 9369 1287
rect 8684 1213 8804 1273
rect 9249 1213 9369 1273
rect 8684 1198 9369 1213
rect 9679 1233 9687 1375
rect 9743 1233 9748 1375
rect 9679 1208 9748 1233
rect 14429 1373 14498 1405
rect 14429 1231 14435 1373
rect 14491 1231 14498 1373
rect 14429 1208 14498 1231
rect 8684 879 8789 1198
rect 9262 1128 9369 1198
rect 8964 1104 9071 1119
rect 8964 1031 8981 1104
rect 9056 1031 9071 1104
rect 8964 1025 9071 1031
rect 9070 932 9140 961
rect 8684 770 8934 879
rect 9070 801 9082 932
rect 9134 801 9140 932
rect 8684 745 8789 770
rect 9070 764 9140 801
rect 9262 746 9280 1128
rect 8678 637 8789 745
rect 9260 708 9280 746
rect 9355 746 9369 1128
rect 9678 1088 9747 1125
rect 9678 946 9685 1088
rect 9741 946 9747 1088
rect 9678 928 9747 946
rect 14428 1106 14497 1125
rect 14428 964 14437 1106
rect 14493 964 14497 1106
rect 14428 928 14497 964
rect 9679 810 9748 845
rect 9355 708 9371 746
rect 9260 658 9371 708
rect 9679 668 9689 810
rect 9745 668 9748 810
rect 9260 637 9501 658
rect 9679 648 9748 668
rect 14428 814 14497 844
rect 14428 672 14437 814
rect 14493 672 14497 814
rect 14428 647 14497 672
rect 8678 619 9501 637
rect 8678 540 8799 619
rect 9247 540 9501 619
rect 8678 531 9501 540
rect 8678 520 9371 531
rect 9679 523 9748 565
rect 4395 270 4465 285
rect 8680 341 8789 520
rect -133 85 -12 218
rect 263 98 4335 164
rect -133 30 -11 85
rect 4538 30 4639 152
rect -133 6 4639 30
rect -133 -43 4637 6
rect -202 -60 4637 -43
rect -206 -61 4637 -60
rect -206 -81 518 -61
rect -206 -137 -78 -81
rect 443 -137 518 -81
rect 1646 -116 2667 -61
rect -206 -154 522 -137
rect -203 -194 522 -154
rect -203 -265 -83 -194
rect 297 -265 522 -194
rect -203 -279 522 -265
rect -119 -283 332 -279
rect 1816 -335 1880 -314
rect 2437 -315 2494 -314
rect 2437 -329 2504 -315
rect 176 -373 252 -353
rect 239 -480 252 -373
rect 176 -501 252 -480
rect 1816 -494 1824 -335
rect 1876 -494 1880 -335
rect 2116 -344 2195 -329
rect 2116 -460 2130 -344
rect 2184 -460 2195 -344
rect 2116 -474 2195 -460
rect 1816 -510 1880 -494
rect 2437 -498 2446 -329
rect 2498 -498 2504 -329
rect 2437 -510 2504 -498
rect 1904 -573 2104 -561
rect -61 -599 42 -584
rect -61 -662 -42 -599
rect 26 -662 42 -599
rect 1904 -638 1925 -573
rect 2091 -638 2104 -573
rect 1904 -649 2104 -638
rect 2207 -570 2407 -559
rect 2207 -632 2230 -570
rect 2392 -632 2407 -570
rect 2207 -648 2407 -632
rect -61 -677 42 -662
rect 2543 -904 4336 -867
rect 2543 -976 2864 -904
rect 4171 -976 4336 -904
rect 2543 -1003 4336 -976
rect -197 -1050 415 -1042
rect -197 -1820 -78 -1050
rect 112 -1067 415 -1050
rect 307 -1217 415 -1067
rect -196 -2705 -78 -1820
rect 112 -1819 415 -1217
rect 2543 -1554 2668 -1003
rect 2791 -1093 2889 -1081
rect 2791 -1158 2805 -1093
rect 2875 -1158 2889 -1093
rect 3332 -1148 3379 -1003
rect 2791 -1164 2889 -1158
rect 3884 -1302 3960 -1287
rect 2905 -1394 2955 -1368
rect 2954 -1533 2955 -1394
rect 3884 -1383 3900 -1302
rect 3952 -1383 3960 -1302
rect 3884 -1400 3960 -1383
rect 2905 -1539 2955 -1533
rect 2942 -1547 2954 -1539
rect 2543 -1607 2777 -1554
rect 2543 -1773 2668 -1607
rect 4197 -1771 4330 -1003
rect 2543 -1774 2670 -1773
rect 4175 -1774 4330 -1771
rect 8680 -1527 8699 341
rect 8773 -1245 8789 341
rect 9261 341 9370 520
rect 9679 381 9689 523
rect 9745 381 9748 523
rect 9679 368 9748 381
rect 14428 535 14497 565
rect 14428 393 14437 535
rect 14493 393 14497 535
rect 14428 368 14497 393
rect 9087 -811 9171 -801
rect 9087 -896 9091 -811
rect 9088 -900 9091 -896
rect 9159 -818 9171 -811
rect 9159 -900 9172 -818
rect 9088 -913 9172 -900
rect 8773 -1354 8941 -1245
rect 8773 -1527 8789 -1354
rect 9261 -1522 9279 341
rect 8680 -1611 8789 -1527
rect 9259 -1527 9279 -1522
rect 9353 -1527 9370 341
rect 9679 246 9748 285
rect 9679 104 9686 246
rect 9742 104 9748 246
rect 9679 88 9748 104
rect 14428 257 14497 285
rect 14428 115 14439 257
rect 14495 115 14497 257
rect 14428 88 14497 115
rect 9679 -36 9748 5
rect 9679 -178 9689 -36
rect 9745 -178 9748 -36
rect 9679 -192 9748 -178
rect 14428 -24 14497 4
rect 14428 -166 14439 -24
rect 14495 -166 14497 -24
rect 14428 -193 14497 -166
rect 14709 -59 14734 2105
rect 14793 -59 14812 2105
rect 9679 -318 9748 -275
rect 9679 -460 9686 -318
rect 9742 -460 9748 -318
rect 9679 -472 9748 -460
rect 14428 -301 14497 -275
rect 14428 -443 14438 -301
rect 14494 -443 14497 -301
rect 14428 -472 14497 -443
rect 9679 -594 9748 -555
rect 9679 -736 9688 -594
rect 9744 -736 9748 -594
rect 9679 -752 9748 -736
rect 14429 -587 14498 -555
rect 14429 -729 14438 -587
rect 14494 -729 14498 -587
rect 14429 -752 14498 -729
rect 9679 -865 9748 -835
rect 9679 -1007 9684 -865
rect 9740 -1007 9748 -865
rect 9679 -1032 9748 -1007
rect 14428 -859 14497 -835
rect 14428 -1001 14437 -859
rect 14493 -1001 14497 -859
rect 14428 -1032 14497 -1001
rect 14709 -1060 14812 -59
rect 14709 -1100 16790 -1060
rect 14709 -1240 15810 -1100
rect 16720 -1240 16790 -1100
rect 14709 -1259 16790 -1240
rect 14770 -1260 16790 -1259
rect 9259 -1534 9370 -1527
rect 9259 -1610 9368 -1534
rect 9236 -1611 9370 -1610
rect 8680 -1630 9370 -1611
rect 8680 -1696 8784 -1630
rect 9254 -1696 9370 -1630
rect 8680 -1710 9370 -1696
rect 2536 -1813 4332 -1774
rect 112 -2420 416 -1819
rect 2536 -1885 2798 -1813
rect 4105 -1885 4332 -1813
rect 112 -2563 410 -2420
rect 2536 -2427 4332 -1885
rect 2534 -2518 4332 -2427
rect 8680 -2501 8808 -1710
rect 9236 -1711 9370 -1710
rect 12280 -1823 14390 -1809
rect 9261 -1948 9370 -1870
rect 12280 -1907 13043 -1823
rect 13641 -1907 14390 -1823
rect 12280 -1909 13052 -1907
rect 13579 -1909 14390 -1907
rect 11892 -1926 11985 -1924
rect 10563 -1928 10955 -1927
rect 11820 -1928 11985 -1926
rect 10563 -1946 11985 -1928
rect 12280 -1931 14390 -1909
rect 9261 -2046 9368 -1948
rect 10563 -1975 10775 -1946
rect 10562 -2000 10775 -1975
rect 11847 -2000 11985 -1946
rect 10562 -2015 11985 -2000
rect 9268 -2235 9368 -2046
rect 10560 -2020 11985 -2015
rect 10560 -2021 11827 -2020
rect 10560 -2077 10660 -2021
rect 9268 -2249 10211 -2235
rect 9268 -2301 9531 -2249
rect 10119 -2301 10211 -2249
rect 9268 -2316 10211 -2301
rect 2534 -2563 4331 -2518
rect 112 -2705 407 -2563
rect -196 -2838 407 -2705
rect -199 -2900 410 -2838
rect 2534 -2900 4327 -2563
rect 8680 -2900 8811 -2501
rect 9268 -2839 9468 -2316
rect 9544 -2454 9621 -2439
rect 9544 -2541 9551 -2454
rect 9610 -2541 9621 -2454
rect 9961 -2450 10039 -2436
rect 9544 -2555 9621 -2541
rect 9753 -2463 9831 -2456
rect 9753 -2548 9765 -2463
rect 9818 -2548 9831 -2463
rect 9753 -2556 9831 -2548
rect 9961 -2536 9974 -2450
rect 10030 -2536 10039 -2450
rect 9961 -2556 10039 -2536
rect 9644 -2623 9736 -2614
rect 9644 -2679 9655 -2623
rect 9726 -2679 9736 -2623
rect 9644 -2690 9736 -2679
rect 9848 -2624 9940 -2614
rect 9848 -2677 9863 -2624
rect 9931 -2677 9940 -2624
rect 9848 -2690 9940 -2677
rect 9268 -2840 10060 -2839
rect 10126 -2840 10210 -2316
rect 9268 -2845 10210 -2840
rect 10562 -2565 10658 -2077
rect 11890 -2109 11985 -2020
rect 11754 -2178 11985 -2109
rect 10937 -2249 11031 -2223
rect 10562 -2616 10771 -2565
rect 10937 -2583 10944 -2249
rect 11020 -2583 11031 -2249
rect 10562 -2839 10658 -2616
rect 10937 -2619 11031 -2583
rect 11210 -2619 11329 -2224
rect 11513 -2257 11634 -2222
rect 11513 -2591 11530 -2257
rect 11606 -2591 11634 -2257
rect 11513 -2618 11634 -2591
rect 11805 -2618 11985 -2178
rect 11240 -2839 11296 -2619
rect 11890 -2839 11985 -2618
rect 10562 -2845 11985 -2839
rect 9268 -2846 11985 -2845
rect 12281 -2032 12400 -1931
rect 13249 -2009 13368 -1931
rect 14279 -1961 14390 -1931
rect 14279 -1966 14391 -1961
rect 12281 -2630 12297 -2032
rect 12381 -2630 12400 -2032
rect 13248 -2103 13371 -2009
rect 12628 -2314 12722 -2301
rect 12628 -2381 12646 -2314
rect 12712 -2381 12722 -2314
rect 12628 -2396 12722 -2381
rect 12945 -2318 13039 -2306
rect 12945 -2389 12960 -2318
rect 13028 -2389 13039 -2318
rect 12945 -2400 13039 -2389
rect 12489 -2462 12545 -2449
rect 12809 -2450 12864 -2445
rect 12489 -2514 12490 -2462
rect 12489 -2530 12545 -2514
rect 12808 -2463 12864 -2450
rect 12808 -2515 12811 -2463
rect 12863 -2515 12864 -2463
rect 12808 -2524 12864 -2515
rect 12809 -2526 12864 -2524
rect 12855 -2528 12864 -2526
rect 13129 -2461 13184 -2447
rect 13129 -2513 13130 -2461
rect 13182 -2513 13184 -2461
rect 13129 -2528 13184 -2513
rect 12489 -2533 12541 -2530
rect 12281 -2750 12400 -2630
rect 13248 -2680 13269 -2103
rect 13249 -2701 13269 -2680
rect 13353 -2701 13371 -2103
rect 14280 -2115 14391 -1966
rect 16590 -2057 16790 -1260
rect 13517 -2180 13580 -2164
rect 13517 -2236 13525 -2180
rect 13577 -2236 13580 -2180
rect 13517 -2251 13580 -2236
rect 13840 -2179 13903 -2163
rect 13840 -2235 13842 -2179
rect 13894 -2235 13903 -2179
rect 13840 -2250 13903 -2235
rect 14160 -2180 14223 -2163
rect 14160 -2236 14164 -2180
rect 14216 -2236 14223 -2180
rect 14160 -2250 14223 -2236
rect 13673 -2462 13740 -2450
rect 13673 -2523 13680 -2462
rect 13732 -2523 13740 -2462
rect 13673 -2536 13740 -2523
rect 13984 -2462 14060 -2451
rect 13984 -2520 13998 -2462
rect 14051 -2520 14060 -2462
rect 13984 -2530 14060 -2520
rect 13249 -2749 13371 -2701
rect 14280 -2713 14294 -2115
rect 14378 -2713 14391 -2115
rect 14627 -2085 16520 -2057
rect 14627 -2140 14914 -2085
rect 15486 -2088 16520 -2085
rect 15486 -2140 15641 -2088
rect 14627 -2143 15641 -2140
rect 16213 -2143 16520 -2088
rect 14627 -2178 16520 -2143
rect 16587 -2170 16790 -2057
rect 16587 -2178 16738 -2170
rect 14280 -2749 14391 -2713
rect 13249 -2750 14391 -2749
rect 12281 -2763 14391 -2750
rect 9268 -2854 12108 -2846
rect 9268 -2859 9533 -2854
rect 9254 -2900 9533 -2859
rect -199 -2902 9533 -2900
rect 10038 -2858 12108 -2854
rect 12281 -2847 13008 -2763
rect 13606 -2847 14391 -2763
rect 12281 -2858 14391 -2847
rect 10038 -2902 10764 -2858
rect -199 -2912 10764 -2902
rect 11836 -2912 12108 -2858
rect 12400 -2860 14391 -2858
rect 14628 -2256 14740 -2178
rect 15364 -2242 15458 -2240
rect 15364 -2244 15379 -2242
rect 14628 -2828 14663 -2256
rect 14718 -2828 14740 -2256
rect 15368 -2266 15379 -2244
rect 15445 -2266 15458 -2242
rect 15447 -2301 15458 -2266
rect 15598 -2253 15712 -2178
rect 16618 -2197 16738 -2178
rect 14965 -2524 15046 -2520
rect 15291 -2521 15372 -2520
rect 14965 -2576 14980 -2524
rect 15033 -2576 15046 -2524
rect 14965 -2588 15046 -2576
rect 15287 -2527 15372 -2521
rect 15287 -2580 15302 -2527
rect 15360 -2580 15372 -2527
rect 15287 -2588 15372 -2580
rect 15287 -2589 15368 -2588
rect 13248 -2861 13370 -2860
rect 14249 -2861 14313 -2860
rect -199 -2940 12108 -2912
rect -199 -2980 690 -2940
rect -210 -3140 690 -2980
rect 4260 -2962 12108 -2940
rect 14628 -2962 14740 -2828
rect 15598 -2825 15625 -2253
rect 15680 -2825 15712 -2253
rect 15859 -2245 15965 -2240
rect 15859 -2297 15872 -2245
rect 15949 -2250 15965 -2245
rect 15949 -2297 15957 -2250
rect 15859 -2301 15957 -2297
rect 15852 -2387 15864 -2386
rect 15805 -2658 15864 -2387
rect 15947 -2570 16032 -2482
rect 15947 -2638 15958 -2570
rect 16026 -2638 16032 -2570
rect 15805 -2660 15868 -2658
rect 15805 -2720 15809 -2660
rect 15863 -2720 15868 -2660
rect 15805 -2722 15868 -2720
rect 15805 -2758 15864 -2722
rect 15947 -2768 16032 -2638
rect 16271 -2580 16350 -2479
rect 16271 -2640 16280 -2580
rect 16344 -2640 16350 -2580
rect 16271 -2669 16350 -2640
rect 15947 -2769 16031 -2768
rect 16271 -2771 16351 -2669
rect 16618 -2769 16645 -2197
rect 16700 -2769 16738 -2197
rect 15598 -2957 15712 -2825
rect 16618 -2957 16738 -2769
rect 15598 -2962 16738 -2957
rect 4260 -2978 16738 -2962
rect 4260 -2985 16039 -2978
rect 4260 -3040 14843 -2985
rect 15415 -3033 16039 -2985
rect 16611 -3019 16738 -2978
rect 16611 -3033 16901 -3019
rect 15415 -3040 16901 -3033
rect 4260 -3140 16901 -3040
rect -210 -3187 16901 -3140
rect -210 -3230 16900 -3187
rect -210 -3440 5410 -3230
rect 16400 -3440 16900 -3230
rect -210 -3480 16900 -3440
<< via1 >>
rect -53 2179 8838 2251
rect -186 -43 -133 2178
rect 9517 2188 14608 2255
rect 4293 1911 4368 1971
rect 111 283 163 1817
rect 297 286 355 1810
rect 442 287 500 1811
rect 642 286 700 1810
rect 783 286 841 1810
rect 980 285 1038 1809
rect 1124 284 1182 1808
rect 1323 284 1381 1808
rect 1467 285 1525 1809
rect 1667 286 1725 1810
rect 1806 286 1864 1810
rect 2008 284 2066 1808
rect 2153 284 2211 1808
rect 2351 285 2409 1809
rect 2490 286 2548 1810
rect 2691 286 2749 1810
rect 2838 283 2896 1807
rect 3036 282 3094 1806
rect 3179 282 3237 1806
rect 3379 283 3437 1807
rect 3519 286 3577 1810
rect 3719 287 3777 1811
rect 3858 288 3916 1812
rect 4062 287 4120 1811
rect 4201 287 4259 1811
rect 4404 285 4462 1809
rect 8741 1806 8793 1862
rect 8900 1810 8952 1865
rect 9691 1790 9743 1941
rect 14440 1788 14497 1950
rect 8800 1626 8883 1689
rect 9683 1515 9739 1657
rect 14438 1505 14495 1667
rect 4977 1310 5029 1420
rect 6717 1140 6769 1210
rect 9687 1233 9743 1375
rect 14435 1231 14491 1373
rect 8981 1031 9056 1104
rect 9082 801 9134 932
rect 9685 946 9741 1088
rect 14437 964 14493 1106
rect 9689 668 9745 810
rect 14437 672 14493 814
rect -78 -137 443 -81
rect -83 -265 297 -194
rect 156 -480 239 -373
rect 1824 -494 1876 -335
rect 2130 -460 2184 -344
rect 2446 -498 2498 -329
rect -42 -662 26 -599
rect 1925 -638 2091 -573
rect 2230 -632 2392 -570
rect -78 -1067 112 -1050
rect -78 -1217 -63 -1067
rect -63 -1217 112 -1067
rect -78 -2705 112 -1217
rect 2805 -1158 2875 -1093
rect 3822 -1134 3878 -1082
rect 3981 -1133 4037 -1081
rect 2902 -1533 2954 -1394
rect 3900 -1383 3952 -1302
rect 3235 -1681 3303 -1624
rect 3405 -1680 3473 -1623
rect 9689 381 9745 523
rect 14437 393 14493 535
rect 9091 -900 9159 -811
rect 9686 104 9742 246
rect 14439 115 14495 257
rect 9689 -178 9745 -36
rect 14439 -166 14495 -24
rect 14734 -59 14793 2105
rect 9686 -460 9742 -318
rect 14438 -443 14494 -301
rect 9688 -736 9744 -594
rect 14438 -729 14494 -587
rect 9684 -1007 9740 -865
rect 14437 -1001 14493 -859
rect 15810 -1240 16720 -1100
rect 13052 -1907 13579 -1841
rect 13052 -1909 13579 -1907
rect 9551 -2541 9610 -2454
rect 9765 -2548 9818 -2463
rect 9974 -2536 10030 -2450
rect 9655 -2679 9726 -2623
rect 9863 -2677 9931 -2624
rect 11097 -2158 11162 -2104
rect 10944 -2583 11020 -2249
rect 11530 -2591 11606 -2257
rect 11392 -2729 11450 -2677
rect 12646 -2381 12712 -2314
rect 12960 -2389 13028 -2318
rect 12490 -2514 12545 -2462
rect 12811 -2515 12863 -2463
rect 13130 -2513 13182 -2461
rect 13525 -2236 13577 -2180
rect 13842 -2235 13894 -2179
rect 14164 -2236 14216 -2180
rect 13680 -2523 13732 -2462
rect 13998 -2520 14051 -2462
rect 15379 -2294 15445 -2242
rect 14980 -2576 15033 -2524
rect 15302 -2580 15360 -2527
rect 690 -3140 4260 -2940
rect 15872 -2297 15949 -2245
rect 15958 -2638 16026 -2570
rect 15809 -2720 15863 -2660
rect 16280 -2640 16344 -2580
rect 5410 -3440 16400 -3230
<< metal2 >>
rect -200 2271 9160 2350
rect -202 2251 9160 2271
rect -202 2179 -53 2251
rect 8838 2179 9160 2251
rect -202 2178 9160 2179
rect -202 1580 -186 2178
rect -133 2160 9160 2178
rect 9437 2268 14757 2270
rect 9437 2255 14812 2268
rect 9437 2188 9517 2255
rect 14608 2188 14812 2255
rect 9437 2161 14812 2188
rect -133 1585 -112 2160
rect 4282 1971 4377 1985
rect 4282 1911 4293 1971
rect 4368 1911 4377 1971
rect 4282 1899 4377 1911
rect 100 1817 170 1840
rect 100 1585 111 1817
rect -133 1580 111 1585
rect -202 1481 -196 1580
rect -119 1481 111 1580
rect -202 -43 -186 1481
rect -133 1470 111 1481
rect -133 -43 -112 1470
rect 100 283 111 1470
rect 163 1585 170 1817
rect 290 1810 363 1841
rect 290 1585 297 1810
rect 163 1470 297 1585
rect 163 283 170 1470
rect 100 244 170 283
rect 290 286 297 1470
rect 355 286 363 1810
rect 290 241 363 286
rect 430 1811 503 1841
rect 430 287 442 1811
rect 500 1577 503 1811
rect 502 1481 503 1577
rect 500 287 503 1481
rect 430 241 503 287
rect 634 1810 707 1842
rect 634 286 642 1810
rect 700 286 707 1810
rect 634 242 707 286
rect 775 1810 848 1842
rect 775 1576 783 1810
rect 775 1480 780 1576
rect 775 286 783 1480
rect 841 286 848 1810
rect 775 242 848 286
rect 972 1809 1045 1842
rect 972 285 980 1809
rect 1038 285 1045 1809
rect 972 242 1045 285
rect 1118 1808 1191 1842
rect 1118 1577 1124 1808
rect 1118 1481 1123 1577
rect 1118 284 1124 1481
rect 1182 284 1191 1808
rect 1118 242 1191 284
rect 1313 1808 1386 1842
rect 1313 687 1323 1808
rect 1381 687 1386 1808
rect 1313 625 1320 687
rect 1382 625 1386 687
rect 1313 390 1323 625
rect 1313 309 1318 390
rect 1313 284 1323 309
rect 1381 284 1386 625
rect 1313 242 1386 284
rect 1459 1809 1532 1842
rect 1459 1575 1467 1809
rect 1459 1479 1463 1575
rect 1459 285 1467 1479
rect 1525 285 1532 1809
rect 1459 242 1532 285
rect 1655 1810 1728 1842
rect 1655 390 1667 1810
rect 1655 309 1663 390
rect 1655 286 1667 309
rect 1725 286 1728 1810
rect 1655 242 1728 286
rect 1800 1810 1873 1842
rect 1800 1575 1806 1810
rect 1800 1479 1804 1575
rect 1800 286 1806 1479
rect 1864 286 1873 1810
rect 1800 242 1873 286
rect 1997 1808 2070 1842
rect 1997 390 2008 1808
rect 1997 309 2004 390
rect 1997 284 2008 309
rect 2066 284 2070 1808
rect 1997 242 2070 284
rect 2144 1808 2217 1842
rect 2144 1576 2153 1808
rect 2144 1480 2148 1576
rect 2144 284 2153 1480
rect 2211 284 2217 1808
rect 2144 242 2217 284
rect 2342 1809 2415 1841
rect 2342 285 2351 1809
rect 2409 285 2415 1809
rect 2342 241 2415 285
rect 2483 1810 2556 1842
rect 2483 1575 2490 1810
rect 2483 1479 2489 1575
rect 2483 286 2490 1479
rect 2548 286 2556 1810
rect 2483 242 2556 286
rect 2685 1810 2758 1841
rect 2685 684 2691 1810
rect 2749 684 2758 1810
rect 2685 602 2690 684
rect 2754 602 2758 684
rect 2685 286 2691 602
rect 2749 390 2758 602
rect 2756 309 2758 390
rect 2749 286 2758 309
rect 2685 241 2758 286
rect 2831 1807 2904 1842
rect 2831 1576 2838 1807
rect 2831 1480 2835 1576
rect 2831 283 2838 1480
rect 2896 283 2904 1807
rect 2831 242 2904 283
rect 3030 1806 3101 1840
rect 3030 681 3036 1806
rect 3030 606 3035 681
rect 3030 391 3036 606
rect 3030 310 3033 391
rect 3030 282 3036 310
rect 3094 282 3101 1806
rect 3030 242 3101 282
rect 3171 1806 3242 1840
rect 3171 1576 3179 1806
rect 3171 1480 3174 1576
rect 3171 282 3179 1480
rect 3237 282 3242 1806
rect 3171 242 3242 282
rect 3371 1807 3442 1840
rect 3371 679 3379 1807
rect 3371 613 3378 679
rect 3371 391 3379 613
rect 3371 310 3375 391
rect 3371 283 3379 310
rect 3437 283 3442 1807
rect 3371 242 3442 283
rect 3511 1810 3582 1841
rect 3511 1575 3519 1810
rect 3511 1479 3514 1575
rect 3511 286 3519 1479
rect 3577 286 3582 1810
rect 3511 243 3582 286
rect 3710 1811 3781 1841
rect 3710 548 3719 1811
rect 3777 548 3781 1811
rect 3710 470 3716 548
rect 3779 470 3781 548
rect 3710 287 3719 470
rect 3777 287 3781 470
rect 3710 243 3781 287
rect 3854 1812 3925 1840
rect 3854 1577 3858 1812
rect 3854 1481 3855 1577
rect 3854 288 3858 1481
rect 3916 288 3925 1812
rect 3854 242 3925 288
rect 4055 1811 4126 1840
rect 4055 1032 4062 1811
rect 4055 958 4061 1032
rect 4055 287 4062 958
rect 4120 287 4126 1811
rect 4055 242 4126 287
rect 4196 1811 4267 1841
rect 4196 287 4201 1811
rect 4259 1583 4267 1811
rect 4396 1809 4467 1840
rect 4396 1583 4404 1809
rect 4259 1508 4404 1583
rect 4259 287 4267 1508
rect 4196 243 4267 287
rect 4396 285 4404 1508
rect 4462 1583 4467 1809
rect 4527 1583 4583 2160
rect 8560 1977 8796 1981
rect 8560 1920 8573 1977
rect 8630 1920 8796 1977
rect 8560 1910 8796 1920
rect 8739 1862 8796 1910
rect 8899 1945 8959 2160
rect 14709 2105 14812 2161
rect 8899 1871 8957 1945
rect 8739 1806 8741 1862
rect 8793 1806 8796 1862
rect 8894 1865 8957 1871
rect 8894 1810 8900 1865
rect 8952 1810 8957 1865
rect 8894 1806 8957 1810
rect 8739 1770 8796 1806
rect 8899 1764 8957 1806
rect 9678 1942 9748 1966
rect 9678 1790 9688 1942
rect 9744 1790 9748 1942
rect 9678 1768 9748 1790
rect 14429 1955 14498 1965
rect 14429 1950 14501 1955
rect 14429 1788 14440 1950
rect 14497 1788 14501 1950
rect 14429 1773 14500 1788
rect 4462 1509 4583 1583
rect 8784 1689 8889 1702
rect 8784 1626 8800 1689
rect 8883 1626 8889 1689
rect 14429 1685 14499 1773
rect 4462 1508 4532 1509
rect 4462 285 4467 1508
rect 4947 1420 5033 1437
rect 4947 1419 4977 1420
rect 4947 1309 4962 1419
rect 5029 1310 5033 1420
rect 5022 1309 5033 1310
rect 4947 1293 5033 1309
rect 8784 1382 8889 1626
rect 9679 1657 9748 1685
rect 14428 1672 14499 1685
rect 14428 1667 14497 1672
rect 9679 1515 9683 1657
rect 9739 1611 9748 1657
rect 13055 1640 13278 1657
rect 9739 1604 9969 1611
rect 9739 1532 9970 1604
rect 10041 1589 10161 1604
rect 9739 1515 9748 1532
rect 9679 1488 9748 1515
rect 8784 1381 9382 1382
rect 8784 1298 9384 1381
rect 6703 1210 6771 1225
rect 6703 1140 6710 1210
rect 6770 1140 6771 1210
rect 6703 1122 6771 1140
rect 8596 1118 9066 1121
rect 8595 1104 9066 1118
rect 8595 1031 8981 1104
rect 9056 1031 9066 1104
rect 8595 1020 9066 1031
rect 8406 791 8490 799
rect 8406 726 8422 791
rect 8480 726 8490 791
rect 8260 627 8341 639
rect 8260 564 8274 627
rect 8334 564 8341 627
rect 8260 478 8341 564
rect 8406 521 8490 726
rect 8406 509 8491 521
rect 8259 429 8341 478
rect 4396 242 4467 285
rect -202 -60 -112 -43
rect -206 -81 518 -60
rect -206 -137 -78 -81
rect 443 -137 518 -81
rect -206 -154 522 -137
rect -203 -194 522 -154
rect -203 -265 -83 -194
rect 297 -265 522 -194
rect -203 -279 522 -265
rect -119 -283 332 -279
rect 1816 -335 1880 -314
rect 2437 -315 2494 -314
rect 2437 -329 2504 -315
rect 134 -367 252 -353
rect 483 -367 587 -365
rect 134 -373 587 -367
rect 134 -480 156 -373
rect 239 -479 587 -373
rect 239 -480 252 -479
rect 134 -500 252 -480
rect -61 -599 42 -584
rect -440 -600 -42 -599
rect -440 -659 -43 -600
rect -370 -660 -43 -659
rect -61 -664 -43 -660
rect 26 -664 42 -599
rect -61 -677 42 -664
rect -195 -1050 410 -950
rect -195 -2705 -78 -1050
rect 112 -2563 410 -1050
rect 483 -1831 587 -479
rect 1619 -434 1699 -431
rect 1816 -434 1824 -335
rect 1619 -493 1824 -434
rect 719 -608 824 -598
rect 719 -665 728 -608
rect 813 -665 824 -608
rect 719 -670 824 -665
rect 720 -1240 824 -670
rect 483 -1926 491 -1831
rect 575 -1926 587 -1831
rect 483 -1933 587 -1926
rect 719 -1326 824 -1240
rect 719 -2135 822 -1326
rect 1619 -1751 1699 -493
rect 1816 -494 1824 -493
rect 1876 -494 1880 -335
rect 2116 -344 2195 -329
rect 2116 -460 2130 -344
rect 2186 -460 2195 -344
rect 2116 -474 2195 -460
rect 1816 -510 1880 -494
rect 2437 -498 2446 -329
rect 2498 -370 2504 -329
rect 2498 -371 4583 -370
rect 2498 -471 4596 -371
rect 2498 -498 2504 -471
rect 2437 -510 2504 -498
rect 1904 -573 2104 -561
rect 1904 -638 1925 -573
rect 2091 -638 2104 -573
rect 1904 -649 2104 -638
rect 2207 -570 2407 -559
rect 2207 -632 2230 -570
rect 2392 -632 2407 -570
rect 2207 -648 2407 -632
rect 1926 -904 2037 -649
rect 1926 -973 1940 -904
rect 2020 -973 2037 -904
rect 1926 -992 2037 -973
rect 2252 -1104 2362 -648
rect 2890 -1021 4060 -1020
rect 2252 -1182 2265 -1104
rect 2350 -1182 2362 -1104
rect 2791 -1072 4060 -1021
rect 2791 -1082 3862 -1072
rect 3983 -1081 4060 -1072
rect 2791 -1093 3822 -1082
rect 2791 -1158 2805 -1093
rect 2875 -1100 3822 -1093
rect 2875 -1158 2959 -1100
rect 3795 -1134 3822 -1100
rect 4037 -1133 4060 -1081
rect 3878 -1134 4060 -1133
rect 3795 -1154 4060 -1134
rect 2791 -1164 2959 -1158
rect 2795 -1165 2959 -1164
rect 2875 -1166 2959 -1165
rect 2252 -1194 2362 -1182
rect 2897 -1215 2959 -1166
rect 3534 -1167 3632 -1166
rect 3534 -1169 3633 -1167
rect 2897 -1394 2957 -1215
rect 3534 -1245 3634 -1169
rect 3536 -1248 3634 -1245
rect 2897 -1533 2902 -1394
rect 2954 -1533 2957 -1394
rect 2897 -1615 2957 -1533
rect 3566 -1518 3633 -1248
rect 3884 -1300 3960 -1287
rect 3884 -1383 3897 -1300
rect 3954 -1383 3960 -1300
rect 3884 -1400 3960 -1383
rect 3566 -1599 3905 -1518
rect 3220 -1615 3480 -1611
rect 2897 -1623 3480 -1615
rect 2897 -1624 3405 -1623
rect 2897 -1681 3235 -1624
rect 3303 -1680 3405 -1624
rect 3473 -1680 3480 -1623
rect 3303 -1681 3480 -1680
rect 2897 -1691 3480 -1681
rect 2897 -1693 3270 -1691
rect 3388 -1694 3480 -1691
rect 1619 -1816 1628 -1751
rect 1697 -1816 1699 -1751
rect 1619 -1828 1699 -1816
rect 719 -2200 734 -2135
rect 812 -2200 822 -2135
rect 719 -2210 822 -2200
rect 112 -2705 407 -2563
rect -195 -2838 407 -2705
rect -199 -2900 410 -2838
rect 3570 -2900 3670 -1599
rect 4495 -2468 4596 -471
rect 8259 -617 8340 429
rect 8259 -669 8272 -617
rect 8260 -674 8272 -669
rect 8335 -674 8341 -617
rect 8260 -682 8341 -674
rect 8410 -718 8491 509
rect 8407 -781 8494 -718
rect 8407 -837 8425 -781
rect 8482 -837 8494 -781
rect 8407 -1527 8494 -837
rect 8407 -1604 8419 -1527
rect 8486 -1604 8494 -1527
rect 8407 -1616 8494 -1604
rect 8595 -1934 8708 1020
rect 9070 954 9140 964
rect 9070 898 9077 954
rect 9135 898 9140 954
rect 9070 801 9082 898
rect 9134 801 9140 898
rect 9070 764 9140 801
rect 9079 -811 9171 -801
rect 9079 -900 9091 -811
rect 9159 -900 9171 -811
rect 9079 -913 9171 -900
rect 8595 -2010 8617 -1934
rect 8700 -2010 8708 -1934
rect 8595 -2033 8708 -2010
rect 8952 -2127 9078 -1410
rect 9299 -1534 9384 1298
rect 9679 1375 9748 1405
rect 9679 1233 9687 1375
rect 9743 1233 9748 1375
rect 9679 1224 9748 1233
rect 9678 1208 9748 1224
rect 9678 1088 9747 1208
rect 9527 976 9595 986
rect 9527 920 9535 976
rect 9591 920 9595 976
rect 9678 946 9685 1088
rect 9741 946 9747 1088
rect 9678 928 9747 946
rect 9527 910 9595 920
rect 9860 919 9970 1532
rect 10039 1582 10161 1589
rect 10039 1480 10053 1582
rect 10149 1480 10161 1582
rect 10039 1468 10161 1480
rect 13055 1488 13088 1640
rect 13251 1488 13278 1640
rect 14428 1505 14438 1667
rect 14495 1505 14497 1667
rect 14428 1488 14497 1505
rect 9527 312 9589 910
rect 9679 810 9748 845
rect 9679 668 9689 810
rect 9745 668 9748 810
rect 9679 652 9748 668
rect 9679 648 9749 652
rect 9680 565 9749 648
rect 9679 543 9749 565
rect 9679 523 9748 543
rect 9679 381 9689 523
rect 9745 381 9748 523
rect 9679 368 9748 381
rect 9527 296 9622 312
rect 9527 239 9540 296
rect 9613 239 9622 296
rect 9527 227 9622 239
rect 9679 246 9748 285
rect 9679 104 9686 246
rect 9742 104 9748 246
rect 9679 -36 9748 104
rect 9679 -178 9689 -36
rect 9745 -178 9748 -36
rect 9679 -192 9748 -178
rect 9679 -318 9748 -275
rect 9679 -460 9686 -318
rect 9742 -460 9748 -318
rect 9483 -619 9560 -562
rect 9483 -675 9494 -619
rect 9550 -675 9560 -619
rect 9483 -682 9560 -675
rect 9679 -594 9748 -460
rect 9679 -736 9688 -594
rect 9744 -736 9748 -594
rect 9679 -752 9748 -736
rect 9861 -824 9969 919
rect 9679 -865 9748 -835
rect 9679 -1007 9684 -865
rect 9740 -1007 9748 -865
rect 9861 -887 9868 -824
rect 9959 -887 9969 -824
rect 9861 -900 9969 -887
rect 9679 -1012 9748 -1007
rect 9679 -1079 9750 -1012
rect 9609 -1097 9750 -1079
rect 9609 -1156 9636 -1097
rect 9730 -1156 9750 -1097
rect 9609 -1173 9750 -1156
rect 9680 -1174 9750 -1173
rect 10039 -1309 10121 1468
rect 13055 1465 13278 1488
rect 11566 -607 11749 -579
rect 11566 -703 11605 -607
rect 11719 -703 11749 -607
rect 11566 -739 11749 -703
rect 10426 -1309 10510 -1300
rect 9300 -1782 9384 -1534
rect 9299 -1864 9384 -1782
rect 9296 -1882 9384 -1864
rect 9753 -1320 9833 -1318
rect 10039 -1320 10120 -1309
rect 9753 -1394 10120 -1320
rect 10426 -1373 10436 -1309
rect 10503 -1373 10510 -1309
rect 9753 -1396 10119 -1394
rect 9296 -2046 9383 -1882
rect 9295 -2126 9383 -2046
rect 9241 -2127 9383 -2126
rect 8952 -2138 9383 -2127
rect 8952 -2203 8963 -2138
rect 9069 -2203 9383 -2138
rect 8952 -2209 9383 -2203
rect 8952 -2211 9379 -2209
rect 8952 -2212 9242 -2211
rect 8952 -2213 9078 -2212
rect 9544 -2454 9621 -2439
rect 4494 -2728 4598 -2468
rect 9544 -2541 9551 -2454
rect 9610 -2541 9621 -2454
rect 9544 -2555 9621 -2541
rect 9753 -2463 9833 -1396
rect 10038 -1397 10119 -1396
rect 10109 -1462 10188 -1458
rect 10109 -1521 10120 -1462
rect 10178 -1521 10188 -1462
rect 10109 -1531 10188 -1521
rect 9753 -2548 9765 -2463
rect 9818 -2548 9833 -2463
rect 9753 -2556 9833 -2548
rect 9961 -2450 10039 -2436
rect 9961 -2536 9974 -2450
rect 10030 -2536 10039 -2450
rect 9961 -2556 10039 -2536
rect 10126 -2614 10184 -1531
rect 9644 -2623 9736 -2614
rect 9644 -2679 9655 -2623
rect 9726 -2679 9736 -2623
rect 9644 -2690 9736 -2679
rect 9848 -2624 10184 -2614
rect 9848 -2677 9863 -2624
rect 9931 -2671 10184 -2624
rect 10245 -1612 10319 -1595
rect 10245 -1669 10258 -1612
rect 10314 -1669 10319 -1612
rect 10245 -1682 10319 -1669
rect 9931 -2672 10177 -2671
rect 9931 -2677 9940 -2672
rect 9848 -2690 9940 -2677
rect 9353 -2728 9467 -2723
rect 4494 -2840 9467 -2728
rect 9660 -2776 9725 -2690
rect 10245 -2776 10304 -1682
rect 10426 -2065 10510 -1373
rect 11649 -1619 11725 -739
rect 11649 -1620 12226 -1619
rect 11649 -1711 12233 -1620
rect 11697 -1769 12029 -1768
rect 11697 -1782 12089 -1769
rect 11697 -1854 11705 -1782
rect 11778 -1854 12089 -1782
rect 11697 -1864 12089 -1854
rect 10426 -2094 10511 -2065
rect 10426 -2161 10439 -2094
rect 10503 -2161 10511 -2094
rect 10426 -2172 10511 -2161
rect 11077 -2098 11311 -2087
rect 11077 -2161 11096 -2098
rect 11164 -2161 11311 -2098
rect 11077 -2174 11311 -2161
rect 11077 -2176 11176 -2174
rect 10924 -2249 11045 -2222
rect 10924 -2480 10944 -2249
rect 11020 -2480 11045 -2249
rect 10924 -2591 10942 -2480
rect 11031 -2591 11045 -2480
rect 10924 -2618 11045 -2591
rect 11244 -2666 11309 -2174
rect 11513 -2240 11634 -2222
rect 11513 -2257 11533 -2240
rect 11513 -2591 11530 -2257
rect 11620 -2325 11634 -2240
rect 11606 -2591 11634 -2325
rect 12029 -2460 12089 -1864
rect 12150 -2164 12233 -1711
rect 13084 -1809 13232 1465
rect 14429 1373 14498 1405
rect 13767 1268 13896 1272
rect 14429 1268 14435 1373
rect 13767 1231 14435 1268
rect 14491 1268 14498 1373
rect 14491 1231 14500 1268
rect 13767 1198 14500 1231
rect 13767 -1473 13896 1198
rect 14428 1106 14497 1125
rect 14428 964 14437 1106
rect 14493 964 14497 1106
rect 14428 942 14497 964
rect 14427 928 14497 942
rect 14427 844 14496 928
rect 14427 833 14497 844
rect 14428 814 14497 833
rect 14428 672 14437 814
rect 14493 672 14497 814
rect 14428 647 14497 672
rect 14428 535 14497 565
rect 14428 393 14437 535
rect 14493 393 14497 535
rect 14131 301 14199 302
rect 14076 287 14202 301
rect 14076 200 14097 287
rect 14192 200 14202 287
rect 14076 184 14202 200
rect 14428 257 14497 393
rect 14131 -912 14199 184
rect 14428 115 14439 257
rect 14495 115 14497 257
rect 14428 88 14497 115
rect 14428 -24 14497 4
rect 14709 -10 14734 2105
rect 14428 -166 14439 -24
rect 14495 -166 14497 -24
rect 14428 -301 14497 -166
rect 14428 -443 14438 -301
rect 14494 -443 14497 -301
rect 14428 -472 14497 -443
rect 14670 -59 14734 -10
rect 14793 -59 14812 2105
rect 14670 -430 14810 -59
rect 14429 -587 14498 -555
rect 14429 -729 14438 -587
rect 14494 -695 14498 -587
rect 14670 -600 15730 -430
rect 14494 -707 15039 -695
rect 14494 -729 14955 -707
rect 14429 -752 14955 -729
rect 14491 -753 14955 -752
rect 14941 -777 14955 -753
rect 15027 -753 15039 -707
rect 15027 -777 15037 -753
rect 14941 -790 15037 -777
rect 14428 -859 14497 -835
rect 14428 -912 14437 -859
rect 14131 -979 14437 -912
rect 14131 -1099 14199 -979
rect 14428 -1001 14437 -979
rect 14493 -1001 14497 -859
rect 14428 -1032 14497 -1001
rect 15560 -1050 15730 -600
rect 14131 -1100 14825 -1099
rect 15194 -1100 15411 -1099
rect 15560 -1100 16910 -1050
rect 14131 -1162 15438 -1100
rect 14131 -1163 15201 -1162
rect 13765 -1481 13903 -1473
rect 13765 -1550 13786 -1481
rect 13893 -1550 13903 -1481
rect 13765 -1564 13903 -1550
rect 14447 -1477 14579 -1470
rect 14447 -1549 14471 -1477
rect 14570 -1541 14579 -1477
rect 14570 -1549 14588 -1541
rect 14447 -1560 14588 -1549
rect 12716 -1841 14136 -1809
rect 12716 -1909 13052 -1841
rect 13579 -1909 14136 -1841
rect 12716 -1931 14136 -1909
rect 14309 -2019 14384 -2017
rect 14124 -2023 14384 -2019
rect 12787 -2088 13081 -2025
rect 13104 -2089 14384 -2023
rect 13104 -2090 14137 -2089
rect 13284 -2093 13376 -2090
rect 14043 -2163 14231 -2160
rect 13517 -2164 14231 -2163
rect 12150 -2179 14231 -2164
rect 12150 -2180 13842 -2179
rect 12150 -2236 13525 -2180
rect 13577 -2235 13842 -2180
rect 13894 -2180 14231 -2179
rect 13894 -2235 14164 -2180
rect 13577 -2236 14164 -2235
rect 14216 -2236 14231 -2180
rect 12150 -2249 14231 -2236
rect 13517 -2250 14231 -2249
rect 13517 -2251 14048 -2250
rect 12628 -2314 12723 -2305
rect 12628 -2381 12646 -2314
rect 12712 -2323 12723 -2314
rect 12945 -2318 13039 -2306
rect 12945 -2323 12960 -2318
rect 12712 -2381 12960 -2323
rect 12628 -2389 12960 -2381
rect 13029 -2389 13039 -2318
rect 12628 -2396 13039 -2389
rect 12945 -2400 13039 -2396
rect 13126 -2460 13195 -2447
rect 12029 -2461 13195 -2460
rect 12029 -2462 13130 -2461
rect 12029 -2514 12490 -2462
rect 12545 -2463 13130 -2462
rect 12545 -2514 12811 -2463
rect 12029 -2515 12811 -2514
rect 12863 -2513 13130 -2463
rect 13182 -2513 13195 -2461
rect 12863 -2515 13195 -2513
rect 12029 -2519 13195 -2515
rect 13126 -2528 13195 -2519
rect 13669 -2450 13757 -2448
rect 13669 -2461 14075 -2450
rect 13669 -2462 13998 -2461
rect 13669 -2523 13680 -2462
rect 13732 -2520 13998 -2462
rect 14054 -2520 14075 -2461
rect 13732 -2523 14075 -2520
rect 13669 -2536 14075 -2523
rect 11513 -2618 11634 -2591
rect 14309 -2597 14384 -2089
rect 14489 -2303 14588 -1560
rect 15369 -2219 15438 -1162
rect 15560 -1240 15810 -1100
rect 16720 -1240 16910 -1100
rect 15560 -1260 16910 -1240
rect 15363 -2224 15457 -2219
rect 15363 -2239 15458 -2224
rect 15363 -2240 15858 -2239
rect 15363 -2242 15965 -2240
rect 15363 -2294 15379 -2242
rect 15445 -2245 15965 -2242
rect 15445 -2294 15872 -2245
rect 15363 -2297 15872 -2294
rect 15949 -2297 15965 -2245
rect 15363 -2300 15965 -2297
rect 15363 -2301 15458 -2300
rect 15851 -2301 15965 -2300
rect 14489 -2326 14589 -2303
rect 14489 -2382 14497 -2326
rect 14582 -2382 14589 -2326
rect 14489 -2389 14589 -2382
rect 14490 -2521 14589 -2389
rect 14965 -2521 15046 -2520
rect 15386 -2521 15588 -2519
rect 14490 -2524 15588 -2521
rect 14490 -2576 14980 -2524
rect 15033 -2527 15588 -2524
rect 15033 -2576 15302 -2527
rect 14490 -2580 15302 -2576
rect 15360 -2578 15588 -2527
rect 15360 -2580 15590 -2578
rect 14490 -2581 15590 -2580
rect 14625 -2582 15590 -2581
rect 14625 -2584 15397 -2582
rect 14965 -2588 15046 -2584
rect 13284 -2604 13376 -2602
rect 13982 -2604 14384 -2597
rect 11376 -2666 11465 -2661
rect 11244 -2677 11465 -2666
rect 11244 -2729 11392 -2677
rect 11450 -2729 11465 -2677
rect 11244 -2745 11465 -2729
rect 11376 -2746 11465 -2745
rect 9660 -2835 10362 -2776
rect 10245 -2836 10304 -2835
rect 4589 -2841 9467 -2840
rect -199 -2940 4320 -2900
rect -199 -2980 690 -2940
rect -210 -3140 690 -2980
rect 4260 -2980 4320 -2940
rect 9353 -2970 9467 -2841
rect 11521 -2970 11620 -2618
rect 12616 -2673 12910 -2610
rect 12952 -2670 14384 -2604
rect 12952 -2671 13985 -2670
rect 15527 -2828 15590 -2582
rect 15805 -2658 15864 -2387
rect 15947 -2570 16035 -2559
rect 15947 -2638 15958 -2570
rect 16026 -2638 16035 -2570
rect 15947 -2650 16035 -2638
rect 16270 -2580 16350 -2564
rect 16270 -2640 16280 -2580
rect 16344 -2640 16350 -2580
rect 16270 -2657 16350 -2640
rect 15805 -2660 15868 -2658
rect 15805 -2675 15809 -2660
rect 15799 -2690 15809 -2675
rect 15863 -2675 15868 -2660
rect 15863 -2690 15870 -2675
rect 15799 -2746 15805 -2690
rect 15865 -2746 15870 -2690
rect 15799 -2760 15870 -2746
rect 16390 -2810 16520 -2800
rect 15527 -2829 16078 -2828
rect 16390 -2829 16410 -2810
rect 15527 -2870 16410 -2829
rect 16500 -2870 16520 -2810
rect 15527 -2889 16520 -2870
rect 16390 -2890 16520 -2889
rect 4260 -3140 9130 -2980
rect 9353 -3066 11621 -2970
rect 9447 -3068 11621 -3066
rect 16580 -3140 16910 -1260
rect -210 -3160 16910 -3140
rect -210 -3230 16900 -3160
rect -210 -3440 5410 -3230
rect 16400 -3440 16900 -3230
rect -210 -3480 16900 -3440
<< via2 >>
rect 4293 1911 4368 1971
rect -196 1481 -186 1580
rect -186 1481 -133 1580
rect -133 1481 -119 1580
rect 443 1481 500 1577
rect 500 1481 502 1577
rect 642 956 700 1030
rect 780 1480 783 1576
rect 783 1480 839 1576
rect 980 957 1038 1031
rect 1123 1481 1124 1577
rect 1124 1481 1182 1577
rect 1320 625 1323 687
rect 1323 625 1381 687
rect 1381 625 1382 687
rect 1318 309 1323 390
rect 1323 309 1378 390
rect 1463 1479 1467 1575
rect 1467 1479 1522 1575
rect 1667 613 1725 679
rect 1663 309 1667 390
rect 1667 309 1723 390
rect 1804 1479 1806 1575
rect 1806 1479 1863 1575
rect 2008 617 2065 674
rect 2004 309 2008 390
rect 2008 309 2064 390
rect 2148 1480 2153 1576
rect 2153 1480 2207 1576
rect 2489 1479 2490 1575
rect 2490 1479 2548 1575
rect 2690 602 2691 684
rect 2691 602 2749 684
rect 2749 602 2754 684
rect 2696 309 2749 390
rect 2749 309 2756 390
rect 2835 1480 2838 1576
rect 2838 1480 2894 1576
rect 3035 606 3036 681
rect 3036 606 3094 681
rect 3033 310 3036 391
rect 3036 310 3093 391
rect 3174 1480 3179 1576
rect 3179 1480 3233 1576
rect 3378 613 3379 679
rect 3379 613 3434 679
rect 3375 310 3379 391
rect 3379 310 3435 391
rect 3514 1479 3519 1575
rect 3519 1479 3573 1575
rect 3716 470 3719 548
rect 3719 470 3777 548
rect 3777 470 3779 548
rect 3855 1481 3858 1577
rect 3858 1481 3914 1577
rect 4061 958 4062 1032
rect 4062 958 4119 1032
rect 8573 1920 8630 1977
rect 9688 1941 9744 1942
rect 9688 1790 9691 1941
rect 9691 1790 9743 1941
rect 9743 1790 9744 1941
rect 4962 1310 4977 1419
rect 4977 1310 5022 1419
rect 4962 1309 5022 1310
rect 6710 1140 6717 1210
rect 6717 1140 6769 1210
rect 6769 1140 6770 1210
rect 7003 719 7066 791
rect 7334 718 7397 790
rect 7662 719 7725 791
rect 7989 719 8052 791
rect 8422 726 8480 791
rect 5259 556 5324 627
rect 5590 557 5655 628
rect 5918 555 5983 626
rect 6244 558 6309 629
rect 8274 564 8334 627
rect 5093 380 5154 450
rect 5427 382 5488 452
rect 5754 380 5815 450
rect 6083 386 6144 456
rect 6385 384 6446 454
rect 6834 379 6895 449
rect 7169 380 7230 450
rect 7497 381 7558 451
rect 7825 383 7886 453
rect 8129 386 8190 456
rect -43 -662 -42 -600
rect -42 -662 26 -600
rect -43 -664 26 -662
rect 728 -665 813 -608
rect 491 -1926 575 -1831
rect 2130 -460 2184 -344
rect 2184 -460 2186 -344
rect 1940 -973 2020 -904
rect 2265 -1182 2350 -1104
rect 3862 -1081 3983 -1072
rect 3862 -1082 3981 -1081
rect 3862 -1133 3878 -1082
rect 3878 -1133 3981 -1082
rect 3981 -1133 3983 -1081
rect 3897 -1302 3954 -1300
rect 3897 -1383 3900 -1302
rect 3900 -1383 3952 -1302
rect 3952 -1383 3954 -1302
rect 1628 -1816 1697 -1751
rect 734 -2200 812 -2135
rect 5095 -532 5155 -436
rect 5425 -530 5485 -434
rect 5754 -529 5814 -433
rect 6083 -530 6143 -434
rect 6389 -530 6449 -434
rect 6835 -528 6900 -444
rect 7167 -529 7232 -445
rect 7496 -531 7561 -447
rect 7826 -529 7891 -445
rect 8129 -528 8194 -444
rect 7004 -674 7069 -618
rect 7335 -675 7400 -619
rect 7662 -676 7727 -620
rect 7988 -676 8053 -620
rect 8272 -674 8335 -617
rect 5265 -842 5323 -778
rect 5592 -843 5650 -779
rect 5920 -843 5978 -779
rect 6247 -843 6305 -779
rect 8425 -837 8482 -781
rect 8419 -1604 8486 -1527
rect 9077 932 9135 954
rect 9077 898 9082 932
rect 9082 898 9134 932
rect 9134 898 9135 932
rect 9091 -900 9159 -811
rect 8617 -2010 8700 -1934
rect 9535 920 9591 976
rect 10053 1480 10149 1582
rect 13088 1488 13251 1640
rect 9540 239 9613 296
rect 9494 -675 9550 -619
rect 9868 -887 9959 -824
rect 9636 -1156 9730 -1097
rect 11605 -703 11719 -607
rect 10436 -1373 10503 -1309
rect 8963 -2203 9069 -2138
rect 9551 -2541 9610 -2454
rect 10120 -1521 10178 -1462
rect 9974 -2536 10030 -2450
rect 10258 -1669 10314 -1612
rect 11705 -1854 11778 -1782
rect 10439 -2161 10503 -2094
rect 11096 -2104 11164 -2098
rect 11096 -2158 11097 -2104
rect 11097 -2158 11162 -2104
rect 11162 -2158 11164 -2104
rect 11096 -2161 11164 -2158
rect 10942 -2583 10944 -2480
rect 10944 -2583 11020 -2480
rect 11020 -2583 11031 -2480
rect 10942 -2591 11031 -2583
rect 11533 -2257 11620 -2240
rect 11533 -2325 11606 -2257
rect 11606 -2325 11620 -2257
rect 14097 200 14192 287
rect 14955 -777 15027 -707
rect 13786 -1550 13893 -1481
rect 14471 -1549 14570 -1477
rect 12960 -2389 13028 -2318
rect 13028 -2389 13029 -2318
rect 13998 -2462 14054 -2461
rect 13998 -2520 14051 -2462
rect 14051 -2520 14054 -2462
rect 14497 -2382 14582 -2326
rect 14904 -2450 14973 -2394
rect 15149 -2442 15218 -2386
rect 15385 -2441 15454 -2385
rect 15958 -2638 16026 -2570
rect 16280 -2640 16344 -2580
rect 15805 -2720 15809 -2690
rect 15809 -2720 15863 -2690
rect 15863 -2720 15865 -2690
rect 15805 -2746 15865 -2720
rect 16410 -2870 16500 -2810
<< metal3 >>
rect 4282 1983 4377 1985
rect 4282 1977 9748 1983
rect 4282 1971 8573 1977
rect 4282 1911 4293 1971
rect 4368 1920 8573 1971
rect 8630 1942 9748 1977
rect 8630 1920 9688 1942
rect 4368 1911 9688 1920
rect 4282 1910 9688 1911
rect 4282 1899 4377 1910
rect 9678 1790 9688 1910
rect 9744 1790 9748 1942
rect 9678 1769 9748 1790
rect 13055 1649 13278 1657
rect 12483 1640 13278 1649
rect 12483 1606 13088 1640
rect 10608 1589 13088 1606
rect 4571 1587 13088 1589
rect -224 1582 13088 1587
rect -224 1580 10053 1582
rect -224 1481 -196 1580
rect -119 1577 10053 1580
rect -119 1481 443 1577
rect 502 1576 1123 1577
rect 502 1481 780 1576
rect -224 1480 780 1481
rect 839 1481 1123 1576
rect 1182 1576 3855 1577
rect 1182 1575 2148 1576
rect 1182 1481 1463 1575
rect 839 1480 1463 1481
rect -224 1479 1463 1480
rect 1522 1479 1804 1575
rect 1863 1480 2148 1575
rect 2207 1575 2835 1576
rect 2207 1480 2489 1575
rect 1863 1479 2489 1480
rect 2548 1480 2835 1575
rect 2894 1480 3174 1576
rect 3233 1575 3855 1576
rect 3233 1480 3514 1575
rect 2548 1479 3514 1480
rect 3573 1481 3855 1575
rect 3914 1494 10053 1577
rect 3914 1481 4892 1494
rect 3573 1479 4892 1481
rect -224 1471 4892 1479
rect 4571 1470 4892 1471
rect 5089 1480 10053 1494
rect 10149 1488 13088 1582
rect 13251 1488 13278 1640
rect 10149 1480 13278 1488
rect 5089 1470 13278 1480
rect 8339 1467 13278 1470
rect 12483 1465 13278 1467
rect 12483 1463 13270 1465
rect 4948 1419 5033 1438
rect 4948 1410 4962 1419
rect -396 1320 4962 1410
rect 4948 1309 4962 1320
rect 5022 1309 5033 1419
rect 4948 1290 5033 1309
rect -396 1210 6781 1220
rect -396 1140 6710 1210
rect 6770 1140 6781 1210
rect -396 1130 6781 1140
rect -442 1032 4168 1038
rect -442 1031 4061 1032
rect -442 1030 980 1031
rect -442 956 642 1030
rect 700 957 980 1030
rect 1038 958 4061 1031
rect 4119 958 4168 1032
rect 9527 976 9595 986
rect 9527 970 9535 976
rect 1038 957 4168 958
rect 700 956 4168 957
rect -442 949 4168 956
rect 9070 954 9535 970
rect -442 78 -366 949
rect 9070 898 9077 954
rect 9135 920 9535 954
rect 9591 920 9595 976
rect 9135 911 9595 920
rect 9135 898 9142 911
rect 9527 910 9595 911
rect 9070 888 9142 898
rect 6980 800 7368 801
rect 8303 800 8447 801
rect 6980 791 8491 800
rect 6980 719 7003 791
rect 7066 790 7662 791
rect 7066 719 7334 790
rect 6980 718 7334 719
rect 7397 719 7662 790
rect 7725 719 7989 791
rect 8052 726 8422 791
rect 8480 726 8491 791
rect 8052 719 8491 726
rect 7397 718 8491 719
rect 6980 711 8491 718
rect 1312 687 1386 698
rect 1312 625 1320 687
rect 1382 676 1386 687
rect 1657 679 1728 689
rect 1657 676 1667 679
rect 1382 625 1667 676
rect 1312 620 1667 625
rect 1312 606 1386 620
rect 1657 613 1667 620
rect 1725 676 1728 679
rect 1999 676 2069 691
rect 2675 684 2758 697
rect 2675 676 2690 684
rect 1725 674 2690 676
rect 1725 620 2008 674
rect 1725 613 1728 620
rect 1657 605 1728 613
rect 1999 617 2008 620
rect 2065 620 2690 674
rect 2065 617 2069 620
rect 1999 606 2069 617
rect 1661 602 1727 605
rect 2675 602 2690 620
rect 2754 676 2758 684
rect 3029 681 3098 693
rect 3029 676 3035 681
rect 2754 620 3035 676
rect 2754 602 2758 620
rect 2675 589 2758 602
rect 3029 606 3035 620
rect 3094 676 3098 681
rect 3366 679 3441 696
rect 3366 676 3378 679
rect 3094 620 3378 676
rect 3094 606 3098 620
rect 3029 594 3098 606
rect 3366 613 3378 620
rect 3434 676 3441 679
rect 3650 676 3921 677
rect 3434 671 3921 676
rect 3434 649 3922 671
rect 3434 620 4871 649
rect 3434 613 3441 620
rect 3735 619 4871 620
rect 3366 601 3441 613
rect 3873 586 4871 619
rect 4600 585 4871 586
rect 5244 629 8341 638
rect 5244 628 6244 629
rect 5244 627 5590 628
rect 3701 548 3790 559
rect 3701 470 3716 548
rect 3779 525 3790 548
rect 3779 524 4384 525
rect 3779 470 4713 524
rect 3701 459 4713 470
rect 4030 458 4713 459
rect 4775 460 4870 585
rect 5244 556 5259 627
rect 5324 557 5590 627
rect 5655 626 6244 628
rect 5655 557 5918 626
rect 5324 556 5918 557
rect 5244 555 5918 556
rect 5983 558 6244 626
rect 6309 627 8341 629
rect 6309 564 8274 627
rect 8334 564 8341 627
rect 6309 558 8341 564
rect 5983 555 8341 558
rect 5244 548 8341 555
rect 8283 547 8341 548
rect 1296 391 4519 400
rect 1296 390 3033 391
rect 1296 309 1318 390
rect 1378 309 1663 390
rect 1723 309 2004 390
rect 2064 309 2696 390
rect 2756 310 3033 390
rect 3093 310 3375 391
rect 3435 310 4519 391
rect 2756 309 4519 310
rect 1296 300 4519 309
rect 4418 231 4518 300
rect 4651 296 4708 458
rect 4775 456 8337 460
rect 4775 452 6083 456
rect 4775 450 5427 452
rect 4775 380 5093 450
rect 5154 382 5427 450
rect 5488 450 6083 452
rect 5488 382 5754 450
rect 5154 380 5754 382
rect 5815 386 6083 450
rect 6144 454 8129 456
rect 6144 386 6385 454
rect 5815 384 6385 386
rect 6446 453 8129 454
rect 6446 451 7825 453
rect 6446 450 7497 451
rect 6446 449 7169 450
rect 6446 384 6834 449
rect 5815 380 6834 384
rect 4775 379 6834 380
rect 6895 380 7169 449
rect 7230 381 7497 450
rect 7558 383 7825 451
rect 7886 386 8129 453
rect 8190 386 8337 456
rect 7886 383 8337 386
rect 7558 381 8337 383
rect 7230 380 8337 381
rect 6895 379 8337 380
rect 4775 371 8337 379
rect 4808 370 8337 371
rect 9527 301 9622 312
rect 9527 299 14202 301
rect 9391 297 14202 299
rect 5080 296 14202 297
rect 4651 241 9540 296
rect 4651 240 6032 241
rect 6448 240 9399 241
rect 1624 79 2158 81
rect -258 78 2195 79
rect -443 3 2195 78
rect -443 0 1676 3
rect -443 -1 1572 0
rect -442 -6 -366 -1
rect 2117 -329 2195 3
rect 4417 -6 4518 231
rect 9527 239 9540 241
rect 9613 287 14202 296
rect 9613 239 14097 287
rect 9527 230 14097 239
rect 9527 227 9622 230
rect 14076 200 14097 230
rect 14192 200 14202 287
rect 14076 184 14202 200
rect 4417 -7 4790 -6
rect 4417 -58 4935 -7
rect 4418 -106 4935 -58
rect 2116 -344 2195 -329
rect 2116 -460 2130 -344
rect 2186 -460 2195 -344
rect 2116 -474 2195 -460
rect 4834 -429 4934 -106
rect 4834 -430 8064 -429
rect 4834 -433 8206 -430
rect 4834 -434 5754 -433
rect 4834 -436 5425 -434
rect 4834 -532 5095 -436
rect 5155 -530 5425 -436
rect 5485 -529 5754 -434
rect 5814 -434 8206 -433
rect 5814 -529 6083 -434
rect 5485 -530 6083 -529
rect 6143 -530 6389 -434
rect 6449 -444 8206 -434
rect 6449 -528 6835 -444
rect 6900 -445 8129 -444
rect 6900 -528 7167 -445
rect 6449 -529 7167 -528
rect 7232 -447 7826 -445
rect 7232 -529 7496 -447
rect 6449 -530 7496 -529
rect 5155 -531 7496 -530
rect 7561 -529 7826 -447
rect 7891 -528 8129 -445
rect 8194 -528 8206 -444
rect 7891 -529 8206 -528
rect 7561 -531 8206 -529
rect 5155 -532 8206 -531
rect 4834 -540 8206 -532
rect 4834 -555 4933 -540
rect -60 -598 42 -583
rect -60 -600 824 -598
rect -60 -664 -43 -600
rect 26 -608 824 -600
rect 11566 -607 11749 -579
rect 8259 -608 8345 -607
rect 11566 -608 11605 -607
rect 26 -664 728 -608
rect -60 -665 728 -664
rect 813 -665 824 -608
rect 8053 -617 11605 -608
rect -60 -670 824 -665
rect 6830 -618 8272 -617
rect -60 -680 42 -670
rect 6830 -674 7004 -618
rect 7069 -619 8272 -618
rect 7069 -674 7335 -619
rect 6830 -675 7335 -674
rect 7400 -620 8272 -619
rect 7400 -675 7662 -620
rect 6830 -676 7662 -675
rect 7727 -676 7988 -620
rect 8053 -674 8272 -620
rect 8335 -619 11605 -617
rect 8335 -674 9494 -619
rect 8053 -675 9494 -674
rect 9550 -675 11605 -619
rect 8053 -676 11605 -675
rect 6830 -680 11605 -676
rect 7925 -681 11605 -680
rect 8259 -682 9560 -681
rect 8259 -684 8345 -682
rect 11566 -703 11605 -681
rect 11719 -703 11749 -607
rect 11566 -739 11749 -703
rect 14940 -707 15037 -695
rect 5241 -769 8367 -768
rect 5241 -778 8492 -769
rect 5241 -842 5265 -778
rect 5323 -779 8492 -778
rect 5323 -842 5592 -779
rect 5241 -843 5592 -842
rect 5650 -843 5920 -779
rect 5978 -843 6247 -779
rect 6305 -781 8492 -779
rect 6305 -837 8425 -781
rect 8482 -837 8492 -781
rect 14940 -777 14955 -707
rect 15027 -777 15037 -707
rect 6305 -843 8492 -837
rect 5241 -849 8492 -843
rect 5365 -850 8492 -849
rect 9079 -811 9171 -801
rect -433 -904 2036 -887
rect -433 -973 1940 -904
rect 2020 -973 2036 -904
rect 9079 -900 9091 -811
rect 9159 -812 9171 -811
rect 9159 -824 9970 -812
rect 9159 -887 9868 -824
rect 9959 -887 9970 -824
rect 9159 -900 9970 -887
rect 9079 -913 9171 -900
rect -433 -988 2036 -973
rect 1926 -990 2036 -988
rect 3803 -1072 4061 -1054
rect -423 -1091 1984 -1089
rect -423 -1104 2360 -1091
rect -423 -1182 2265 -1104
rect 2350 -1182 2360 -1104
rect 3803 -1133 3862 -1072
rect 3983 -1078 4061 -1072
rect 3983 -1079 4066 -1078
rect 3983 -1097 9750 -1079
rect 3983 -1133 9636 -1097
rect 3803 -1146 9636 -1133
rect 4035 -1148 9636 -1146
rect 9609 -1156 9636 -1148
rect 9730 -1156 9750 -1097
rect 9609 -1173 9750 -1156
rect -423 -1191 2360 -1182
rect 1847 -1193 2360 -1191
rect 3884 -1295 3960 -1287
rect 3884 -1296 9370 -1295
rect 3884 -1300 10511 -1296
rect 10570 -1299 10645 -1298
rect 14940 -1299 15037 -777
rect 3884 -1383 3897 -1300
rect 3954 -1309 10511 -1300
rect 3954 -1373 10436 -1309
rect 10503 -1373 10511 -1309
rect 3954 -1383 10511 -1373
rect 3884 -1387 10511 -1383
rect 10569 -1300 10897 -1299
rect 11540 -1300 15037 -1299
rect 10569 -1319 15037 -1300
rect 15553 -1319 15621 -1317
rect 10569 -1387 15621 -1319
rect 3884 -1400 3960 -1387
rect 10569 -1389 15037 -1387
rect 10569 -1390 11546 -1389
rect 10112 -1457 10190 -1453
rect 10570 -1457 10645 -1390
rect 14940 -1392 15037 -1389
rect 10109 -1462 10645 -1457
rect 8407 -1520 8495 -1518
rect 9946 -1520 10042 -1518
rect 8407 -1527 10042 -1520
rect 8407 -1604 8419 -1527
rect 8486 -1604 10042 -1527
rect 10109 -1521 10120 -1462
rect 10178 -1521 10645 -1462
rect 14471 -1472 14587 -1471
rect 13765 -1474 13903 -1473
rect 14078 -1474 14590 -1472
rect 10703 -1476 14590 -1474
rect 10109 -1531 10645 -1521
rect 10702 -1477 14590 -1476
rect 10702 -1481 14471 -1477
rect 10702 -1550 13786 -1481
rect 13893 -1549 14471 -1481
rect 14570 -1549 14590 -1477
rect 13893 -1550 14590 -1549
rect 10702 -1560 14590 -1550
rect 10702 -1562 14577 -1560
rect 10702 -1564 14105 -1562
rect 10702 -1594 10779 -1564
rect 10312 -1595 10779 -1594
rect 8407 -1615 10042 -1604
rect 8407 -1616 8495 -1615
rect 1620 -1744 4897 -1743
rect 1620 -1746 5667 -1744
rect 9158 -1746 9235 -1744
rect 1620 -1751 9235 -1746
rect 482 -1831 591 -1813
rect 1620 -1816 1628 -1751
rect 1697 -1816 9235 -1751
rect 1620 -1823 9235 -1816
rect 3011 -1824 9235 -1823
rect 482 -1926 491 -1831
rect 575 -1920 591 -1831
rect 575 -1926 8708 -1920
rect 482 -1934 8708 -1926
rect 482 -2010 8617 -1934
rect 8700 -2010 8708 -1934
rect 482 -2032 8708 -2010
rect 585 -2033 8708 -2032
rect 9158 -2004 9235 -1824
rect 9946 -1770 10042 -1615
rect 10245 -1612 10779 -1595
rect 10245 -1669 10258 -1612
rect 10314 -1669 10779 -1612
rect 10245 -1671 10703 -1669
rect 10245 -1682 10319 -1671
rect 10370 -1770 11785 -1769
rect 9946 -1782 11785 -1770
rect 9946 -1854 11705 -1782
rect 11778 -1854 11785 -1782
rect 15553 -1839 15621 -1387
rect 9946 -1866 11785 -1854
rect 9946 -1869 10042 -1866
rect 15551 -1906 16587 -1839
rect 719 -2127 8916 -2126
rect 719 -2135 9079 -2127
rect 719 -2200 734 -2135
rect 812 -2138 9079 -2135
rect 812 -2200 8963 -2138
rect 719 -2203 8963 -2200
rect 9069 -2203 9079 -2138
rect 719 -2208 9079 -2203
rect 1693 -2209 9079 -2208
rect 1693 -2210 7945 -2209
rect 8122 -2212 9079 -2209
rect 9158 -2211 9237 -2004
rect 11521 -2021 14410 -2020
rect 14819 -2021 14886 -2020
rect 10426 -2065 10504 -2064
rect 10426 -2084 10511 -2065
rect 10425 -2094 11174 -2084
rect 10425 -2161 10439 -2094
rect 10503 -2098 11175 -2094
rect 10503 -2161 11096 -2098
rect 11164 -2161 11175 -2098
rect 10425 -2166 11175 -2161
rect 9160 -2307 9237 -2211
rect 9157 -2314 9237 -2307
rect 10426 -2176 11175 -2166
rect 11521 -2123 14921 -2021
rect 11521 -2124 14410 -2123
rect 9157 -2372 9239 -2314
rect 10426 -2317 10504 -2176
rect 11521 -2222 11625 -2124
rect 9154 -2717 9239 -2372
rect 9551 -2385 10504 -2317
rect 11513 -2240 11636 -2222
rect 11513 -2325 11533 -2240
rect 11620 -2325 11636 -2240
rect 11513 -2342 11636 -2325
rect 12947 -2318 13042 -2307
rect 9551 -2390 10040 -2385
rect 10426 -2386 10504 -2385
rect 10440 -2388 10504 -2386
rect 9551 -2404 9622 -2390
rect 9544 -2440 9622 -2404
rect 9544 -2454 9621 -2440
rect 9544 -2541 9551 -2454
rect 9610 -2541 9621 -2454
rect 9544 -2555 9621 -2541
rect 9961 -2447 10040 -2390
rect 12947 -2389 12960 -2318
rect 13029 -2319 13042 -2318
rect 13029 -2326 14632 -2319
rect 13029 -2382 14497 -2326
rect 14582 -2382 14632 -2326
rect 14819 -2358 14921 -2123
rect 13029 -2389 14632 -2382
rect 14818 -2385 15528 -2358
rect 16520 -2374 16587 -1906
rect 16520 -2376 16611 -2374
rect 14818 -2386 15385 -2385
rect 12947 -2399 13042 -2389
rect 14818 -2394 15149 -2386
rect 9961 -2450 10039 -2447
rect 14818 -2450 14904 -2394
rect 14973 -2442 15149 -2394
rect 15218 -2441 15385 -2386
rect 15454 -2441 15528 -2385
rect 15218 -2442 15528 -2441
rect 14973 -2450 15528 -2442
rect 9961 -2536 9974 -2450
rect 10030 -2536 10039 -2450
rect 13982 -2461 14079 -2450
rect 14818 -2461 15528 -2450
rect 9961 -2556 10039 -2536
rect 10925 -2480 11042 -2463
rect 10925 -2591 10942 -2480
rect 11031 -2591 11042 -2480
rect 10925 -2614 11042 -2591
rect 13982 -2520 13998 -2461
rect 14054 -2520 14079 -2461
rect 14819 -2464 14921 -2461
rect 16519 -2463 17075 -2376
rect 15947 -2481 16035 -2480
rect 13982 -2580 14079 -2520
rect 15655 -2559 16035 -2481
rect 15655 -2580 15734 -2559
rect 10925 -2717 11041 -2614
rect 13982 -2658 15734 -2580
rect 15947 -2569 16035 -2559
rect 15947 -2570 16361 -2569
rect 16523 -2570 16611 -2463
rect 15947 -2638 15958 -2570
rect 16026 -2580 16611 -2570
rect 16026 -2638 16280 -2580
rect 15947 -2640 16280 -2638
rect 16344 -2640 16611 -2580
rect 15947 -2649 16611 -2640
rect 16780 -2640 17080 -2550
rect 15947 -2650 16525 -2649
rect 13982 -2659 15523 -2658
rect 15655 -2659 15734 -2658
rect 9154 -2718 11041 -2717
rect 15799 -2690 15870 -2675
rect 15799 -2718 15805 -2690
rect 9154 -2746 15805 -2718
rect 15865 -2746 15870 -2690
rect 9154 -2806 15870 -2746
rect 16780 -2800 16870 -2640
rect 9154 -2808 9281 -2806
rect 16390 -2810 16870 -2800
rect 16390 -2870 16410 -2810
rect 16500 -2870 16870 -2810
rect 16390 -2890 16870 -2870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  gf180mcu_fd_sc_mcu7t5v0__inv_1_0 ~/conda-gf180mcu-env/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1757859342
transform 1 0 -119 0 1 -1023
box -86 -86 534 870
use nfet_03v3_1_028  nfet_03v3_1_028_0
timestamp 1757730057
transform 1 0 8873 0 1 694
box 0 0 280 416
use nfet_03v3_2_2_028  nfet_03v3_2_2_028_0
timestamp 1757729720
transform -1 0 3575 0 -1 -1071
box 0 0 440 622
use nfet_03v3_2_2_028  nfet_03v3_2_2_028_1
timestamp 1757729720
transform 1 0 3700 0 1 -1693
box 0 0 440 622
use nfet_03v3_2_028  nfet_03v3_2_028_0
timestamp 1757729325
transform 1 0 2700 0 1 -1678
box 0 0 280 593
use nfet_03v3_2_028  nfet_03v3_2_028_1
timestamp 1757729325
transform -1 0 10980 0 -1 -2152
box 0 0 280 593
use nfet_03v3_2_028  nfet_03v3_2_028_2
timestamp 1757729325
transform 1 0 10988 0 1 -2688
box 0 0 280 593
use nfet_03v3_2_028  nfet_03v3_2_028_3
timestamp 1757729325
transform -1 0 11560 0 -1 -2153
box 0 0 280 593
use nfet_03v3_2_028  nfet_03v3_2_028_4
timestamp 1757729325
transform 1 0 11572 0 1 -2691
box 0 0 280 593
use nfet_03v3_4_2_08  nfet_03v3_4_2_08_0
timestamp 1757728578
transform 1 0 14789 0 1 -2834
box 0 0 760 591
use nfet_03v3_4_2_08  nfet_03v3_4_2_08_1
timestamp 1757728578
transform 1 0 15769 0 1 -2839
box 0 0 760 591
use nfet_03v3_05_05  nfet_03v3_05_05_0
timestamp 1757727608
transform -1 0 10028 0 -1 -2414
box -28 -26 501 285
use nfet_03v3_8_028  nfet_03v3_8_028_0
timestamp 1757730643
transform 1 0 8880 0 1 -1423
box 0 -97 280 1816
use pfet_03v3_1_1  pfet_03v3_1_1_0
timestamp 1757817671
transform -1 0 2581 0 -1 -182
box -117 -108 982 654
use pfet_03v3_1_028  pfet_03v3_1_028_0
timestamp 1757722512
transform -1 0 9000 0 -1 2060
box -151 -136 513 649
use pfet_03v3_2_24_03  pfet_03v3_2_24_03_0
timestamp 1757727097
transform 1 0 4994 0 1 104
box -334 -2650 3601 2164
use pfet_03v3_4_8_028  pfet_03v3_4_8_028_0
timestamp 1757847982
transform 1 0 12390 0 1 -2677
box 0 0 884 660
use pfet_03v3_4_8_028  pfet_03v3_4_8_028_1
timestamp 1757847982
transform 1 0 13420 0 1 -2679
box 0 0 884 660
use pfet_03v3_8_05  pfet_03v3_8_05_0
timestamp 1757750971
transform 1 0 111 0 1 170
box -111 -170 4560 1880
use ppolyf_res  ppolyf_res_0
timestamp 1757840551
transform 0 -1 14686 1 0 -1210
box -60 -60 3412 5256
<< labels >>
flabel metal3 -393 1324 -300 1406 0 FreeSans 160 0 0 0 IN_P
flabel metal3 -390 1135 -297 1217 0 FreeSans 160 0 0 0 IN_N
flabel metal2 -436 -657 -365 -604 0 FreeSans 160 0 0 0 EN
flabel metal3 -425 -984 -335 -896 0 FreeSans 160 0 0 0 CAL_P
flabel metal3 -415 -1183 -325 -1095 0 FreeSans 160 0 0 0 CAL_N
flabel metal3 16940 -2460 17070 -2380 0 FreeSans 160 0 0 0 OUT_N
flabel metal3 16940 -2640 17070 -2550 0 FreeSans 160 0 0 0 OUT_P
flabel metal2 -200 2160 130 2350 0 FreeSans 320 0 0 0 VDD
flabel metal2 -90 -1810 240 -1620 0 FreeSans 320 0 0 0 VSS
<< end >>
