magic
tech gf180mcuD
magscale 1 10
timestamp 1757239750
<< nwell >>
rect 2721 2575 3605 4676
rect 2721 2574 3606 2575
rect 2720 2376 3606 2574
rect 2722 2308 3606 2376
rect 2722 2306 3603 2308
<< pwell >>
rect 3683 4674 4444 4676
rect 3619 4402 4444 4674
rect 3619 4363 4009 4402
rect 4112 4363 4444 4402
rect 3619 3641 4444 4363
rect 3619 2578 4812 3641
rect 3619 2404 4831 2578
rect 3619 2307 4812 2404
rect 4423 2305 4812 2307
rect 2088 11 2091 1074
rect 2088 -262 2091 -163
<< nmos >>
rect 3793 2695 3849 4295
rect 3953 2695 4009 4295
rect 4113 2695 4169 4295
rect 4273 2695 4329 4295
rect 4591 2707 4647 3507
<< pmos >>
rect 2895 2697 2951 4297
rect 3055 2697 3111 4297
rect 3215 2697 3271 4297
rect 3375 2697 3431 4297
<< ndiff >>
rect 3705 4282 3793 4295
rect 3705 2708 3718 4282
rect 3764 2708 3793 4282
rect 3705 2695 3793 2708
rect 3849 4282 3953 4295
rect 3849 2708 3878 4282
rect 3924 2708 3953 4282
rect 3849 2695 3953 2708
rect 4009 4282 4113 4295
rect 4009 2708 4038 4282
rect 4084 2708 4113 4282
rect 4009 2695 4113 2708
rect 4169 4282 4273 4295
rect 4169 2708 4198 4282
rect 4244 2708 4273 4282
rect 4169 2695 4273 2708
rect 4329 4282 4417 4295
rect 4329 2708 4358 4282
rect 4404 2708 4417 4282
rect 4329 2695 4417 2708
rect 4491 3487 4591 3507
rect 4491 2726 4510 3487
rect 4557 2726 4591 3487
rect 4491 2707 4591 2726
rect 4647 3488 4747 3507
rect 4647 2727 4681 3488
rect 4728 2727 4747 3488
rect 4647 2707 4747 2727
<< pdiff >>
rect 2807 4284 2895 4297
rect 2807 2710 2820 4284
rect 2866 2710 2895 4284
rect 2807 2697 2895 2710
rect 2951 4284 3055 4297
rect 2951 2710 2980 4284
rect 3026 2710 3055 4284
rect 2951 2697 3055 2710
rect 3111 4284 3215 4297
rect 3111 2710 3140 4284
rect 3186 2710 3215 4284
rect 3111 2697 3215 2710
rect 3271 4284 3375 4297
rect 3271 2710 3300 4284
rect 3346 2710 3375 4284
rect 3271 2697 3375 2710
rect 3431 4284 3519 4297
rect 3431 2710 3460 4284
rect 3506 2710 3519 4284
rect 3431 2697 3519 2710
<< ndiffc >>
rect 3718 2708 3764 4282
rect 3878 2708 3924 4282
rect 4038 2708 4084 4282
rect 4198 2708 4244 4282
rect 4358 2708 4404 4282
rect 4510 2726 4557 3487
rect 4681 2727 4728 3488
<< pdiffc >>
rect 2820 2710 2866 4284
rect 2980 2710 3026 4284
rect 3140 2710 3186 4284
rect 3300 2710 3346 4284
rect 3460 2710 3506 4284
<< psubdiff >>
rect 4414 2577 4831 2578
rect 3656 2532 4831 2577
rect 3656 2439 3761 2532
rect 4378 2439 4831 2532
rect 3656 2409 4831 2439
rect 4414 2404 4831 2409
<< nsubdiff >>
rect 2791 4609 3558 4652
rect 2791 4517 2849 4609
rect 3454 4517 3558 4609
rect 2791 4485 3558 4517
<< psubdiffcont >>
rect 3761 2439 4378 2532
<< nsubdiffcont >>
rect 2849 4517 3454 4609
<< polysilicon >>
rect 2895 4337 3431 4386
rect 2895 4297 2951 4337
rect 3055 4297 3111 4337
rect 3215 4297 3271 4337
rect 3375 4297 3431 4337
rect 3793 4337 4009 4386
rect 4112 4337 4329 4386
rect 3793 4295 3849 4337
rect 3953 4295 4009 4337
rect 4113 4295 4169 4337
rect 4273 4295 4329 4337
rect 2895 2653 2951 2697
rect 3055 2653 3111 2697
rect 3215 2653 3271 2697
rect 3375 2653 3431 2697
rect 4562 3549 4671 3622
rect 4591 3507 4647 3549
rect 3793 2651 3849 2695
rect 3953 2651 4009 2695
rect 4113 2651 4169 2695
rect 4273 2651 4329 2695
rect 4591 2661 4647 2707
<< metal1 >>
rect 2791 4609 3558 4652
rect 2791 4517 2849 4609
rect 3454 4517 3558 4609
rect 2791 4485 3558 4517
rect 2820 4284 2866 4295
rect 2980 4284 3026 4295
rect 2866 4242 2873 4254
rect 2872 4167 2873 4242
rect 2866 4154 2873 4167
rect 2820 2699 2866 2710
rect 3140 4284 3186 4295
rect 3300 4284 3346 4295
rect 3186 4242 3193 4254
rect 3192 4167 3193 4242
rect 3026 2820 3037 2833
rect 3036 2749 3037 2820
rect 3026 2737 3037 2749
rect 2980 2699 3026 2710
rect 3186 4154 3193 4167
rect 3140 2699 3186 2710
rect 3460 4284 3506 4295
rect 3718 4282 3764 4293
rect 3506 4232 3513 4244
rect 3346 2819 3356 2833
rect 3346 2735 3356 2748
rect 3300 2699 3346 2710
rect 3506 4143 3513 4157
rect 3460 2699 3506 2710
rect 3878 4282 3924 4293
rect 3764 2822 3780 2836
rect 3774 2751 3780 2822
rect 3764 2738 3780 2751
rect 3718 2697 3764 2708
rect 3878 2697 3924 2708
rect 4038 4282 4084 4293
rect 4198 4282 4244 4293
rect 4084 2827 4095 2841
rect 4094 2756 4095 2827
rect 4084 2743 4095 2756
rect 4038 2697 4084 2708
rect 4198 2697 4244 2708
rect 4358 4282 4404 4293
rect 4515 3499 4581 3500
rect 4502 3487 4581 3499
rect 4404 2828 4415 2842
rect 4413 2757 4415 2828
rect 4404 2744 4415 2757
rect 4502 2726 4510 3487
rect 4557 2726 4581 3487
rect 4502 2709 4581 2726
rect 4657 3488 4736 3505
rect 4657 2727 4681 3488
rect 4728 2847 4736 3488
rect 4728 2832 4739 2847
rect 4737 2761 4739 2832
rect 4728 2750 4739 2761
rect 4728 2749 4737 2750
rect 4728 2727 4736 2749
rect 4657 2715 4736 2727
rect 4657 2714 4723 2715
rect 4358 2697 4404 2708
rect 4414 2577 4831 2578
rect 3656 2532 4831 2577
rect 3656 2439 3761 2532
rect 4378 2439 4831 2532
rect 3656 2409 4831 2439
rect 4414 2404 4831 2409
<< via1 >>
rect 2820 4167 2866 4242
rect 2866 4167 2872 4242
rect 3140 4167 3186 4242
rect 3186 4167 3192 4242
rect 2981 2749 3026 2820
rect 3026 2749 3036 2820
rect 3461 4157 3506 4232
rect 3506 4157 3513 4232
rect 3301 2748 3346 2819
rect 3346 2748 3356 2819
rect 3719 2751 3764 2822
rect 3764 2751 3774 2822
rect 4039 2756 4084 2827
rect 4084 2756 4094 2827
rect 4358 2757 4404 2828
rect 4404 2757 4413 2828
rect 4682 2761 4728 2832
rect 4728 2761 4737 2832
<< metal2 >>
rect 2808 4242 3524 4245
rect 2808 4167 2820 4242
rect 2872 4167 3140 4242
rect 3192 4232 3524 4242
rect 3192 4167 3461 4232
rect 2808 4157 3461 4167
rect 3513 4157 3524 4232
rect 2808 4146 3524 4157
rect 2970 2832 4754 2844
rect 2970 2828 4682 2832
rect 2970 2827 4358 2828
rect 2970 2822 4039 2827
rect 2970 2820 3719 2822
rect 2970 2749 2981 2820
rect 3036 2819 3719 2820
rect 3036 2749 3301 2819
rect 2970 2748 3301 2749
rect 3356 2751 3719 2819
rect 3774 2756 4039 2822
rect 4094 2757 4358 2827
rect 4413 2761 4682 2828
rect 4737 2761 4754 2832
rect 4413 2757 4754 2761
rect 4094 2756 4754 2757
rect 3774 2751 4754 2756
rect 3356 2748 4754 2751
rect 2970 2737 4754 2748
<< labels >>
flabel metal1 3880 2901 3922 3499 0 FreeSans 320 0 0 0 VCM
port 1 nsew
flabel metal1 4200 2893 4242 3499 0 FreeSans 160 0 0 0 VREF_GND
port 2 nsew
flabel metal1 4509 2870 4573 3412 0 FreeSans 160 0 0 0 VIN
port 3 nsew
flabel metal2 2880 4166 3400 4223 0 FreeSans 320 0 0 0 VREF
port 4 nsew
flabel polysilicon 3796 4339 4007 4382 0 FreeSans 160 0 0 0 EN_VCM
port 5 nsew
flabel polysilicon 2906 4340 3426 4382 0 FreeSans 160 0 0 0 EN_VREF_Z
port 6 nsew
flabel metal2 3242 2745 3982 2827 0 FreeSans 320 0 0 0 Cbtm
port 7 nsew
flabel metal1 2826 4500 3534 4631 0 FreeSans 320 0 0 0 VDD
port 8 nsew
flabel polysilicon 4123 4344 4324 4383 0 FreeSans 160 0 0 0 EN_VSS
port 9 nsew
flabel polysilicon 4567 3554 4667 3618 0 FreeSans 160 0 0 0 EN_VIN
port 10 nsew
flabel metal1 3767 2420 4635 2539 0 FreeSans 320 0 0 0 VSS
port 11 nsew
<< end >>
