magic
tech gf180mcuD
magscale 1 10
timestamp 1757514455
<< nwell >>
rect -1250 -3442 1250 3442
<< pmos >>
rect -1000 1232 1000 3232
rect -1000 -1000 1000 1000
rect -1000 -3232 1000 -1232
<< pdiff >>
rect -1088 3219 -1000 3232
rect -1088 1245 -1075 3219
rect -1029 1245 -1000 3219
rect -1088 1232 -1000 1245
rect 1000 3219 1088 3232
rect 1000 1245 1029 3219
rect 1075 1245 1088 3219
rect 1000 1232 1088 1245
rect -1088 987 -1000 1000
rect -1088 -987 -1075 987
rect -1029 -987 -1000 987
rect -1088 -1000 -1000 -987
rect 1000 987 1088 1000
rect 1000 -987 1029 987
rect 1075 -987 1088 987
rect 1000 -1000 1088 -987
rect -1088 -1245 -1000 -1232
rect -1088 -3219 -1075 -1245
rect -1029 -3219 -1000 -1245
rect -1088 -3232 -1000 -3219
rect 1000 -1245 1088 -1232
rect 1000 -3219 1029 -1245
rect 1075 -3219 1088 -1245
rect 1000 -3232 1088 -3219
<< pdiffc >>
rect -1075 1245 -1029 3219
rect 1029 1245 1075 3219
rect -1075 -987 -1029 987
rect 1029 -987 1075 987
rect -1075 -3219 -1029 -1245
rect 1029 -3219 1075 -1245
<< nsubdiff >>
rect -1226 3346 1226 3418
rect -1226 3302 -1154 3346
rect -1226 -3302 -1213 3302
rect -1167 -3302 -1154 3302
rect 1154 3302 1226 3346
rect -1226 -3346 -1154 -3302
rect 1154 -3302 1167 3302
rect 1213 -3302 1226 3302
rect 1154 -3346 1226 -3302
rect -1226 -3418 1226 -3346
<< nsubdiffcont >>
rect -1213 -3302 -1167 3302
rect 1167 -3302 1213 3302
<< polysilicon >>
rect -1000 3311 1000 3324
rect -1000 3265 -987 3311
rect 987 3265 1000 3311
rect -1000 3232 1000 3265
rect -1000 1199 1000 1232
rect -1000 1153 -987 1199
rect 987 1153 1000 1199
rect -1000 1140 1000 1153
rect -1000 1079 1000 1092
rect -1000 1033 -987 1079
rect 987 1033 1000 1079
rect -1000 1000 1000 1033
rect -1000 -1033 1000 -1000
rect -1000 -1079 -987 -1033
rect 987 -1079 1000 -1033
rect -1000 -1092 1000 -1079
rect -1000 -1153 1000 -1140
rect -1000 -1199 -987 -1153
rect 987 -1199 1000 -1153
rect -1000 -1232 1000 -1199
rect -1000 -3265 1000 -3232
rect -1000 -3311 -987 -3265
rect 987 -3311 1000 -3265
rect -1000 -3324 1000 -3311
<< polycontact >>
rect -987 3265 987 3311
rect -987 1153 987 1199
rect -987 1033 987 1079
rect -987 -1079 987 -1033
rect -987 -1199 987 -1153
rect -987 -3311 987 -3265
<< metal1 >>
rect -1213 3359 1213 3405
rect -1213 3302 -1167 3359
rect -998 3265 -987 3311
rect 987 3265 998 3311
rect 1167 3302 1213 3359
rect -1075 3219 -1029 3230
rect -1075 1234 -1029 1245
rect 1029 3219 1075 3230
rect 1029 1234 1075 1245
rect -998 1153 -987 1199
rect 987 1153 998 1199
rect -998 1033 -987 1079
rect 987 1033 998 1079
rect -1075 987 -1029 998
rect -1075 -998 -1029 -987
rect 1029 987 1075 998
rect 1029 -998 1075 -987
rect -998 -1079 -987 -1033
rect 987 -1079 998 -1033
rect -998 -1199 -987 -1153
rect 987 -1199 998 -1153
rect -1075 -1245 -1029 -1234
rect -1075 -3230 -1029 -3219
rect 1029 -1245 1075 -1234
rect 1029 -3230 1075 -3219
rect -1213 -3359 -1167 -3302
rect -998 -3311 -987 -3265
rect 987 -3311 998 -3265
rect 1167 -3359 1213 -3302
rect -1213 -3405 1213 -3359
<< properties >>
string FIXED_BBOX -1190 -3382 1190 3382
string gencell pfet_03v3
string library gf180mcu
string parameters w 10 l 10 m 3 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {pfet_03v3 pfet_06v0}
<< end >>
