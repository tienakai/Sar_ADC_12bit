magic
tech gf180mcuD
magscale 1 10
timestamp 1757722512
<< nwell >>
rect -151 -136 513 649
<< nsubdiff >>
rect -123 570 440 590
rect -123 523 -14 570
rect 355 523 440 570
rect -123 510 440 523
rect -123 476 -41 510
rect -123 -12 -110 476
rect -56 -12 -41 476
rect 361 473 440 510
rect -123 -31 -41 -12
rect 361 30 378 473
rect 424 30 440 473
rect 361 -31 440 30
rect -123 -45 440 -31
rect -123 -92 -14 -45
rect 355 -92 440 -45
rect -123 -105 440 -92
<< nsubdiffcont >>
rect -14 523 355 570
rect -110 -12 -56 476
rect 378 30 424 473
rect -14 -92 355 -45
<< polysilicon >>
rect 120 413 201 428
rect 120 367 135 413
rect 188 367 201 413
rect 120 355 201 367
rect 130 354 201 355
rect 130 340 186 354
<< polycontact >>
rect 135 367 188 413
<< metal1 >>
rect -123 570 440 590
rect -123 523 -14 570
rect 355 523 440 570
rect -123 510 440 523
rect -123 476 -41 510
rect -123 -12 -110 476
rect -56 -12 -41 476
rect 361 473 440 510
rect 113 413 205 445
rect 113 367 135 413
rect 188 367 205 413
rect 113 360 205 367
rect -123 -31 -41 -12
rect 361 30 378 473
rect 424 30 440 473
rect 361 -31 440 30
rect -123 -45 440 -31
rect -123 -92 -14 -45
rect 355 -92 440 -45
rect -123 -105 440 -92
use pfet_03v3_9MEGGS  pfet_03v3_9MEGGS_0
timestamp 1757722512
transform 1 0 158 0 1 199
box -202 -230 202 230
<< end >>
