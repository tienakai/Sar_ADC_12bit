magic
tech gf180mcuD
magscale 1 10
timestamp 1757654639
<< nwell >>
rect 2044 8986 10762 9646
rect 2044 6460 9136 8986
rect 9306 7736 9710 8862
rect 9878 7786 10762 8986
rect 14288 5848 17036 10282
<< pwell >>
rect 10850 7584 12406 9560
rect 9368 6648 11916 7584
rect 9658 5872 11916 6648
rect 14124 5885 14134 5985
rect 9658 5848 12384 5872
rect 11764 5845 12384 5848
rect 11778 5806 12384 5845
rect 11778 5803 11844 5806
<< nmos >>
rect 9480 6716 9536 7516
rect 9770 5916 9826 7516
rect 10372 5916 10428 7516
rect 10532 5916 10588 7516
rect 10820 5916 10876 7516
rect 10980 5916 11036 7516
rect 11268 5916 11324 7516
rect 11428 5916 11484 7516
rect 11588 5916 11644 7516
rect 11748 5916 11804 7516
<< pmos >>
rect 2218 8088 5538 9468
rect 5642 8088 8962 9468
rect 9480 9116 9536 9516
rect 2218 6638 5538 8018
rect 5642 6638 8962 8018
rect 9480 7932 9536 8732
rect 10052 7916 10108 9516
rect 10212 7916 10268 9516
rect 10372 7916 10428 9516
rect 10532 7916 10588 9516
rect 14462 8104 16862 10104
rect 14462 6026 16862 8026
<< mvnmos >>
rect 10970 7884 11150 9484
rect 11254 7884 11434 9484
rect 11538 7884 11718 9484
rect 11822 7884 12002 9484
rect 12106 7884 12286 9484
<< ndiff >>
rect 9392 7503 9480 7516
rect 9392 6729 9405 7503
rect 9451 6729 9480 7503
rect 9392 6716 9480 6729
rect 9536 7503 9624 7516
rect 9536 6729 9565 7503
rect 9611 6729 9624 7503
rect 9536 6716 9624 6729
rect 9682 7503 9770 7516
rect 9682 5929 9695 7503
rect 9741 5929 9770 7503
rect 9682 5916 9770 5929
rect 9826 7503 9914 7516
rect 9826 5929 9855 7503
rect 9901 5929 9914 7503
rect 10284 7503 10372 7516
rect 9826 5916 9914 5929
rect 10284 5929 10297 7503
rect 10343 5929 10372 7503
rect 10284 5916 10372 5929
rect 10428 7503 10532 7516
rect 10428 5929 10457 7503
rect 10503 5929 10532 7503
rect 10428 5916 10532 5929
rect 10588 7503 10676 7516
rect 10588 5929 10617 7503
rect 10663 5929 10676 7503
rect 10588 5916 10676 5929
rect 10732 7503 10820 7516
rect 10732 5929 10745 7503
rect 10791 5929 10820 7503
rect 10732 5916 10820 5929
rect 10876 7503 10980 7516
rect 10876 5929 10905 7503
rect 10951 5929 10980 7503
rect 10876 5916 10980 5929
rect 11036 7503 11124 7516
rect 11036 5929 11065 7503
rect 11111 5929 11124 7503
rect 11036 5916 11124 5929
rect 11180 7503 11268 7516
rect 11180 5929 11193 7503
rect 11239 5929 11268 7503
rect 11180 5916 11268 5929
rect 11324 7503 11428 7516
rect 11324 5929 11353 7503
rect 11399 5929 11428 7503
rect 11324 5916 11428 5929
rect 11484 7503 11588 7516
rect 11484 5929 11513 7503
rect 11559 5929 11588 7503
rect 11484 5916 11588 5929
rect 11644 7503 11748 7516
rect 11644 5929 11673 7503
rect 11719 5929 11748 7503
rect 11644 5916 11748 5929
rect 11804 7503 11892 7516
rect 11804 5929 11833 7503
rect 11879 5929 11892 7503
rect 11804 5916 11892 5929
<< pdiff >>
rect 14374 10091 14462 10104
rect 2130 9455 2218 9468
rect 2130 8101 2143 9455
rect 2189 8101 2218 9455
rect 2130 8088 2218 8101
rect 5538 9455 5642 9468
rect 5538 8101 5567 9455
rect 5613 8101 5642 9455
rect 5538 8088 5642 8101
rect 8962 9455 9050 9468
rect 8962 8101 8991 9455
rect 9037 8101 9050 9455
rect 9392 9503 9480 9516
rect 9392 9129 9405 9503
rect 9451 9129 9480 9503
rect 9392 9116 9480 9129
rect 9536 9503 9624 9516
rect 9536 9129 9565 9503
rect 9611 9129 9624 9503
rect 9964 9503 10052 9516
rect 9536 9116 9624 9129
rect 8962 8088 9050 8101
rect 9392 8719 9480 8732
rect 2130 8005 2218 8018
rect 2130 6651 2143 8005
rect 2189 6651 2218 8005
rect 2130 6638 2218 6651
rect 5538 8005 5642 8018
rect 5538 6651 5567 8005
rect 5613 6651 5642 8005
rect 5538 6638 5642 6651
rect 8962 8005 9050 8018
rect 8962 6651 8991 8005
rect 9037 6651 9050 8005
rect 9392 7945 9405 8719
rect 9451 7945 9480 8719
rect 9392 7932 9480 7945
rect 9536 8719 9624 8732
rect 9536 7945 9565 8719
rect 9611 7945 9624 8719
rect 9536 7932 9624 7945
rect 9964 7929 9977 9503
rect 10023 7929 10052 9503
rect 9964 7916 10052 7929
rect 10108 9503 10212 9516
rect 10108 7929 10137 9503
rect 10183 7929 10212 9503
rect 10108 7916 10212 7929
rect 10268 9503 10372 9516
rect 10268 7929 10297 9503
rect 10343 7929 10372 9503
rect 10268 7916 10372 7929
rect 10428 9503 10532 9516
rect 10428 7929 10457 9503
rect 10503 7929 10532 9503
rect 10428 7916 10532 7929
rect 10588 9503 10676 9516
rect 10588 7929 10617 9503
rect 10663 7929 10676 9503
rect 10588 7916 10676 7929
rect 14374 8117 14387 10091
rect 14433 8117 14462 10091
rect 14374 8104 14462 8117
rect 16862 10091 16950 10104
rect 16862 8117 16891 10091
rect 16937 8117 16950 10091
rect 16862 8104 16950 8117
rect 14374 8013 14462 8026
rect 8962 6638 9050 6651
rect 14374 6039 14387 8013
rect 14433 6039 14462 8013
rect 14374 6026 14462 6039
rect 16862 8013 16950 8026
rect 16862 6039 16891 8013
rect 16937 6039 16950 8013
rect 16862 6026 16950 6039
<< mvndiff >>
rect 10882 9471 10970 9484
rect 10882 7897 10895 9471
rect 10941 7897 10970 9471
rect 10882 7884 10970 7897
rect 11150 9471 11254 9484
rect 11150 7897 11179 9471
rect 11225 7897 11254 9471
rect 11150 7884 11254 7897
rect 11434 9471 11538 9484
rect 11434 7897 11463 9471
rect 11509 7897 11538 9471
rect 11434 7884 11538 7897
rect 11718 9471 11822 9484
rect 11718 7897 11747 9471
rect 11793 7897 11822 9471
rect 11718 7884 11822 7897
rect 12002 9471 12106 9484
rect 12002 7897 12031 9471
rect 12077 7897 12106 9471
rect 12002 7884 12106 7897
rect 12286 9471 12374 9484
rect 12286 7897 12315 9471
rect 12361 7897 12374 9471
rect 12286 7884 12374 7897
<< ndiffc >>
rect 9405 6729 9451 7503
rect 9565 6729 9611 7503
rect 9695 5929 9741 7503
rect 9855 5929 9901 7503
rect 10297 5929 10343 7503
rect 10457 5929 10503 7503
rect 10617 5929 10663 7503
rect 10745 5929 10791 7503
rect 10905 5929 10951 7503
rect 11065 5929 11111 7503
rect 11193 5929 11239 7503
rect 11353 5929 11399 7503
rect 11513 5929 11559 7503
rect 11673 5929 11719 7503
rect 11833 5929 11879 7503
<< pdiffc >>
rect 2143 8101 2189 9455
rect 5567 8101 5613 9455
rect 8991 8101 9037 9455
rect 9405 9129 9451 9503
rect 9565 9129 9611 9503
rect 2143 6651 2189 8005
rect 5567 6651 5613 8005
rect 8991 6651 9037 8005
rect 9405 7945 9451 8719
rect 9565 7945 9611 8719
rect 9977 7929 10023 9503
rect 10137 7929 10183 9503
rect 10297 7929 10343 9503
rect 10457 7929 10503 9503
rect 10617 7929 10663 9503
rect 14387 8117 14433 10091
rect 16891 8117 16937 10091
rect 14387 6039 14433 8013
rect 16891 6039 16937 8013
<< mvndiffc >>
rect 10895 7897 10941 9471
rect 11179 7897 11225 9471
rect 11463 7897 11509 9471
rect 11747 7897 11793 9471
rect 12031 7897 12077 9471
rect 12315 7897 12361 9471
<< psubdiff >>
rect 14028 7653 14128 7673
rect 14028 7592 14054 7653
rect 14114 7592 14128 7653
rect 14028 7573 14128 7592
rect 10065 7526 10165 7552
rect 10065 7480 10094 7526
rect 10140 7480 10165 7526
rect 10065 7452 10165 7480
rect 10067 6966 10167 6994
rect 10067 6920 10094 6966
rect 10140 6920 10167 6966
rect 10067 6894 10167 6920
rect 10067 5949 10167 5977
rect 10067 5903 10093 5949
rect 10139 5903 10167 5949
rect 14025 5960 14134 5985
rect 10067 5877 10167 5903
rect 14025 5900 14045 5960
rect 14114 5900 14134 5960
rect 14025 5885 14134 5900
<< nsubdiff >>
rect 9160 9503 9260 9530
rect 9160 9457 9187 9503
rect 9233 9457 9260 9503
rect 9160 9430 9260 9457
rect 9760 9503 9860 9530
rect 9760 9457 9787 9503
rect 9833 9457 9860 9503
rect 9760 9430 9860 9457
rect 9338 7837 9438 7864
rect 9338 7788 9366 7837
rect 9415 7788 9438 7837
rect 9338 7764 9438 7788
rect 13644 8554 13744 8576
rect 13644 8494 13663 8554
rect 13730 8494 13744 8554
rect 13644 8476 13744 8494
rect 12106 6804 12206 6829
rect 12106 6756 12129 6804
rect 12183 6756 12206 6804
rect 12106 6729 12206 6756
rect 14316 5944 14416 5970
rect 14316 5898 14341 5944
rect 14387 5898 14416 5944
rect 14316 5872 14416 5898
<< psubdiffcont >>
rect 14054 7592 14114 7653
rect 10094 7480 10140 7526
rect 10094 6920 10140 6966
rect 10093 5903 10139 5949
rect 14045 5900 14114 5960
<< nsubdiffcont >>
rect 9187 9457 9233 9503
rect 9787 9457 9833 9503
rect 9366 7788 9415 7837
rect 13663 8494 13730 8554
rect 12129 6756 12183 6804
rect 14341 5898 14387 5944
<< polysilicon >>
rect 14462 10183 16862 10196
rect 14462 10137 14475 10183
rect 16849 10137 16862 10183
rect 14462 10104 16862 10137
rect 11650 9730 11930 9750
rect 11650 9620 11690 9730
rect 11910 9620 11930 9730
rect 11650 9590 11930 9620
rect 2218 9547 8962 9560
rect 2218 9501 2231 9547
rect 5525 9502 5655 9547
rect 5525 9501 5538 9502
rect 2218 9468 5538 9501
rect 5642 9501 5655 9502
rect 8949 9501 8962 9547
rect 5642 9468 8962 9501
rect 9480 9516 9536 9560
rect 10052 9516 10108 9560
rect 10212 9516 10268 9560
rect 10372 9516 10428 9560
rect 10532 9516 10588 9560
rect 10970 9550 12286 9590
rect 9480 9069 9536 9116
rect 9480 9030 9578 9069
rect 9498 8989 9578 9030
rect 9480 8732 9536 8776
rect 2218 8018 5538 8088
rect 5642 8018 8962 8088
rect 9480 7516 9536 7932
rect 10970 9484 11150 9550
rect 11254 9484 11434 9550
rect 11538 9484 11718 9550
rect 11822 9484 12002 9550
rect 12106 9484 12286 9550
rect 10052 7872 10108 7916
rect 10212 7872 10268 7916
rect 10372 7872 10428 7916
rect 10532 7872 10588 7916
rect 14462 8026 16862 8104
rect 10052 7837 10588 7872
rect 10970 7840 11150 7884
rect 11254 7840 11434 7884
rect 11538 7840 11718 7884
rect 11822 7840 12002 7884
rect 12106 7840 12286 7884
rect 10052 7791 10069 7837
rect 10115 7836 10588 7837
rect 10115 7791 10132 7836
rect 10052 7774 10132 7791
rect 10440 7637 10520 7654
rect 10440 7596 10457 7637
rect 10372 7591 10457 7596
rect 10503 7596 10520 7637
rect 10503 7591 10588 7596
rect 10372 7560 10588 7591
rect 9770 7516 9826 7560
rect 9480 6672 9536 6716
rect 9468 6655 9548 6672
rect 2218 6605 5538 6638
rect 2218 6559 2231 6605
rect 5525 6604 5538 6605
rect 5642 6605 8962 6638
rect 5642 6604 5655 6605
rect 5525 6559 5655 6604
rect 8949 6559 8962 6605
rect 9468 6609 9485 6655
rect 9531 6609 9548 6655
rect 9468 6592 9548 6609
rect 2218 6546 8962 6559
rect 10372 7516 10428 7560
rect 10532 7516 10588 7560
rect 10820 7516 10876 7560
rect 10980 7516 11036 7560
rect 11268 7516 11324 7560
rect 11428 7516 11484 7560
rect 11588 7516 11644 7560
rect 11748 7516 11804 7560
rect 9770 5872 9826 5916
rect 14462 5993 16862 6026
rect 10372 5872 10428 5916
rect 10532 5872 10588 5916
rect 10820 5872 10876 5916
rect 10980 5872 11036 5916
rect 11268 5872 11324 5916
rect 11428 5872 11484 5916
rect 11588 5872 11644 5916
rect 11748 5872 11804 5916
rect 14462 5947 14475 5993
rect 16849 5947 16862 5993
rect 14462 5934 16862 5947
rect 9758 5855 9838 5872
rect 9758 5809 9776 5855
rect 9822 5809 9838 5855
rect 10820 5869 11804 5872
rect 10820 5852 11844 5869
rect 10820 5836 11781 5852
rect 9758 5792 9838 5809
rect 11764 5806 11781 5836
rect 11827 5806 11844 5852
rect 11764 5790 11844 5806
<< polycontact >>
rect 14475 10137 16849 10183
rect 11690 9620 11910 9730
rect 2231 9501 5525 9547
rect 5655 9501 8949 9547
rect 10069 7791 10115 7837
rect 10457 7591 10503 7637
rect 2231 6559 5525 6605
rect 5655 6559 8949 6605
rect 9485 6609 9531 6655
rect 14475 5947 16849 5993
rect 9776 5809 9822 5855
rect 11781 5806 11827 5852
<< metal1 >>
rect 1713 10497 17738 10672
rect 2220 9501 2231 9547
rect 5525 9501 5536 9547
rect 5644 9501 5655 9547
rect 8949 9501 8960 9547
rect 9172 9506 9248 9518
rect 2143 9455 2189 9466
rect 2142 8665 2143 8885
rect 5567 9455 5613 9466
rect 2189 8665 5567 8885
rect 2143 8005 2189 8101
rect 8991 9455 9037 9466
rect 8976 9440 8991 9452
rect 9172 9454 9184 9506
rect 9236 9454 9248 9506
rect 9037 9440 9052 9452
rect 9172 9442 9248 9454
rect 9405 9503 9451 10497
rect 11650 9730 11930 10497
rect 11650 9620 11690 9730
rect 11910 9620 11930 9730
rect 11650 9600 11930 9620
rect 8976 9388 8988 9440
rect 9040 9388 9052 9440
rect 8976 9376 8991 9388
rect 5613 8665 8991 8885
rect 5567 8005 5613 8101
rect 2189 7145 5567 7365
rect 2143 6640 2189 6651
rect 9037 9376 9052 9388
rect 8991 8005 9037 8101
rect 5613 7145 8991 7365
rect 5567 6640 5613 6651
rect 9550 9503 9626 9514
rect 9550 9502 9565 9503
rect 9611 9502 9626 9503
rect 9550 9450 9562 9502
rect 9614 9450 9626 9502
rect 9550 9446 9565 9450
rect 9405 8719 9451 9129
rect 9611 9446 9626 9450
rect 9772 9506 9848 9518
rect 9772 9454 9784 9506
rect 9836 9454 9848 9506
rect 9772 9442 9848 9454
rect 9962 9503 10038 9514
rect 9962 9502 9977 9503
rect 10023 9502 10038 9503
rect 9962 9450 9974 9502
rect 10026 9450 10038 9502
rect 9962 9446 9977 9450
rect 9565 9118 9611 9129
rect 9498 9055 9578 9069
rect 9498 9003 9512 9055
rect 9564 9003 9578 9055
rect 9498 8989 9578 9003
rect 9405 7864 9451 7945
rect 9338 7837 9451 7864
rect 9338 7788 9366 7837
rect 9415 7788 9451 7837
rect 9338 7764 9451 7788
rect 9565 8719 9611 8730
rect 9565 7837 9611 7945
rect 10023 9446 10038 9450
rect 10137 9503 10183 9514
rect 10122 9053 10137 9065
rect 10282 9503 10358 9514
rect 10282 9502 10297 9503
rect 10343 9502 10358 9503
rect 10282 9450 10294 9502
rect 10346 9450 10358 9502
rect 10282 9446 10297 9450
rect 10183 9053 10198 9065
rect 10122 9001 10134 9053
rect 10186 9001 10198 9053
rect 10122 8989 10137 9001
rect 10122 8570 10137 8582
rect 10183 8989 10198 9001
rect 10183 8570 10198 8582
rect 10122 8518 10134 8570
rect 10186 8518 10198 8570
rect 10122 8506 10137 8518
rect 9977 7918 10023 7929
rect 10183 8506 10198 8518
rect 10137 7918 10183 7929
rect 10343 9446 10358 9450
rect 10457 9503 10503 9514
rect 10442 9053 10457 9065
rect 10602 9503 10678 9514
rect 10602 9502 10617 9503
rect 10663 9502 10678 9503
rect 10602 9450 10614 9502
rect 10666 9450 10678 9502
rect 10602 9446 10617 9450
rect 10503 9053 10518 9065
rect 10442 9001 10454 9053
rect 10506 9001 10518 9053
rect 10442 8989 10457 9001
rect 10442 8570 10457 8582
rect 10503 8989 10518 9001
rect 10503 8570 10518 8582
rect 10442 8518 10454 8570
rect 10506 8518 10518 8570
rect 10442 8506 10457 8518
rect 10297 7918 10343 7929
rect 10503 8506 10518 8518
rect 10457 7916 10503 7929
rect 10663 9446 10678 9450
rect 10880 9471 10956 9482
rect 10880 9470 10895 9471
rect 10941 9470 10956 9471
rect 10880 9418 10892 9470
rect 10944 9418 10956 9470
rect 10880 9414 10895 9418
rect 10880 8570 10895 8582
rect 10941 9414 10956 9418
rect 11179 9471 11225 9482
rect 10941 8570 10956 8582
rect 10880 8518 10892 8570
rect 10944 8518 10956 8570
rect 10880 8506 10895 8518
rect 10617 7918 10663 7929
rect 10941 8506 10956 8518
rect 10895 7886 10941 7897
rect 11164 7950 11179 7954
rect 11448 9471 11524 9482
rect 11448 9470 11463 9471
rect 11509 9470 11524 9471
rect 11448 9418 11460 9470
rect 11512 9418 11524 9470
rect 11448 9414 11463 9418
rect 11448 8570 11463 8582
rect 11509 9414 11524 9418
rect 11747 9471 11793 9482
rect 11509 8570 11524 8582
rect 11448 8518 11460 8570
rect 11512 8518 11524 8570
rect 11448 8506 11463 8518
rect 11225 7950 11240 7954
rect 11164 7898 11176 7950
rect 11228 7898 11240 7950
rect 11164 7897 11179 7898
rect 11225 7897 11240 7898
rect 11164 7886 11240 7897
rect 11509 8506 11524 8518
rect 11463 7886 11509 7897
rect 11732 7950 11747 7954
rect 12016 9471 12092 9482
rect 12016 9470 12031 9471
rect 12077 9470 12092 9471
rect 12016 9418 12028 9470
rect 12080 9418 12092 9470
rect 12016 9414 12031 9418
rect 12016 8570 12031 8582
rect 12077 9414 12092 9418
rect 12315 9471 12361 9482
rect 12077 8570 12092 8582
rect 12016 8518 12028 8570
rect 12080 8518 12092 8570
rect 12016 8506 12031 8518
rect 11793 7950 11808 7954
rect 11732 7898 11744 7950
rect 11796 7898 11808 7950
rect 11732 7897 11747 7898
rect 11793 7897 11808 7898
rect 11732 7886 11808 7897
rect 12077 8506 12092 8518
rect 12031 7886 12077 7897
rect 13644 8586 13744 10497
rect 14464 10137 14475 10183
rect 16849 10137 16937 10183
rect 14387 10091 14433 10102
rect 13700 8554 13767 8586
rect 13730 8494 13767 8554
rect 13700 8466 13767 8494
rect 12361 8090 12654 8172
rect 16891 10091 16937 10137
rect 16876 9470 16891 9482
rect 16937 9470 16952 9482
rect 16876 9418 16888 9470
rect 16940 9418 16952 9470
rect 16876 9414 16891 9418
rect 14387 8013 14433 8117
rect 12315 7886 12361 7897
rect 12838 7941 12914 7954
rect 12838 7889 12850 7941
rect 12902 7889 12914 7941
rect 12838 7877 12914 7889
rect 10052 7837 10132 7854
rect 9565 7791 10069 7837
rect 10115 7791 10132 7837
rect 9565 7514 9611 7791
rect 10052 7774 10132 7791
rect 14154 7682 14205 7683
rect 10440 7640 10520 7654
rect 14080 7653 14205 7682
rect 10440 7588 10454 7640
rect 10506 7588 10520 7640
rect 14114 7592 14205 7653
rect 10440 7574 10520 7588
rect 14080 7562 14205 7592
rect 10093 7526 10140 7552
rect 8991 6640 9037 6651
rect 9374 7503 9466 7514
rect 9374 7502 9405 7503
rect 9451 7502 9466 7503
rect 9374 7450 9402 7502
rect 9454 7450 9466 7502
rect 9374 6729 9405 7450
rect 9451 7446 9466 7450
rect 9565 7503 9741 7514
rect 9374 6718 9451 6729
rect 9611 7422 9695 7503
rect 9565 6718 9611 6729
rect 2220 6559 2231 6605
rect 5525 6559 5536 6605
rect 5644 6559 5655 6605
rect 8949 6594 8960 6605
rect 9374 6594 9420 6718
rect 8949 6559 9420 6594
rect 9468 6655 9548 6672
rect 9468 6609 9485 6655
rect 9531 6609 9548 6655
rect 9468 6592 9548 6609
rect 8915 6548 9420 6559
rect 9485 6347 9532 6592
rect 9471 6343 9547 6347
rect 9471 6291 9483 6343
rect 9535 6291 9547 6343
rect 9471 6287 9547 6291
rect 9840 7503 9916 7514
rect 9840 7502 9855 7503
rect 9901 7502 9916 7503
rect 9840 7450 9852 7502
rect 9904 7450 9916 7502
rect 9840 7446 9855 7450
rect 9695 5918 9741 5929
rect 9901 7446 9916 7450
rect 10093 7480 10094 7526
rect 10093 6966 10140 7480
rect 10093 6920 10094 6966
rect 10093 5977 10140 6920
rect 10297 7503 10343 7514
rect 10282 5982 10297 5986
rect 10442 7503 10518 7514
rect 10442 7502 10457 7503
rect 10503 7502 10518 7503
rect 10442 7450 10454 7502
rect 10506 7450 10518 7502
rect 10442 7446 10457 7450
rect 10343 5982 10358 5986
rect 9855 5918 9901 5929
rect 10067 5949 10167 5977
rect 10067 5903 10093 5949
rect 10139 5903 10167 5949
rect 10282 5930 10294 5982
rect 10346 5930 10358 5982
rect 10282 5929 10297 5930
rect 10343 5929 10358 5930
rect 10282 5918 10358 5929
rect 10503 7446 10518 7450
rect 10617 7503 10663 7514
rect 10457 5918 10503 5929
rect 10602 5982 10617 5986
rect 10730 7503 10806 7514
rect 10730 7502 10745 7503
rect 10791 7502 10806 7503
rect 10730 7450 10742 7502
rect 10794 7450 10806 7502
rect 10730 7446 10745 7450
rect 10663 5982 10678 5986
rect 10602 5930 10614 5982
rect 10666 5930 10678 5982
rect 10602 5929 10617 5930
rect 10663 5929 10678 5930
rect 10602 5918 10678 5929
rect 10791 7446 10806 7450
rect 10905 7503 10951 7514
rect 10745 5918 10791 5929
rect 10890 5982 10905 5986
rect 11048 7503 11124 7514
rect 11048 7502 11065 7503
rect 11111 7502 11124 7503
rect 11048 7450 11060 7502
rect 11112 7450 11124 7502
rect 11048 7446 11065 7450
rect 10951 5982 10966 5986
rect 10890 5930 10902 5982
rect 10954 5930 10966 5982
rect 10890 5929 10905 5930
rect 10951 5929 10966 5930
rect 10890 5918 10966 5929
rect 11111 7446 11124 7450
rect 11180 7503 11256 7514
rect 11180 7502 11193 7503
rect 11239 7502 11256 7503
rect 11180 7450 11192 7502
rect 11244 7450 11256 7502
rect 11180 7446 11193 7450
rect 11065 5918 11111 5929
rect 11239 7446 11256 7450
rect 11353 7503 11399 7514
rect 11193 5918 11239 5929
rect 11338 5982 11353 5986
rect 11498 7503 11574 7514
rect 11498 7502 11513 7503
rect 11559 7502 11574 7503
rect 11498 7450 11510 7502
rect 11562 7450 11574 7502
rect 11498 7446 11513 7450
rect 11399 5982 11414 5986
rect 11338 5930 11350 5982
rect 11402 5930 11414 5982
rect 11338 5929 11353 5930
rect 11399 5929 11414 5930
rect 11338 5918 11414 5929
rect 11559 7446 11574 7450
rect 11673 7503 11719 7514
rect 11513 5918 11559 5929
rect 11658 5982 11673 5986
rect 11818 7503 11894 7514
rect 11818 7502 11833 7503
rect 11879 7502 11894 7503
rect 11818 7450 11830 7502
rect 11882 7450 11894 7502
rect 11818 7446 11833 7450
rect 11719 5982 11734 5986
rect 11658 5930 11670 5982
rect 11722 5930 11734 5982
rect 11658 5929 11673 5930
rect 11719 5929 11734 5930
rect 11658 5918 11734 5929
rect 11879 7446 11894 7450
rect 12978 7147 13054 7315
rect 12190 6348 12916 6358
rect 12190 6296 12208 6348
rect 12260 6296 12916 6348
rect 12190 6287 12916 6296
rect 12322 6133 12398 6181
rect 12322 6081 12334 6133
rect 12386 6081 12398 6133
rect 12322 6069 12398 6081
rect 14154 5994 14205 7562
rect 14079 5960 14205 5994
rect 14341 6039 14387 6169
rect 14341 6028 14433 6039
rect 16937 9414 16952 9418
rect 16891 8013 16937 8117
rect 14341 5970 14387 6028
rect 16891 5993 16937 6039
rect 11833 5918 11879 5929
rect 11353 5916 11399 5918
rect 10067 5877 10167 5903
rect 14114 5900 14205 5960
rect 9758 5855 9838 5872
rect 9758 5809 9776 5855
rect 9822 5809 9838 5855
rect 9758 5792 9838 5809
rect 9776 5734 9822 5792
rect 9760 5726 9836 5734
rect 9760 5674 9773 5726
rect 9825 5674 9836 5726
rect 9760 5666 9836 5674
rect 10093 5315 10139 5877
rect 14079 5874 14205 5900
rect 11284 5853 11360 5862
rect 11284 5801 11296 5853
rect 11348 5801 11360 5853
rect 11284 5790 11360 5801
rect 11764 5855 11844 5869
rect 11764 5803 11778 5855
rect 11830 5803 11844 5855
rect 11764 5790 11844 5803
rect 11299 5315 11345 5790
rect 14097 5315 14205 5874
rect 14316 5944 14398 5970
rect 14464 5947 14475 5993
rect 16849 5947 16937 5993
rect 14316 5898 14341 5944
rect 14387 5898 14398 5944
rect 14316 5872 14398 5898
rect 14341 5734 14387 5872
rect 14326 5726 14402 5734
rect 14326 5674 14338 5726
rect 14390 5674 14402 5726
rect 14326 5666 14402 5674
rect 1597 5140 17622 5315
<< via1 >>
rect 9184 9503 9236 9506
rect 9184 9457 9187 9503
rect 9187 9457 9233 9503
rect 9233 9457 9236 9503
rect 9184 9454 9236 9457
rect 8988 9388 8991 9440
rect 8991 9388 9037 9440
rect 9037 9388 9040 9440
rect 9562 9450 9565 9502
rect 9565 9450 9611 9502
rect 9611 9450 9614 9502
rect 9784 9503 9836 9506
rect 9784 9457 9787 9503
rect 9787 9457 9833 9503
rect 9833 9457 9836 9503
rect 9784 9454 9836 9457
rect 9974 9450 9977 9502
rect 9977 9450 10023 9502
rect 10023 9450 10026 9502
rect 9512 9003 9564 9055
rect 10294 9450 10297 9502
rect 10297 9450 10343 9502
rect 10343 9450 10346 9502
rect 10134 9001 10137 9053
rect 10137 9001 10183 9053
rect 10183 9001 10186 9053
rect 10134 8518 10137 8570
rect 10137 8518 10183 8570
rect 10183 8518 10186 8570
rect 10614 9450 10617 9502
rect 10617 9450 10663 9502
rect 10663 9450 10666 9502
rect 10454 9001 10457 9053
rect 10457 9001 10503 9053
rect 10503 9001 10506 9053
rect 10454 8518 10457 8570
rect 10457 8518 10503 8570
rect 10503 8518 10506 8570
rect 10892 9418 10895 9470
rect 10895 9418 10941 9470
rect 10941 9418 10944 9470
rect 10892 8518 10895 8570
rect 10895 8518 10941 8570
rect 10941 8518 10944 8570
rect 11460 9418 11463 9470
rect 11463 9418 11509 9470
rect 11509 9418 11512 9470
rect 11460 8518 11463 8570
rect 11463 8518 11509 8570
rect 11509 8518 11512 8570
rect 11176 7898 11179 7950
rect 11179 7898 11225 7950
rect 11225 7898 11228 7950
rect 12028 9418 12031 9470
rect 12031 9418 12077 9470
rect 12077 9418 12080 9470
rect 12028 8518 12031 8570
rect 12031 8518 12077 8570
rect 12077 8518 12080 8570
rect 11744 7898 11747 7950
rect 11747 7898 11793 7950
rect 11793 7898 11796 7950
rect 13672 8498 13724 8550
rect 16888 9418 16891 9470
rect 16891 9418 16937 9470
rect 16937 9418 16940 9470
rect 12850 7889 12902 7941
rect 10454 7637 10506 7640
rect 10454 7591 10457 7637
rect 10457 7591 10503 7637
rect 10503 7591 10506 7637
rect 10454 7588 10506 7591
rect 9402 7450 9405 7502
rect 9405 7450 9451 7502
rect 9451 7450 9454 7502
rect 9483 6291 9535 6343
rect 9852 7450 9855 7502
rect 9855 7450 9901 7502
rect 9901 7450 9904 7502
rect 10454 7450 10457 7502
rect 10457 7450 10503 7502
rect 10503 7450 10506 7502
rect 10294 5930 10297 5982
rect 10297 5930 10343 5982
rect 10343 5930 10346 5982
rect 10742 7450 10745 7502
rect 10745 7450 10791 7502
rect 10791 7450 10794 7502
rect 10614 5930 10617 5982
rect 10617 5930 10663 5982
rect 10663 5930 10666 5982
rect 11060 7450 11065 7502
rect 11065 7450 11111 7502
rect 11111 7450 11112 7502
rect 10902 5930 10905 5982
rect 10905 5930 10951 5982
rect 10951 5930 10954 5982
rect 11192 7450 11193 7502
rect 11193 7450 11239 7502
rect 11239 7450 11244 7502
rect 11510 7450 11513 7502
rect 11513 7450 11559 7502
rect 11559 7450 11562 7502
rect 11350 5930 11353 5982
rect 11353 5930 11399 5982
rect 11399 5930 11402 5982
rect 11830 7450 11833 7502
rect 11833 7450 11879 7502
rect 11879 7450 11882 7502
rect 11670 5930 11673 5982
rect 11673 5930 11719 5982
rect 11719 5930 11722 5982
rect 12850 7207 12902 7259
rect 13671 6749 13723 6801
rect 12208 6296 12260 6348
rect 12334 6081 12386 6133
rect 9773 5674 9825 5726
rect 11296 5801 11348 5853
rect 11778 5852 11830 5855
rect 11778 5806 11781 5852
rect 11781 5806 11827 5852
rect 11827 5806 11830 5852
rect 11778 5803 11830 5806
rect 14338 5674 14390 5726
<< metal2 >>
rect 8976 9506 10678 9514
rect 8976 9454 9184 9506
rect 9236 9502 9784 9506
rect 9236 9454 9562 9502
rect 8976 9450 9562 9454
rect 9614 9454 9784 9502
rect 9836 9502 10678 9506
rect 9836 9454 9974 9502
rect 9614 9450 9974 9454
rect 10026 9450 10294 9502
rect 10346 9450 10614 9502
rect 10666 9450 10678 9502
rect 8976 9446 10678 9450
rect 10880 9470 16952 9482
rect 8976 9440 9052 9446
rect 8976 9388 8988 9440
rect 9040 9388 9052 9440
rect 10880 9418 10892 9470
rect 10944 9418 11460 9470
rect 11512 9418 12028 9470
rect 12080 9418 16888 9470
rect 16940 9418 16952 9470
rect 10880 9414 16952 9418
rect 8976 9376 9052 9388
rect 9498 9065 9578 9069
rect 9498 9055 10518 9065
rect 9498 9003 9512 9055
rect 9564 9053 10518 9055
rect 9564 9003 10134 9053
rect 9498 9001 10134 9003
rect 10186 9001 10454 9053
rect 10506 9001 10518 9053
rect 9498 8989 10518 9001
rect 10122 8570 12092 8582
rect 10122 8518 10134 8570
rect 10186 8518 10454 8570
rect 10506 8518 10892 8570
rect 10944 8518 11460 8570
rect 11512 8518 12028 8570
rect 12080 8518 12092 8570
rect 10122 8506 12092 8518
rect 13644 8550 13744 8586
rect 10440 7640 10520 8506
rect 13644 8498 13672 8550
rect 13724 8498 13744 8550
rect 11164 7950 11808 7954
rect 11164 7898 11176 7950
rect 11228 7898 11744 7950
rect 11796 7898 11808 7950
rect 11164 7886 11808 7898
rect 12838 7941 12914 7954
rect 12838 7889 12850 7941
rect 12902 7889 12914 7941
rect 10440 7588 10454 7640
rect 10506 7588 10520 7640
rect 10440 7574 10520 7588
rect 11510 7514 11613 7886
rect 9390 7502 11124 7514
rect 9390 7450 9402 7502
rect 9454 7450 9852 7502
rect 9904 7450 10454 7502
rect 10506 7450 10742 7502
rect 10794 7450 11060 7502
rect 11112 7450 11124 7502
rect 9390 7446 11124 7450
rect 11180 7502 11894 7514
rect 11180 7450 11192 7502
rect 11244 7450 11510 7502
rect 11562 7450 11830 7502
rect 11882 7450 11894 7502
rect 11180 7446 11894 7450
rect 12838 7259 12914 7889
rect 12838 7207 12850 7259
rect 12902 7207 12914 7259
rect 12838 7198 12914 7207
rect 13644 6801 13744 8498
rect 13644 6749 13671 6801
rect 13723 6749 13744 6801
rect 13644 6658 13744 6749
rect 9471 6348 12271 6358
rect 9471 6343 12208 6348
rect 9471 6291 9483 6343
rect 9535 6296 12208 6343
rect 12260 6296 12271 6348
rect 9535 6291 12271 6296
rect 9471 6287 12271 6291
rect 12322 6133 12398 6145
rect 12322 6081 12334 6133
rect 12386 6081 12398 6133
rect 10282 5982 10678 5986
rect 10282 5930 10294 5982
rect 10346 5930 10614 5982
rect 10666 5930 10678 5982
rect 10282 5917 10678 5930
rect 10890 5982 11734 5986
rect 10890 5930 10902 5982
rect 10954 5930 11350 5982
rect 11402 5930 11670 5982
rect 11722 5930 11734 5982
rect 10890 5918 11734 5930
rect 11290 5862 11353 5918
rect 12322 5872 12398 6081
rect 11844 5869 12398 5872
rect 11284 5853 11360 5862
rect 11284 5801 11296 5853
rect 11348 5801 11360 5853
rect 11284 5790 11360 5801
rect 11764 5855 12398 5869
rect 11764 5803 11778 5855
rect 11830 5806 12398 5855
rect 11830 5803 11844 5806
rect 11764 5790 11844 5803
rect 9760 5726 14402 5734
rect 9760 5674 9773 5726
rect 9825 5674 14338 5726
rect 14390 5674 14402 5726
rect 9760 5666 14402 5674
use gf180mcu_fd_sc_mcu7t5v0__inv_4  gf180mcu_fd_sc_mcu7t5v0__inv_4_0 ~/conda-gf180mcu-env/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 12580 0 1 7742
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  gf180mcu_fd_sc_mcu7t5v0__inv_8_0 ~/conda-gf180mcu-env/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 12064 0 -1 7622
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  gf180mcu_fd_sc_mcu7t5v0__inv_8_1
timestamp 1753044640
transform 1 0 12064 0 1 5934
box -86 -86 2102 870
<< labels >>
flabel metal1 2142 8665 9032 8885 1 FreeSans 3200 0 0 0 Vtop
flabel metal1 9405 9118 9451 9514 1 FreeSans 400 0 0 0 VDD
flabel nwell 9405 7932 9451 8732 1 FreeSans 400 0 0 0 VDD
flabel metal2 8976 9446 10678 9514 1 FreeSans 800 0 0 0 Vtop
flabel nwell 10052 7836 10588 7872 1 FreeSans 400 0 0 0 EN_Z_LVL_SHFT
flabel metal1 9565 7791 10069 7837 1 FreeSans 400 0 0 0 EN_Z_LVL_SHFT
flabel polysilicon 10970 9550 12002 9590 1 FreeSans 400 0 0 0 VDD
flabel pwell 9374 6718 9451 7514 1 FreeSans 400 0 0 0 Vbottom
flabel polysilicon 10820 5836 11036 5872 1 FreeSans 400 0 0 0 EN_Z
flabel polysilicon 11268 5836 11804 5872 1 FreeSans 400 0 0 0 EN_Z
flabel metal2 10890 5918 11734 5986 1 FreeSans 400 0 0 0 VSS
flabel metal2 10282 5917 10678 5986 1 FreeSans 400 0 0 0 VIN
port 3 n
flabel metal2 10518 7446 11124 7514 1 FreeSans 400 0 0 0 Vbottom
flabel metal2 9825 5666 14338 5734 1 FreeSans 800 0 0 0 VGATE
port 6 n
flabel metal1 1713 10497 17738 10672 1 FreeSans 3200 0 0 0 VDD
port 1 n
flabel metal1 1597 5140 17622 5315 1 FreeSans 3200 0 0 0 VSS
port 2 n
flabel metal1 12978 7147 13054 7315 1 FreeSans 400 0 0 0 SW_ON
port 4 n
flabel metal1 12190 6287 12916 6358 1 FreeSans 400 0 0 0 EN
port 5 n
<< end >>
