magic
tech gf180mcuD
magscale 1 10
timestamp 1757847982
<< nwell >>
rect 324 570 409 657
rect 640 570 725 657
rect 162 4 247 90
rect 481 3 566 90
<< polysilicon >>
rect 324 570 409 657
rect 640 570 725 657
rect 162 4 247 90
rect 481 3 566 90
<< metal1 >>
rect 324 644 409 657
rect 324 592 340 644
rect 396 592 409 644
rect 324 577 409 592
rect 640 644 725 657
rect 640 592 652 644
rect 708 592 725 644
rect 640 577 725 592
rect 162 74 247 84
rect 162 19 178 74
rect 237 19 247 74
rect 162 4 247 19
rect 481 71 566 83
rect 481 18 494 71
rect 555 18 566 71
rect 481 3 566 18
<< via1 >>
rect 340 592 396 644
rect 652 592 708 644
rect 178 19 237 74
rect 494 18 555 71
<< metal2 >>
rect 324 644 409 657
rect 324 592 340 644
rect 396 592 409 644
rect 324 577 409 592
rect 640 644 725 657
rect 640 592 652 644
rect 708 592 725 644
rect 640 577 725 592
rect 162 74 247 84
rect 162 19 178 74
rect 237 19 247 74
rect 162 4 247 19
rect 481 71 566 83
rect 481 18 494 71
rect 555 18 566 71
rect 481 3 566 18
use pfet_03v3_9DSAFW  pfet_03v3_9DSAFW_0
timestamp 1757847982
transform 1 0 442 0 1 330
box -442 -330 442 330
<< end >>
