magic
tech gf180mcuD
magscale 1 10
timestamp 1757817671
<< nwell >>
rect -117 653 69 654
rect -117 -107 982 653
rect -105 -108 982 -107
<< nsubdiff >>
rect -84 587 935 608
rect -84 539 41 587
rect 843 539 935 587
rect -84 526 935 539
rect -84 481 0 526
rect -84 43 -67 481
rect -13 43 0 481
rect 850 492 935 526
rect -84 0 0 43
rect 850 54 864 492
rect 918 54 935 492
rect 850 0 935 54
rect -84 -14 935 0
rect -84 -62 28 -14
rect 830 -62 935 -14
rect -84 -81 935 -62
<< nsubdiffcont >>
rect 41 539 843 587
rect -67 43 -13 481
rect 864 54 918 492
rect 28 -62 830 -14
<< polysilicon >>
rect 175 438 374 459
rect 175 385 217 438
rect 341 385 374 438
rect 175 360 374 385
rect 478 442 677 459
rect 478 390 507 442
rect 659 390 677 442
rect 478 360 677 390
<< polycontact >>
rect 217 385 341 438
rect 507 390 659 442
<< metal1 >>
rect -84 587 935 608
rect -84 539 41 587
rect 843 539 935 587
rect -84 526 935 539
rect -84 481 0 526
rect -84 43 -67 481
rect -13 43 0 481
rect 850 492 935 526
rect 179 450 371 451
rect 179 438 374 450
rect 179 385 217 438
rect 341 385 374 438
rect 179 379 374 385
rect 478 442 677 450
rect 478 390 507 442
rect 659 390 677 442
rect 478 379 677 390
rect 179 378 371 379
rect -84 0 0 43
rect 850 54 864 492
rect 918 54 935 492
rect 850 0 935 54
rect -84 -14 935 0
rect -84 -62 28 -14
rect 830 -62 935 -14
rect -84 -81 935 -62
use pfet_03v3_US4NEC  pfet_03v3_US4NEC_0
timestamp 1757723484
transform 1 0 426 0 1 230
box -426 -230 426 230
<< end >>
