magic
tech gf180mcuD
magscale 1 10
timestamp 1757235355
<< nwell >>
rect -762 -930 762 930
<< pmos >>
rect -588 -800 -532 800
rect -428 -800 -372 800
rect -268 -800 -212 800
rect -108 -800 -52 800
rect 52 -800 108 800
rect 212 -800 268 800
rect 372 -800 428 800
rect 532 -800 588 800
<< pdiff >>
rect -676 787 -588 800
rect -676 -787 -663 787
rect -617 -787 -588 787
rect -676 -800 -588 -787
rect -532 787 -428 800
rect -532 -787 -503 787
rect -457 -787 -428 787
rect -532 -800 -428 -787
rect -372 787 -268 800
rect -372 -787 -343 787
rect -297 -787 -268 787
rect -372 -800 -268 -787
rect -212 787 -108 800
rect -212 -787 -183 787
rect -137 -787 -108 787
rect -212 -800 -108 -787
rect -52 787 52 800
rect -52 -787 -23 787
rect 23 -787 52 787
rect -52 -800 52 -787
rect 108 787 212 800
rect 108 -787 137 787
rect 183 -787 212 787
rect 108 -800 212 -787
rect 268 787 372 800
rect 268 -787 297 787
rect 343 -787 372 787
rect 268 -800 372 -787
rect 428 787 532 800
rect 428 -787 457 787
rect 503 -787 532 787
rect 428 -800 532 -787
rect 588 787 676 800
rect 588 -787 617 787
rect 663 -787 676 787
rect 588 -800 676 -787
<< pdiffc >>
rect -663 -787 -617 787
rect -503 -787 -457 787
rect -343 -787 -297 787
rect -183 -787 -137 787
rect -23 -787 23 787
rect 137 -787 183 787
rect 297 -787 343 787
rect 457 -787 503 787
rect 617 -787 663 787
<< polysilicon >>
rect -588 800 -532 844
rect -428 800 -372 844
rect -268 800 -212 844
rect -108 800 -52 844
rect 52 800 108 844
rect 212 800 268 844
rect 372 800 428 844
rect 532 800 588 844
rect -588 -844 -532 -800
rect -428 -844 -372 -800
rect -268 -844 -212 -800
rect -108 -844 -52 -800
rect 52 -844 108 -800
rect 212 -844 268 -800
rect 372 -844 428 -800
rect 532 -844 588 -800
<< metal1 >>
rect -663 787 -617 798
rect -663 -798 -617 -787
rect -503 787 -457 798
rect -503 -798 -457 -787
rect -343 787 -297 798
rect -343 -798 -297 -787
rect -183 787 -137 798
rect -183 -798 -137 -787
rect -23 787 23 798
rect -23 -798 23 -787
rect 137 787 183 798
rect 137 -798 183 -787
rect 297 787 343 798
rect 297 -798 343 -787
rect 457 787 503 798
rect 457 -798 503 -787
rect 617 787 663 798
rect 617 -798 663 -787
<< properties >>
string gencell pfet_03v3
string library gf180mcu
string parameters w 8 l 0.280 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {pfet_03v3 pfet_06v0}
<< end >>
