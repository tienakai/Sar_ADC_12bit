magic
tech gf180mcuD
magscale 1 10
timestamp 1757690107
<< psubdiff >>
rect 130 260 15320 280
rect 130 209 150 260
rect 15260 209 15320 260
rect 130 190 15320 209
rect 0 130 80 150
rect 0 -32110 14 130
rect 65 -32110 80 130
rect 0 -32130 80 -32110
rect 130 -32192 15320 -32179
rect 130 -32257 150 -32192
rect 445 -32193 15320 -32192
rect 15300 -32257 15320 -32193
rect 130 -32270 15320 -32257
<< psubdiffcont >>
rect 150 209 15260 260
rect 14 -32110 65 130
rect 150 -32193 445 -32192
rect 150 -32257 15300 -32193
<< metal1 >>
rect 79 651 320 660
rect 79 590 89 651
rect 150 590 250 651
rect 311 590 320 651
rect 79 580 320 590
rect 15110 609 15452 622
rect 169 527 230 580
rect 15110 551 15128 609
rect 15201 551 15359 609
rect 15432 551 15452 609
rect 15110 540 15452 551
rect 169 280 231 527
rect 15249 280 15321 540
rect 130 275 15321 280
rect 130 261 15320 275
rect 130 209 150 261
rect 15260 209 15320 261
rect 130 190 15320 209
rect 0 130 80 150
rect 0 -32110 14 130
rect 66 -32110 80 130
rect 0 -32130 80 -32110
rect 130 -32192 15320 -32179
rect 130 -32257 150 -32192
rect 445 -32193 15320 -32192
rect 15300 -32257 15320 -32193
rect 130 -32270 15320 -32257
<< via1 >>
rect 89 590 150 651
rect 250 590 311 651
rect 15128 551 15201 609
rect 15359 551 15432 609
rect 150 260 15260 261
rect 150 209 15260 260
rect 14 -32110 65 130
rect 65 -32110 66 130
rect 150 -32257 15300 -32193
<< metal2 >>
rect 78 651 320 660
rect 78 590 89 651
rect 150 590 250 651
rect 311 590 320 651
rect 78 580 320 590
rect 15110 611 15452 622
rect 168 448 231 580
rect 15110 551 15127 611
rect 15201 551 15358 611
rect 15432 551 15452 611
rect 15110 540 15452 551
rect 15249 450 15321 540
rect 1370 440 1770 450
rect 1370 380 1380 440
rect 1440 380 1700 440
rect 1760 380 1770 440
rect 1370 270 1770 380
rect 1826 440 2226 450
rect 1826 380 1836 440
rect 1896 380 2156 440
rect 2216 380 2226 440
rect 1826 270 2226 380
rect 2282 440 2682 450
rect 2282 380 2292 440
rect 2352 380 2612 440
rect 2672 380 2682 440
rect 2282 280 2682 380
rect 2740 440 3140 450
rect 2740 380 2750 440
rect 2810 380 3070 440
rect 3130 380 3140 440
rect 2740 280 3140 380
rect 2282 270 3140 280
rect 3196 440 3596 450
rect 3196 380 3206 440
rect 3266 380 3526 440
rect 3586 380 3596 440
rect 3196 270 3596 380
rect 3652 440 4052 450
rect 3652 380 3662 440
rect 3722 380 3982 440
rect 4042 380 4052 440
rect 3652 270 4052 380
rect 4110 440 4510 450
rect 4110 380 4120 440
rect 4180 380 4440 440
rect 4500 380 4510 440
rect 4110 270 4510 380
rect 4566 440 4966 450
rect 4566 380 4576 440
rect 4636 380 4896 440
rect 4956 380 4966 440
rect 4566 270 4966 380
rect 5022 440 5422 450
rect 5022 380 5032 440
rect 5092 380 5352 440
rect 5412 380 5422 440
rect 5022 270 5422 380
rect 5480 440 5880 450
rect 5480 380 5490 440
rect 5550 380 5810 440
rect 5870 380 5880 440
rect 5480 270 5880 380
rect 5936 440 6336 450
rect 5936 380 5946 440
rect 6006 380 6266 440
rect 6326 380 6336 440
rect 5936 270 6336 380
rect 6392 440 6792 450
rect 6392 380 6402 440
rect 6462 380 6722 440
rect 6782 380 6792 440
rect 6392 270 6792 380
rect 6850 440 7250 450
rect 6850 380 6860 440
rect 6920 380 7180 440
rect 7240 380 7250 440
rect 6850 270 7250 380
rect 7306 440 7706 450
rect 7306 380 7316 440
rect 7376 380 7636 440
rect 7696 380 7706 440
rect 7306 270 7706 380
rect 7762 440 8162 450
rect 7762 380 7772 440
rect 7832 380 8092 440
rect 8152 380 8162 440
rect 7762 270 8162 380
rect 8236 440 8636 450
rect 8236 380 8246 440
rect 8306 380 8566 440
rect 8626 380 8636 440
rect 8236 270 8636 380
rect 8692 440 9092 450
rect 8692 380 8702 440
rect 8762 380 9022 440
rect 9082 380 9092 440
rect 8692 270 9092 380
rect 9150 440 9550 450
rect 9150 380 9160 440
rect 9220 380 9480 440
rect 9540 380 9550 440
rect 9150 270 9550 380
rect 9606 440 10006 450
rect 9606 380 9616 440
rect 9676 380 9936 440
rect 9996 380 10006 440
rect 9606 270 10006 380
rect 10062 440 10462 450
rect 10062 380 10072 440
rect 10132 380 10392 440
rect 10452 380 10462 440
rect 10062 280 10462 380
rect 10520 440 10920 450
rect 10520 380 10530 440
rect 10590 380 10850 440
rect 10910 380 10920 440
rect 10520 280 10920 380
rect 10062 270 10920 280
rect 10976 440 11376 450
rect 10976 380 10986 440
rect 11046 380 11306 440
rect 11366 380 11376 440
rect 10976 270 11376 380
rect 11432 440 11832 450
rect 11432 380 11442 440
rect 11502 380 11762 440
rect 11822 380 11832 440
rect 11432 270 11832 380
rect 11890 440 12290 450
rect 11890 380 11900 440
rect 11960 380 12220 440
rect 12280 380 12290 440
rect 11890 270 12290 380
rect 12346 440 12746 450
rect 12346 380 12356 440
rect 12416 380 12676 440
rect 12736 380 12746 440
rect 12346 270 12746 380
rect 12802 440 13202 450
rect 12802 380 12812 440
rect 12872 380 13132 440
rect 13192 380 13202 440
rect 12802 270 13202 380
rect 13260 440 13660 450
rect 13260 380 13270 440
rect 13330 380 13590 440
rect 13650 380 13660 440
rect 13260 270 13660 380
rect 13716 440 14116 450
rect 13716 380 13726 440
rect 13786 380 14046 440
rect 14106 380 14116 440
rect 13716 270 14116 380
rect 14172 440 14572 450
rect 14172 380 14182 440
rect 14242 380 14502 440
rect 14562 380 14572 440
rect 14172 270 14572 380
rect 14630 440 15030 450
rect 14630 380 14640 440
rect 14700 380 14960 440
rect 15020 380 15030 440
rect 14630 270 15030 380
rect 15086 440 15486 450
rect 15086 380 15096 440
rect 15156 380 15416 440
rect 15476 380 15486 440
rect 15086 270 15486 380
rect 375 269 489 270
rect 820 269 934 270
rect 1270 269 15486 270
rect 335 261 15486 269
rect 15260 209 15486 261
rect 335 199 15486 209
rect 0 130 80 150
rect 0 -52 14 130
rect 66 -42 80 130
rect 1370 90 1770 199
rect 1370 30 1380 90
rect 1440 30 1700 90
rect 1760 30 1770 90
rect 1370 20 1770 30
rect 1826 90 2226 199
rect 1826 30 1836 90
rect 1896 30 2156 90
rect 2216 30 2226 90
rect 1826 20 2226 30
rect 2282 190 3140 199
rect 2282 90 2682 190
rect 2282 30 2292 90
rect 2352 30 2612 90
rect 2672 30 2682 90
rect 2282 20 2682 30
rect 2740 90 3140 190
rect 2740 30 2750 90
rect 2810 30 3070 90
rect 3130 30 3140 90
rect 2740 20 3140 30
rect 3196 90 3596 199
rect 3196 30 3206 90
rect 3266 30 3526 90
rect 3586 30 3596 90
rect 3196 20 3596 30
rect 3652 90 4052 199
rect 3652 30 3662 90
rect 3722 30 3982 90
rect 4042 30 4052 90
rect 3652 20 4052 30
rect 4110 90 4510 199
rect 4110 30 4120 90
rect 4180 30 4440 90
rect 4500 30 4510 90
rect 4110 20 4510 30
rect 4566 90 4966 199
rect 4566 30 4576 90
rect 4636 30 4896 90
rect 4956 30 4966 90
rect 4566 20 4966 30
rect 5022 90 5422 199
rect 5022 30 5032 90
rect 5092 30 5352 90
rect 5412 30 5422 90
rect 5022 20 5422 30
rect 5480 90 5880 199
rect 5480 30 5490 90
rect 5550 30 5810 90
rect 5870 30 5880 90
rect 5480 20 5880 30
rect 5936 90 6336 199
rect 5936 30 5946 90
rect 6006 30 6266 90
rect 6326 30 6336 90
rect 5936 20 6336 30
rect 6392 90 6792 199
rect 6392 30 6402 90
rect 6462 30 6722 90
rect 6782 30 6792 90
rect 6392 20 6792 30
rect 6850 90 7250 199
rect 6850 30 6860 90
rect 6920 30 7180 90
rect 7240 30 7250 90
rect 6850 20 7250 30
rect 7306 90 7706 199
rect 7306 30 7316 90
rect 7376 30 7636 90
rect 7696 30 7706 90
rect 7306 20 7706 30
rect 7762 90 8162 199
rect 7762 30 7772 90
rect 7832 30 8092 90
rect 8152 30 8162 90
rect 7762 20 8162 30
rect 8236 90 8636 199
rect 8236 30 8246 90
rect 8306 30 8566 90
rect 8626 30 8636 90
rect 8236 20 8636 30
rect 8692 90 9092 199
rect 8692 30 8702 90
rect 8762 30 9022 90
rect 9082 30 9092 90
rect 8692 20 9092 30
rect 9150 90 9550 199
rect 9150 30 9160 90
rect 9220 30 9480 90
rect 9540 30 9550 90
rect 9150 20 9550 30
rect 9606 90 10006 199
rect 9606 30 9616 90
rect 9676 30 9936 90
rect 9996 30 10006 90
rect 9606 20 10006 30
rect 10062 190 10920 199
rect 10062 90 10462 190
rect 10062 30 10072 90
rect 10132 30 10392 90
rect 10452 30 10462 90
rect 10062 20 10462 30
rect 10520 90 10920 190
rect 10520 30 10530 90
rect 10590 30 10850 90
rect 10910 30 10920 90
rect 10520 20 10920 30
rect 10976 90 11376 199
rect 10976 30 10986 90
rect 11046 30 11306 90
rect 11366 30 11376 90
rect 10976 20 11376 30
rect 11432 90 11832 199
rect 11432 30 11442 90
rect 11502 30 11762 90
rect 11822 30 11832 90
rect 11432 20 11832 30
rect 11890 90 12290 199
rect 11890 30 11900 90
rect 11960 30 12220 90
rect 12280 30 12290 90
rect 11890 20 12290 30
rect 12346 90 12746 199
rect 12346 30 12356 90
rect 12416 30 12676 90
rect 12736 30 12746 90
rect 12346 20 12746 30
rect 12802 90 13202 199
rect 12802 30 12812 90
rect 12872 30 13132 90
rect 13192 30 13202 90
rect 12802 20 13202 30
rect 13260 90 13660 199
rect 13260 30 13270 90
rect 13330 30 13590 90
rect 13650 30 13660 90
rect 13260 20 13660 30
rect 13716 90 14116 199
rect 13716 30 13726 90
rect 13786 30 14046 90
rect 14106 30 14116 90
rect 13716 20 14116 30
rect 14172 90 14572 199
rect 14172 30 14182 90
rect 14242 30 14502 90
rect 14562 30 14572 90
rect 14172 20 14572 30
rect 14630 90 15030 199
rect 14630 30 14640 90
rect 14700 30 14960 90
rect 15020 30 15030 90
rect 14630 20 15030 30
rect 15086 90 15486 199
rect 15086 30 15096 90
rect 15156 30 15416 90
rect 15476 30 15486 90
rect 15086 20 15486 30
rect 66 -52 400 -42
rect 0 -112 10 -52
rect 70 -112 330 -52
rect 390 -112 400 -52
rect 0 -402 14 -112
rect 66 -402 400 -112
rect 0 -462 10 -402
rect 70 -462 330 -402
rect 390 -462 400 -402
rect 0 -554 14 -462
rect 66 -472 400 -462
rect 456 -52 856 -42
rect 456 -112 466 -52
rect 526 -112 786 -52
rect 846 -112 856 -52
rect 456 -222 856 -112
rect 912 -52 1312 -42
rect 912 -112 922 -52
rect 982 -112 1242 -52
rect 1302 -112 1312 -52
rect 912 -222 1312 -112
rect 1370 -52 1770 -42
rect 1370 -112 1380 -52
rect 1440 -112 1700 -52
rect 1760 -112 1770 -52
rect 1370 -222 1770 -112
rect 1826 -52 2226 -42
rect 1826 -112 1836 -52
rect 1896 -112 2156 -52
rect 2216 -112 2226 -52
rect 1826 -222 2226 -112
rect 2282 -52 2682 -42
rect 2282 -112 2292 -52
rect 2352 -112 2612 -52
rect 2672 -112 2682 -52
rect 2282 -222 2682 -112
rect 456 -223 2682 -222
rect 2740 -52 3140 -42
rect 2740 -112 2750 -52
rect 2810 -112 3070 -52
rect 3130 -112 3140 -52
rect 2740 -222 3140 -112
rect 3196 -52 3596 -42
rect 3196 -112 3206 -52
rect 3266 -112 3526 -52
rect 3586 -112 3596 -52
rect 3196 -222 3596 -112
rect 3652 -52 4052 -42
rect 3652 -112 3662 -52
rect 3722 -112 3982 -52
rect 4042 -112 4052 -52
rect 3652 -222 4052 -112
rect 4110 -52 4510 -42
rect 4110 -112 4120 -52
rect 4180 -112 4440 -52
rect 4500 -112 4510 -52
rect 4110 -222 4510 -112
rect 4566 -52 4966 -42
rect 4566 -112 4576 -52
rect 4636 -112 4896 -52
rect 4956 -112 4966 -52
rect 4566 -222 4966 -112
rect 5022 -52 5422 -42
rect 5022 -112 5032 -52
rect 5092 -112 5352 -52
rect 5412 -112 5422 -52
rect 5022 -222 5422 -112
rect 5480 -52 5880 -42
rect 5480 -112 5490 -52
rect 5550 -112 5810 -52
rect 5870 -112 5880 -52
rect 5480 -222 5880 -112
rect 5936 -52 6336 -42
rect 5936 -112 5946 -52
rect 6006 -112 6266 -52
rect 6326 -112 6336 -52
rect 5936 -222 6336 -112
rect 6392 -52 6792 -42
rect 6392 -112 6402 -52
rect 6462 -112 6722 -52
rect 6782 -112 6792 -52
rect 6392 -222 6792 -112
rect 6850 -52 7250 -42
rect 6850 -112 6860 -52
rect 6920 -112 7180 -52
rect 7240 -112 7250 -52
rect 6850 -222 7250 -112
rect 7306 -52 7706 -42
rect 7306 -112 7316 -52
rect 7376 -112 7636 -52
rect 7696 -112 7706 -52
rect 7306 -222 7706 -112
rect 7762 -52 8162 -42
rect 7762 -112 7772 -52
rect 7832 -112 8092 -52
rect 8152 -112 8162 -52
rect 7762 -222 8162 -112
rect 8236 -52 8636 -42
rect 8236 -112 8246 -52
rect 8306 -112 8566 -52
rect 8626 -112 8636 -52
rect 8236 -222 8636 -112
rect 8692 -52 9092 -42
rect 8692 -112 8702 -52
rect 8762 -112 9022 -52
rect 9082 -112 9092 -52
rect 8692 -222 9092 -112
rect 9150 -52 9550 -42
rect 9150 -112 9160 -52
rect 9220 -112 9480 -52
rect 9540 -112 9550 -52
rect 9150 -222 9550 -112
rect 9606 -52 10006 -42
rect 9606 -112 9616 -52
rect 9676 -112 9936 -52
rect 9996 -112 10006 -52
rect 9606 -222 10006 -112
rect 10062 -52 10462 -42
rect 10062 -112 10072 -52
rect 10132 -112 10392 -52
rect 10452 -112 10462 -52
rect 10062 -222 10462 -112
rect 2740 -223 10462 -222
rect 10520 -52 10920 -42
rect 10520 -112 10530 -52
rect 10590 -112 10850 -52
rect 10910 -112 10920 -52
rect 10520 -222 10920 -112
rect 10976 -52 11376 -42
rect 10976 -112 10986 -52
rect 11046 -112 11306 -52
rect 11366 -112 11376 -52
rect 10976 -222 11376 -112
rect 11432 -52 11832 -42
rect 11432 -112 11442 -52
rect 11502 -112 11762 -52
rect 11822 -112 11832 -52
rect 11432 -222 11832 -112
rect 11890 -52 12290 -42
rect 11890 -112 11900 -52
rect 11960 -112 12220 -52
rect 12280 -112 12290 -52
rect 11890 -222 12290 -112
rect 12346 -52 12746 -42
rect 12346 -112 12356 -52
rect 12416 -112 12676 -52
rect 12736 -112 12746 -52
rect 12346 -222 12746 -112
rect 12802 -52 13202 -42
rect 12802 -112 12812 -52
rect 12872 -112 13132 -52
rect 13192 -112 13202 -52
rect 12802 -222 13202 -112
rect 13260 -52 13660 -42
rect 13260 -112 13270 -52
rect 13330 -112 13590 -52
rect 13650 -112 13660 -52
rect 13260 -222 13660 -112
rect 13716 -52 14116 -42
rect 13716 -112 13726 -52
rect 13786 -112 14046 -52
rect 14106 -112 14116 -52
rect 13716 -222 14116 -112
rect 14172 -52 14572 -42
rect 14172 -112 14182 -52
rect 14242 -112 14502 -52
rect 14562 -112 14572 -52
rect 14172 -222 14572 -112
rect 14630 -52 15030 -42
rect 14630 -112 14640 -52
rect 14700 -112 14960 -52
rect 15020 -112 15030 -52
rect 14630 -222 15030 -112
rect 15086 -52 15486 -42
rect 15086 -112 15096 -52
rect 15156 -112 15416 -52
rect 15476 -112 15486 -52
rect 15086 -222 15486 -112
rect 10520 -223 15486 -222
rect 456 -293 15486 -223
rect 456 -402 856 -293
rect 456 -462 466 -402
rect 526 -462 786 -402
rect 846 -462 856 -402
rect 456 -472 856 -462
rect 912 -402 1312 -293
rect 912 -462 922 -402
rect 982 -462 1242 -402
rect 1302 -462 1312 -402
rect 912 -472 1312 -462
rect 1370 -402 1770 -293
rect 1370 -462 1380 -402
rect 1440 -462 1700 -402
rect 1760 -462 1770 -402
rect 1370 -472 1770 -462
rect 1826 -402 2226 -293
rect 1826 -462 1836 -402
rect 1896 -462 2156 -402
rect 2216 -462 2226 -402
rect 1826 -472 2226 -462
rect 2282 -402 2682 -293
rect 2282 -462 2292 -402
rect 2352 -462 2612 -402
rect 2672 -462 2682 -402
rect 2282 -472 2682 -462
rect 2740 -402 3140 -293
rect 2740 -462 2750 -402
rect 2810 -462 3070 -402
rect 3130 -462 3140 -402
rect 2740 -472 3140 -462
rect 3196 -402 3596 -293
rect 3196 -462 3206 -402
rect 3266 -462 3526 -402
rect 3586 -462 3596 -402
rect 3196 -472 3596 -462
rect 3652 -402 4052 -293
rect 3652 -462 3662 -402
rect 3722 -462 3982 -402
rect 4042 -462 4052 -402
rect 3652 -472 4052 -462
rect 4110 -402 4510 -293
rect 4110 -462 4120 -402
rect 4180 -462 4440 -402
rect 4500 -462 4510 -402
rect 4110 -472 4510 -462
rect 4566 -402 4966 -293
rect 4566 -462 4576 -402
rect 4636 -462 4896 -402
rect 4956 -462 4966 -402
rect 4566 -472 4966 -462
rect 5022 -402 5422 -293
rect 5022 -462 5032 -402
rect 5092 -462 5352 -402
rect 5412 -462 5422 -402
rect 5022 -472 5422 -462
rect 5480 -402 5880 -293
rect 5480 -462 5490 -402
rect 5550 -462 5810 -402
rect 5870 -462 5880 -402
rect 5480 -472 5880 -462
rect 5936 -402 6336 -293
rect 5936 -462 5946 -402
rect 6006 -462 6266 -402
rect 6326 -462 6336 -402
rect 5936 -472 6336 -462
rect 6392 -402 6792 -293
rect 6392 -462 6402 -402
rect 6462 -462 6722 -402
rect 6782 -462 6792 -402
rect 6392 -472 6792 -462
rect 6850 -402 7250 -293
rect 6850 -462 6860 -402
rect 6920 -462 7180 -402
rect 7240 -462 7250 -402
rect 6850 -472 7250 -462
rect 7306 -402 7706 -293
rect 7306 -462 7316 -402
rect 7376 -462 7636 -402
rect 7696 -462 7706 -402
rect 7306 -472 7706 -462
rect 7762 -402 8162 -293
rect 7762 -462 7772 -402
rect 7832 -462 8092 -402
rect 8152 -462 8162 -402
rect 7762 -472 8162 -462
rect 8236 -402 8636 -293
rect 8236 -462 8246 -402
rect 8306 -462 8566 -402
rect 8626 -462 8636 -402
rect 8236 -472 8636 -462
rect 8692 -402 9092 -293
rect 8692 -462 8702 -402
rect 8762 -462 9022 -402
rect 9082 -462 9092 -402
rect 8692 -472 9092 -462
rect 9150 -402 9550 -293
rect 9150 -462 9160 -402
rect 9220 -462 9480 -402
rect 9540 -462 9550 -402
rect 9150 -472 9550 -462
rect 9606 -402 10006 -293
rect 9606 -462 9616 -402
rect 9676 -462 9936 -402
rect 9996 -462 10006 -402
rect 9606 -472 10006 -462
rect 10062 -402 10462 -293
rect 10062 -462 10072 -402
rect 10132 -462 10392 -402
rect 10452 -462 10462 -402
rect 10062 -472 10462 -462
rect 10520 -402 10920 -293
rect 10520 -462 10530 -402
rect 10590 -462 10850 -402
rect 10910 -462 10920 -402
rect 10520 -472 10920 -462
rect 10976 -402 11376 -293
rect 10976 -462 10986 -402
rect 11046 -462 11306 -402
rect 11366 -462 11376 -402
rect 10976 -472 11376 -462
rect 11432 -402 11832 -293
rect 11432 -462 11442 -402
rect 11502 -462 11762 -402
rect 11822 -462 11832 -402
rect 11432 -472 11832 -462
rect 11890 -402 12290 -293
rect 11890 -462 11900 -402
rect 11960 -462 12220 -402
rect 12280 -462 12290 -402
rect 11890 -472 12290 -462
rect 12346 -402 12746 -293
rect 12346 -462 12356 -402
rect 12416 -462 12676 -402
rect 12736 -462 12746 -402
rect 12346 -472 12746 -462
rect 12802 -402 13202 -293
rect 12802 -462 12812 -402
rect 12872 -462 13132 -402
rect 13192 -462 13202 -402
rect 12802 -472 13202 -462
rect 13260 -402 13660 -293
rect 13260 -462 13270 -402
rect 13330 -462 13590 -402
rect 13650 -462 13660 -402
rect 13260 -472 13660 -462
rect 13716 -402 14116 -293
rect 13716 -462 13726 -402
rect 13786 -462 14046 -402
rect 14106 -462 14116 -402
rect 13716 -472 14116 -462
rect 14172 -402 14572 -293
rect 14172 -462 14182 -402
rect 14242 -462 14502 -402
rect 14562 -462 14572 -402
rect 14172 -472 14572 -462
rect 14630 -402 15030 -293
rect 14630 -462 14640 -402
rect 14700 -462 14960 -402
rect 15020 -462 15030 -402
rect 14630 -472 15030 -462
rect 15086 -402 15486 -293
rect 15086 -462 15096 -402
rect 15156 -462 15416 -402
rect 15476 -462 15486 -402
rect 15086 -472 15486 -462
rect 66 -544 80 -472
rect 456 -544 526 -472
rect 912 -544 983 -472
rect 1370 -544 1441 -472
rect 1826 -544 1897 -472
rect 2282 -544 2353 -472
rect 2740 -544 2811 -472
rect 3196 -544 3267 -472
rect 3652 -544 3723 -472
rect 4110 -544 4181 -472
rect 4566 -544 4637 -472
rect 5022 -544 5093 -472
rect 5480 -544 5551 -472
rect 5936 -544 6007 -472
rect 6392 -544 6463 -472
rect 6850 -544 6921 -472
rect 7306 -544 7377 -472
rect 7762 -544 7833 -472
rect 8236 -544 8307 -472
rect 8692 -544 8763 -472
rect 9150 -544 9221 -472
rect 9606 -544 9677 -472
rect 10062 -544 10133 -472
rect 10520 -544 10591 -472
rect 10976 -544 11047 -472
rect 11432 -544 11503 -472
rect 11890 -544 11961 -472
rect 12346 -544 12417 -472
rect 12802 -544 12873 -472
rect 13260 -544 13331 -472
rect 13716 -544 13787 -472
rect 14172 -544 14243 -472
rect 14630 -544 14701 -472
rect 66 -554 400 -544
rect 0 -614 10 -554
rect 70 -614 330 -554
rect 390 -614 400 -554
rect 0 -904 14 -614
rect 66 -904 400 -614
rect 0 -964 10 -904
rect 70 -964 330 -904
rect 390 -964 400 -904
rect 0 -1046 14 -964
rect 66 -974 400 -964
rect 456 -554 856 -544
rect 456 -614 466 -554
rect 526 -614 786 -554
rect 846 -614 856 -554
rect 456 -724 856 -614
rect 912 -554 1312 -544
rect 912 -614 922 -554
rect 982 -614 1242 -554
rect 1302 -614 1312 -554
rect 912 -724 1312 -614
rect 1370 -554 1770 -544
rect 1370 -614 1380 -554
rect 1440 -614 1700 -554
rect 1760 -614 1770 -554
rect 1370 -724 1770 -614
rect 1826 -554 2226 -544
rect 1826 -614 1836 -554
rect 1896 -614 2156 -554
rect 2216 -614 2226 -554
rect 1826 -724 2226 -614
rect 2282 -554 2682 -544
rect 2282 -614 2292 -554
rect 2352 -614 2612 -554
rect 2672 -614 2682 -554
rect 2282 -724 2682 -614
rect 2740 -554 3140 -544
rect 2740 -614 2750 -554
rect 2810 -614 3070 -554
rect 3130 -614 3140 -554
rect 2740 -724 3140 -614
rect 3196 -554 3596 -544
rect 3196 -614 3206 -554
rect 3266 -614 3526 -554
rect 3586 -614 3596 -554
rect 3196 -724 3596 -614
rect 3652 -554 4052 -544
rect 3652 -614 3662 -554
rect 3722 -614 3982 -554
rect 4042 -614 4052 -554
rect 3652 -724 4052 -614
rect 4110 -554 4510 -544
rect 4110 -614 4120 -554
rect 4180 -614 4440 -554
rect 4500 -614 4510 -554
rect 4110 -724 4510 -614
rect 4566 -554 4966 -544
rect 4566 -614 4576 -554
rect 4636 -614 4896 -554
rect 4956 -614 4966 -554
rect 4566 -724 4966 -614
rect 5022 -554 5422 -544
rect 5022 -614 5032 -554
rect 5092 -614 5352 -554
rect 5412 -614 5422 -554
rect 5022 -724 5422 -614
rect 5480 -554 5880 -544
rect 5480 -614 5490 -554
rect 5550 -614 5810 -554
rect 5870 -614 5880 -554
rect 5480 -724 5880 -614
rect 5936 -554 6336 -544
rect 5936 -614 5946 -554
rect 6006 -614 6266 -554
rect 6326 -614 6336 -554
rect 5936 -724 6336 -614
rect 6392 -554 6792 -544
rect 6392 -614 6402 -554
rect 6462 -614 6722 -554
rect 6782 -614 6792 -554
rect 6392 -724 6792 -614
rect 6850 -554 7250 -544
rect 6850 -614 6860 -554
rect 6920 -614 7180 -554
rect 7240 -614 7250 -554
rect 6850 -724 7250 -614
rect 7306 -554 7706 -544
rect 7306 -614 7316 -554
rect 7376 -614 7636 -554
rect 7696 -614 7706 -554
rect 7306 -724 7706 -614
rect 7762 -554 8162 -544
rect 7762 -614 7772 -554
rect 7832 -614 8092 -554
rect 8152 -614 8162 -554
rect 7762 -724 8162 -614
rect 8236 -554 8636 -544
rect 8236 -614 8246 -554
rect 8306 -614 8566 -554
rect 8626 -614 8636 -554
rect 8236 -724 8636 -614
rect 8692 -554 9092 -544
rect 8692 -614 8702 -554
rect 8762 -614 9022 -554
rect 9082 -614 9092 -554
rect 8692 -724 9092 -614
rect 9150 -554 9550 -544
rect 9150 -614 9160 -554
rect 9220 -614 9480 -554
rect 9540 -614 9550 -554
rect 9150 -724 9550 -614
rect 9606 -554 10006 -544
rect 9606 -614 9616 -554
rect 9676 -614 9936 -554
rect 9996 -614 10006 -554
rect 9606 -724 10006 -614
rect 10062 -554 10462 -544
rect 10062 -614 10072 -554
rect 10132 -614 10392 -554
rect 10452 -614 10462 -554
rect 10062 -724 10462 -614
rect 10520 -554 10920 -544
rect 10520 -614 10530 -554
rect 10590 -614 10850 -554
rect 10910 -614 10920 -554
rect 10520 -724 10920 -614
rect 10976 -554 11376 -544
rect 10976 -614 10986 -554
rect 11046 -614 11306 -554
rect 11366 -614 11376 -554
rect 10976 -724 11376 -614
rect 11432 -554 11832 -544
rect 11432 -614 11442 -554
rect 11502 -614 11762 -554
rect 11822 -614 11832 -554
rect 11432 -724 11832 -614
rect 11890 -554 12290 -544
rect 11890 -614 11900 -554
rect 11960 -614 12220 -554
rect 12280 -614 12290 -554
rect 11890 -724 12290 -614
rect 12346 -554 12746 -544
rect 12346 -614 12356 -554
rect 12416 -614 12676 -554
rect 12736 -614 12746 -554
rect 12346 -724 12746 -614
rect 12802 -554 13202 -544
rect 12802 -614 12812 -554
rect 12872 -614 13132 -554
rect 13192 -614 13202 -554
rect 12802 -724 13202 -614
rect 13260 -554 13660 -544
rect 13260 -614 13270 -554
rect 13330 -614 13590 -554
rect 13650 -614 13660 -554
rect 13260 -724 13660 -614
rect 13716 -554 14116 -544
rect 13716 -614 13726 -554
rect 13786 -614 14046 -554
rect 14106 -614 14116 -554
rect 13716 -724 14116 -614
rect 14172 -554 14572 -544
rect 14172 -614 14182 -554
rect 14242 -614 14502 -554
rect 14562 -614 14572 -554
rect 14172 -724 14572 -614
rect 14630 -554 15030 -544
rect 14630 -614 14640 -554
rect 14700 -614 14960 -554
rect 15020 -614 15030 -554
rect 14630 -724 15030 -614
rect 15086 -554 15486 -544
rect 15086 -614 15096 -554
rect 15156 -614 15416 -554
rect 15476 -614 15486 -554
rect 15086 -724 15486 -614
rect 456 -794 15486 -724
rect 456 -904 856 -794
rect 456 -964 466 -904
rect 526 -964 786 -904
rect 846 -964 856 -904
rect 456 -974 856 -964
rect 912 -904 1312 -794
rect 912 -964 922 -904
rect 982 -964 1242 -904
rect 1302 -964 1312 -904
rect 912 -974 1312 -964
rect 1370 -904 1770 -794
rect 1370 -964 1380 -904
rect 1440 -964 1700 -904
rect 1760 -964 1770 -904
rect 1370 -974 1770 -964
rect 1826 -904 2226 -794
rect 1826 -964 1836 -904
rect 1896 -964 2156 -904
rect 2216 -964 2226 -904
rect 1826 -974 2226 -964
rect 2282 -904 2682 -794
rect 2282 -964 2292 -904
rect 2352 -964 2612 -904
rect 2672 -964 2682 -904
rect 2282 -974 2682 -964
rect 2740 -904 3140 -794
rect 2740 -964 2750 -904
rect 2810 -964 3070 -904
rect 3130 -964 3140 -904
rect 2740 -974 3140 -964
rect 3196 -904 3596 -794
rect 3196 -964 3206 -904
rect 3266 -964 3526 -904
rect 3586 -964 3596 -904
rect 3196 -974 3596 -964
rect 3652 -904 4052 -794
rect 3652 -964 3662 -904
rect 3722 -964 3982 -904
rect 4042 -964 4052 -904
rect 3652 -974 4052 -964
rect 4110 -904 4510 -794
rect 4110 -964 4120 -904
rect 4180 -964 4440 -904
rect 4500 -964 4510 -904
rect 4110 -974 4510 -964
rect 4566 -904 4966 -794
rect 4566 -964 4576 -904
rect 4636 -964 4896 -904
rect 4956 -964 4966 -904
rect 4566 -974 4966 -964
rect 5022 -904 5422 -794
rect 5022 -964 5032 -904
rect 5092 -964 5352 -904
rect 5412 -964 5422 -904
rect 5022 -974 5422 -964
rect 5480 -904 5880 -794
rect 5480 -964 5490 -904
rect 5550 -964 5810 -904
rect 5870 -964 5880 -904
rect 5480 -974 5880 -964
rect 5936 -904 6336 -794
rect 5936 -964 5946 -904
rect 6006 -964 6266 -904
rect 6326 -964 6336 -904
rect 5936 -974 6336 -964
rect 6392 -904 6792 -794
rect 6392 -964 6402 -904
rect 6462 -964 6722 -904
rect 6782 -964 6792 -904
rect 6392 -974 6792 -964
rect 6850 -904 7250 -794
rect 6850 -964 6860 -904
rect 6920 -964 7180 -904
rect 7240 -964 7250 -904
rect 6850 -974 7250 -964
rect 7306 -904 7706 -794
rect 7306 -964 7316 -904
rect 7376 -964 7636 -904
rect 7696 -964 7706 -904
rect 7306 -974 7706 -964
rect 7762 -904 8162 -794
rect 7762 -964 7772 -904
rect 7832 -964 8092 -904
rect 8152 -964 8162 -904
rect 7762 -974 8162 -964
rect 8236 -904 8636 -794
rect 8236 -964 8246 -904
rect 8306 -964 8566 -904
rect 8626 -964 8636 -904
rect 8236 -974 8636 -964
rect 8692 -904 9092 -794
rect 8692 -964 8702 -904
rect 8762 -964 9022 -904
rect 9082 -964 9092 -904
rect 8692 -974 9092 -964
rect 9150 -904 9550 -794
rect 9150 -964 9160 -904
rect 9220 -964 9480 -904
rect 9540 -964 9550 -904
rect 9150 -974 9550 -964
rect 9606 -904 10006 -794
rect 9606 -964 9616 -904
rect 9676 -964 9936 -904
rect 9996 -964 10006 -904
rect 9606 -974 10006 -964
rect 10062 -904 10462 -794
rect 10062 -964 10072 -904
rect 10132 -964 10392 -904
rect 10452 -964 10462 -904
rect 10062 -974 10462 -964
rect 10520 -904 10920 -794
rect 10520 -964 10530 -904
rect 10590 -964 10850 -904
rect 10910 -964 10920 -904
rect 10520 -974 10920 -964
rect 10976 -904 11376 -794
rect 10976 -964 10986 -904
rect 11046 -964 11306 -904
rect 11366 -964 11376 -904
rect 10976 -974 11376 -964
rect 11432 -904 11832 -794
rect 11432 -964 11442 -904
rect 11502 -964 11762 -904
rect 11822 -964 11832 -904
rect 11432 -974 11832 -964
rect 11890 -904 12290 -794
rect 11890 -964 11900 -904
rect 11960 -964 12220 -904
rect 12280 -964 12290 -904
rect 11890 -974 12290 -964
rect 12346 -904 12746 -794
rect 12346 -964 12356 -904
rect 12416 -964 12676 -904
rect 12736 -964 12746 -904
rect 12346 -974 12746 -964
rect 12802 -904 13202 -794
rect 12802 -964 12812 -904
rect 12872 -964 13132 -904
rect 13192 -964 13202 -904
rect 12802 -974 13202 -964
rect 13260 -904 13660 -794
rect 13260 -964 13270 -904
rect 13330 -964 13590 -904
rect 13650 -964 13660 -904
rect 13260 -974 13660 -964
rect 13716 -904 14116 -794
rect 13716 -964 13726 -904
rect 13786 -964 14046 -904
rect 14106 -964 14116 -904
rect 13716 -974 14116 -964
rect 14172 -904 14572 -794
rect 14172 -964 14182 -904
rect 14242 -964 14502 -904
rect 14562 -964 14572 -904
rect 14172 -974 14572 -964
rect 14630 -904 15030 -794
rect 14630 -964 14640 -904
rect 14700 -964 14960 -904
rect 15020 -964 15030 -904
rect 14630 -974 15030 -964
rect 15086 -904 15486 -794
rect 15086 -964 15096 -904
rect 15156 -964 15416 -904
rect 15476 -964 15486 -904
rect 15086 -974 15486 -964
rect 66 -1036 80 -974
rect 456 -1036 527 -974
rect 912 -1036 983 -974
rect 1370 -1036 1441 -974
rect 1826 -1036 1897 -974
rect 2282 -1036 2353 -974
rect 2740 -1036 2810 -974
rect 3196 -1036 3266 -974
rect 3652 -1036 3722 -974
rect 4110 -1036 4180 -974
rect 4566 -1036 4636 -974
rect 5022 -1036 5092 -974
rect 5480 -1036 5550 -974
rect 5936 -1036 6006 -974
rect 6392 -1036 6462 -974
rect 6850 -1036 6920 -974
rect 7306 -1036 7376 -974
rect 7762 -1036 7832 -974
rect 8236 -1036 8306 -974
rect 8692 -1036 8762 -974
rect 9150 -1036 9220 -974
rect 9606 -1036 9676 -974
rect 10062 -1036 10132 -974
rect 10520 -1036 10590 -974
rect 10976 -1036 11046 -974
rect 11432 -1036 11502 -974
rect 11890 -1036 11960 -974
rect 12346 -1036 12416 -974
rect 12802 -1036 12872 -974
rect 13260 -1036 13330 -974
rect 13716 -1036 13786 -974
rect 14172 -1036 14242 -974
rect 14630 -1036 14700 -974
rect 66 -1046 400 -1036
rect 0 -1106 10 -1046
rect 70 -1106 330 -1046
rect 390 -1106 400 -1046
rect 0 -1396 14 -1106
rect 66 -1396 400 -1106
rect 0 -1456 10 -1396
rect 70 -1456 330 -1396
rect 390 -1456 400 -1396
rect 0 -1562 14 -1456
rect 66 -1466 400 -1456
rect 456 -1046 856 -1036
rect 456 -1106 466 -1046
rect 526 -1106 786 -1046
rect 846 -1106 856 -1046
rect 456 -1216 856 -1106
rect 912 -1046 1312 -1036
rect 912 -1106 922 -1046
rect 982 -1106 1242 -1046
rect 1302 -1106 1312 -1046
rect 912 -1216 1312 -1106
rect 1370 -1046 1770 -1036
rect 1370 -1106 1380 -1046
rect 1440 -1106 1700 -1046
rect 1760 -1106 1770 -1046
rect 1370 -1216 1770 -1106
rect 1826 -1046 2226 -1036
rect 1826 -1106 1836 -1046
rect 1896 -1106 2156 -1046
rect 2216 -1106 2226 -1046
rect 1826 -1216 2226 -1106
rect 2282 -1046 2682 -1036
rect 2282 -1106 2292 -1046
rect 2352 -1106 2612 -1046
rect 2672 -1106 2682 -1046
rect 2282 -1216 2682 -1106
rect 2740 -1046 3140 -1036
rect 2740 -1106 2750 -1046
rect 2810 -1106 3070 -1046
rect 3130 -1106 3140 -1046
rect 2740 -1216 3140 -1106
rect 3196 -1046 3596 -1036
rect 3196 -1106 3206 -1046
rect 3266 -1106 3526 -1046
rect 3586 -1106 3596 -1046
rect 3196 -1216 3596 -1106
rect 3652 -1046 4052 -1036
rect 3652 -1106 3662 -1046
rect 3722 -1106 3982 -1046
rect 4042 -1106 4052 -1046
rect 3652 -1216 4052 -1106
rect 4110 -1046 4510 -1036
rect 4110 -1106 4120 -1046
rect 4180 -1106 4440 -1046
rect 4500 -1106 4510 -1046
rect 4110 -1216 4510 -1106
rect 4566 -1046 4966 -1036
rect 4566 -1106 4576 -1046
rect 4636 -1106 4896 -1046
rect 4956 -1106 4966 -1046
rect 4566 -1216 4966 -1106
rect 5022 -1046 5422 -1036
rect 5022 -1106 5032 -1046
rect 5092 -1106 5352 -1046
rect 5412 -1106 5422 -1046
rect 5022 -1216 5422 -1106
rect 5480 -1046 5880 -1036
rect 5480 -1106 5490 -1046
rect 5550 -1106 5810 -1046
rect 5870 -1106 5880 -1046
rect 5480 -1216 5880 -1106
rect 5936 -1046 6336 -1036
rect 5936 -1106 5946 -1046
rect 6006 -1106 6266 -1046
rect 6326 -1106 6336 -1046
rect 5936 -1216 6336 -1106
rect 6392 -1046 6792 -1036
rect 6392 -1106 6402 -1046
rect 6462 -1106 6722 -1046
rect 6782 -1106 6792 -1046
rect 6392 -1216 6792 -1106
rect 6850 -1046 7250 -1036
rect 6850 -1106 6860 -1046
rect 6920 -1106 7180 -1046
rect 7240 -1106 7250 -1046
rect 6850 -1216 7250 -1106
rect 7306 -1046 7706 -1036
rect 7306 -1106 7316 -1046
rect 7376 -1106 7636 -1046
rect 7696 -1106 7706 -1046
rect 7306 -1216 7706 -1106
rect 7762 -1046 8162 -1036
rect 7762 -1106 7772 -1046
rect 7832 -1106 8092 -1046
rect 8152 -1106 8162 -1046
rect 7762 -1216 8162 -1106
rect 8236 -1046 8636 -1036
rect 8236 -1106 8246 -1046
rect 8306 -1106 8566 -1046
rect 8626 -1106 8636 -1046
rect 8236 -1216 8636 -1106
rect 8692 -1046 9092 -1036
rect 8692 -1106 8702 -1046
rect 8762 -1106 9022 -1046
rect 9082 -1106 9092 -1046
rect 8692 -1216 9092 -1106
rect 9150 -1046 9550 -1036
rect 9150 -1106 9160 -1046
rect 9220 -1106 9480 -1046
rect 9540 -1106 9550 -1046
rect 9150 -1216 9550 -1106
rect 9606 -1046 10006 -1036
rect 9606 -1106 9616 -1046
rect 9676 -1106 9936 -1046
rect 9996 -1106 10006 -1046
rect 9606 -1216 10006 -1106
rect 10062 -1046 10462 -1036
rect 10062 -1106 10072 -1046
rect 10132 -1106 10392 -1046
rect 10452 -1106 10462 -1046
rect 10062 -1216 10462 -1106
rect 10520 -1046 10920 -1036
rect 10520 -1106 10530 -1046
rect 10590 -1106 10850 -1046
rect 10910 -1106 10920 -1046
rect 10520 -1216 10920 -1106
rect 10976 -1046 11376 -1036
rect 10976 -1106 10986 -1046
rect 11046 -1106 11306 -1046
rect 11366 -1106 11376 -1046
rect 10976 -1216 11376 -1106
rect 11432 -1046 11832 -1036
rect 11432 -1106 11442 -1046
rect 11502 -1106 11762 -1046
rect 11822 -1106 11832 -1046
rect 11432 -1216 11832 -1106
rect 11890 -1046 12290 -1036
rect 11890 -1106 11900 -1046
rect 11960 -1106 12220 -1046
rect 12280 -1106 12290 -1046
rect 11890 -1216 12290 -1106
rect 12346 -1046 12746 -1036
rect 12346 -1106 12356 -1046
rect 12416 -1106 12676 -1046
rect 12736 -1106 12746 -1046
rect 12346 -1216 12746 -1106
rect 12802 -1046 13202 -1036
rect 12802 -1106 12812 -1046
rect 12872 -1106 13132 -1046
rect 13192 -1106 13202 -1046
rect 12802 -1216 13202 -1106
rect 13260 -1046 13660 -1036
rect 13260 -1106 13270 -1046
rect 13330 -1106 13590 -1046
rect 13650 -1106 13660 -1046
rect 13260 -1216 13660 -1106
rect 13716 -1046 14116 -1036
rect 13716 -1106 13726 -1046
rect 13786 -1106 14046 -1046
rect 14106 -1106 14116 -1046
rect 13716 -1216 14116 -1106
rect 14172 -1046 14572 -1036
rect 14172 -1106 14182 -1046
rect 14242 -1106 14502 -1046
rect 14562 -1106 14572 -1046
rect 14172 -1216 14572 -1106
rect 14630 -1046 15030 -1036
rect 14630 -1106 14640 -1046
rect 14700 -1106 14960 -1046
rect 15020 -1106 15030 -1046
rect 14630 -1216 15030 -1106
rect 15086 -1046 15486 -1036
rect 15086 -1106 15096 -1046
rect 15156 -1106 15416 -1046
rect 15476 -1106 15486 -1046
rect 15086 -1216 15486 -1106
rect 456 -1286 15486 -1216
rect 456 -1396 856 -1286
rect 456 -1456 466 -1396
rect 526 -1456 786 -1396
rect 846 -1456 856 -1396
rect 456 -1466 856 -1456
rect 912 -1396 1312 -1286
rect 912 -1456 922 -1396
rect 982 -1456 1242 -1396
rect 1302 -1456 1312 -1396
rect 912 -1466 1312 -1456
rect 1370 -1396 1770 -1286
rect 1370 -1456 1380 -1396
rect 1440 -1456 1700 -1396
rect 1760 -1456 1770 -1396
rect 1370 -1466 1770 -1456
rect 1826 -1396 2226 -1286
rect 1826 -1456 1836 -1396
rect 1896 -1456 2156 -1396
rect 2216 -1456 2226 -1396
rect 1826 -1466 2226 -1456
rect 2282 -1396 2682 -1286
rect 2282 -1456 2292 -1396
rect 2352 -1456 2612 -1396
rect 2672 -1456 2682 -1396
rect 2282 -1466 2682 -1456
rect 2740 -1396 3140 -1286
rect 2740 -1456 2750 -1396
rect 2810 -1456 3070 -1396
rect 3130 -1456 3140 -1396
rect 2740 -1466 3140 -1456
rect 3196 -1396 3596 -1286
rect 3196 -1456 3206 -1396
rect 3266 -1456 3526 -1396
rect 3586 -1456 3596 -1396
rect 3196 -1466 3596 -1456
rect 3652 -1396 4052 -1286
rect 3652 -1456 3662 -1396
rect 3722 -1456 3982 -1396
rect 4042 -1456 4052 -1396
rect 3652 -1466 4052 -1456
rect 4110 -1396 4510 -1286
rect 4110 -1456 4120 -1396
rect 4180 -1456 4440 -1396
rect 4500 -1456 4510 -1396
rect 4110 -1466 4510 -1456
rect 4566 -1396 4966 -1286
rect 4566 -1456 4576 -1396
rect 4636 -1456 4896 -1396
rect 4956 -1456 4966 -1396
rect 4566 -1466 4966 -1456
rect 5022 -1396 5422 -1286
rect 5022 -1456 5032 -1396
rect 5092 -1456 5352 -1396
rect 5412 -1456 5422 -1396
rect 5022 -1466 5422 -1456
rect 5480 -1396 5880 -1286
rect 5480 -1456 5490 -1396
rect 5550 -1456 5810 -1396
rect 5870 -1456 5880 -1396
rect 5480 -1466 5880 -1456
rect 5936 -1396 6336 -1286
rect 5936 -1456 5946 -1396
rect 6006 -1456 6266 -1396
rect 6326 -1456 6336 -1396
rect 5936 -1466 6336 -1456
rect 6392 -1396 6792 -1286
rect 6392 -1456 6402 -1396
rect 6462 -1456 6722 -1396
rect 6782 -1456 6792 -1396
rect 6392 -1466 6792 -1456
rect 6850 -1396 7250 -1286
rect 6850 -1456 6860 -1396
rect 6920 -1456 7180 -1396
rect 7240 -1456 7250 -1396
rect 6850 -1466 7250 -1456
rect 7306 -1396 7706 -1286
rect 7306 -1456 7316 -1396
rect 7376 -1456 7636 -1396
rect 7696 -1456 7706 -1396
rect 7306 -1466 7706 -1456
rect 7762 -1396 8162 -1286
rect 7762 -1456 7772 -1396
rect 7832 -1456 8092 -1396
rect 8152 -1456 8162 -1396
rect 7762 -1466 8162 -1456
rect 8236 -1396 8636 -1286
rect 8236 -1456 8246 -1396
rect 8306 -1456 8566 -1396
rect 8626 -1456 8636 -1396
rect 8236 -1466 8636 -1456
rect 8692 -1396 9092 -1286
rect 8692 -1456 8702 -1396
rect 8762 -1456 9022 -1396
rect 9082 -1456 9092 -1396
rect 8692 -1466 9092 -1456
rect 9150 -1396 9550 -1286
rect 9150 -1456 9160 -1396
rect 9220 -1456 9480 -1396
rect 9540 -1456 9550 -1396
rect 9150 -1466 9550 -1456
rect 9606 -1396 10006 -1286
rect 9606 -1456 9616 -1396
rect 9676 -1456 9936 -1396
rect 9996 -1456 10006 -1396
rect 9606 -1466 10006 -1456
rect 10062 -1396 10462 -1286
rect 10062 -1456 10072 -1396
rect 10132 -1456 10392 -1396
rect 10452 -1456 10462 -1396
rect 10062 -1466 10462 -1456
rect 10520 -1396 10920 -1286
rect 10520 -1456 10530 -1396
rect 10590 -1456 10850 -1396
rect 10910 -1456 10920 -1396
rect 10520 -1466 10920 -1456
rect 10976 -1396 11376 -1286
rect 10976 -1456 10986 -1396
rect 11046 -1456 11306 -1396
rect 11366 -1456 11376 -1396
rect 10976 -1466 11376 -1456
rect 11432 -1396 11832 -1286
rect 11432 -1456 11442 -1396
rect 11502 -1456 11762 -1396
rect 11822 -1456 11832 -1396
rect 11432 -1466 11832 -1456
rect 11890 -1396 12290 -1286
rect 11890 -1456 11900 -1396
rect 11960 -1456 12220 -1396
rect 12280 -1456 12290 -1396
rect 11890 -1466 12290 -1456
rect 12346 -1396 12746 -1286
rect 12346 -1456 12356 -1396
rect 12416 -1456 12676 -1396
rect 12736 -1456 12746 -1396
rect 12346 -1466 12746 -1456
rect 12802 -1396 13202 -1286
rect 12802 -1456 12812 -1396
rect 12872 -1456 13132 -1396
rect 13192 -1456 13202 -1396
rect 12802 -1466 13202 -1456
rect 13260 -1396 13660 -1286
rect 13260 -1456 13270 -1396
rect 13330 -1456 13590 -1396
rect 13650 -1456 13660 -1396
rect 13260 -1466 13660 -1456
rect 13716 -1396 14116 -1286
rect 13716 -1456 13726 -1396
rect 13786 -1456 14046 -1396
rect 14106 -1456 14116 -1396
rect 13716 -1466 14116 -1456
rect 14172 -1396 14572 -1286
rect 14172 -1456 14182 -1396
rect 14242 -1456 14502 -1396
rect 14562 -1456 14572 -1396
rect 14172 -1466 14572 -1456
rect 14630 -1396 15030 -1286
rect 14630 -1456 14640 -1396
rect 14700 -1456 14960 -1396
rect 15020 -1456 15030 -1396
rect 14630 -1466 15030 -1456
rect 15086 -1396 15486 -1286
rect 15086 -1456 15096 -1396
rect 15156 -1456 15416 -1396
rect 15476 -1456 15486 -1396
rect 15086 -1466 15486 -1456
rect 66 -1552 80 -1466
rect 456 -1552 526 -1466
rect 912 -1552 982 -1466
rect 1370 -1552 1440 -1466
rect 1826 -1552 1896 -1466
rect 2282 -1552 2352 -1466
rect 2740 -1552 2810 -1466
rect 3196 -1552 3266 -1466
rect 3652 -1552 3722 -1466
rect 4110 -1552 4180 -1466
rect 4566 -1552 4636 -1466
rect 5022 -1552 5092 -1466
rect 5480 -1552 5550 -1466
rect 5936 -1552 6006 -1466
rect 6392 -1552 6462 -1466
rect 6850 -1552 6920 -1466
rect 7306 -1552 7376 -1466
rect 7762 -1552 7832 -1466
rect 8236 -1552 8306 -1466
rect 8692 -1552 8762 -1466
rect 9150 -1552 9220 -1466
rect 9606 -1552 9676 -1466
rect 10062 -1552 10132 -1466
rect 10520 -1552 10590 -1466
rect 10976 -1552 11046 -1466
rect 11432 -1552 11502 -1466
rect 11890 -1552 11960 -1466
rect 12346 -1552 12416 -1466
rect 12802 -1552 12872 -1466
rect 13260 -1552 13330 -1466
rect 13716 -1552 13786 -1466
rect 14172 -1552 14242 -1466
rect 14630 -1552 14700 -1466
rect 66 -1562 400 -1552
rect 0 -1622 10 -1562
rect 70 -1622 330 -1562
rect 390 -1622 400 -1562
rect 0 -1912 14 -1622
rect 66 -1912 400 -1622
rect 0 -1972 10 -1912
rect 70 -1972 330 -1912
rect 390 -1972 400 -1912
rect 0 -2064 14 -1972
rect 66 -1982 400 -1972
rect 456 -1562 856 -1552
rect 456 -1622 466 -1562
rect 526 -1622 786 -1562
rect 846 -1622 856 -1562
rect 456 -1732 856 -1622
rect 912 -1562 1312 -1552
rect 912 -1622 922 -1562
rect 982 -1622 1242 -1562
rect 1302 -1622 1312 -1562
rect 912 -1732 1312 -1622
rect 1370 -1562 1770 -1552
rect 1370 -1622 1380 -1562
rect 1440 -1622 1700 -1562
rect 1760 -1622 1770 -1562
rect 1370 -1732 1770 -1622
rect 1826 -1562 2226 -1552
rect 1826 -1622 1836 -1562
rect 1896 -1622 2156 -1562
rect 2216 -1622 2226 -1562
rect 1826 -1732 2226 -1622
rect 2282 -1562 2682 -1552
rect 2282 -1622 2292 -1562
rect 2352 -1622 2612 -1562
rect 2672 -1622 2682 -1562
rect 2282 -1732 2682 -1622
rect 2740 -1562 3140 -1552
rect 2740 -1622 2750 -1562
rect 2810 -1622 3070 -1562
rect 3130 -1622 3140 -1562
rect 2740 -1732 3140 -1622
rect 3196 -1562 3596 -1552
rect 3196 -1622 3206 -1562
rect 3266 -1622 3526 -1562
rect 3586 -1622 3596 -1562
rect 3196 -1732 3596 -1622
rect 3652 -1562 4052 -1552
rect 3652 -1622 3662 -1562
rect 3722 -1622 3982 -1562
rect 4042 -1622 4052 -1562
rect 3652 -1732 4052 -1622
rect 4110 -1562 4510 -1552
rect 4110 -1622 4120 -1562
rect 4180 -1622 4440 -1562
rect 4500 -1622 4510 -1562
rect 4110 -1732 4510 -1622
rect 4566 -1562 4966 -1552
rect 4566 -1622 4576 -1562
rect 4636 -1622 4896 -1562
rect 4956 -1622 4966 -1562
rect 4566 -1732 4966 -1622
rect 5022 -1562 5422 -1552
rect 5022 -1622 5032 -1562
rect 5092 -1622 5352 -1562
rect 5412 -1622 5422 -1562
rect 5022 -1732 5422 -1622
rect 5480 -1562 5880 -1552
rect 5480 -1622 5490 -1562
rect 5550 -1622 5810 -1562
rect 5870 -1622 5880 -1562
rect 5480 -1732 5880 -1622
rect 5936 -1562 6336 -1552
rect 5936 -1622 5946 -1562
rect 6006 -1622 6266 -1562
rect 6326 -1622 6336 -1562
rect 5936 -1732 6336 -1622
rect 6392 -1562 6792 -1552
rect 6392 -1622 6402 -1562
rect 6462 -1622 6722 -1562
rect 6782 -1622 6792 -1562
rect 6392 -1732 6792 -1622
rect 6850 -1562 7250 -1552
rect 6850 -1622 6860 -1562
rect 6920 -1622 7180 -1562
rect 7240 -1622 7250 -1562
rect 6850 -1732 7250 -1622
rect 7306 -1562 7706 -1552
rect 7306 -1622 7316 -1562
rect 7376 -1622 7636 -1562
rect 7696 -1622 7706 -1562
rect 7306 -1732 7706 -1622
rect 7762 -1562 8162 -1552
rect 7762 -1622 7772 -1562
rect 7832 -1622 8092 -1562
rect 8152 -1622 8162 -1562
rect 7762 -1732 8162 -1622
rect 8236 -1562 8636 -1552
rect 8236 -1622 8246 -1562
rect 8306 -1622 8566 -1562
rect 8626 -1622 8636 -1562
rect 8236 -1732 8636 -1622
rect 8692 -1562 9092 -1552
rect 8692 -1622 8702 -1562
rect 8762 -1622 9022 -1562
rect 9082 -1622 9092 -1562
rect 8692 -1732 9092 -1622
rect 9150 -1562 9550 -1552
rect 9150 -1622 9160 -1562
rect 9220 -1622 9480 -1562
rect 9540 -1622 9550 -1562
rect 9150 -1732 9550 -1622
rect 9606 -1562 10006 -1552
rect 9606 -1622 9616 -1562
rect 9676 -1622 9936 -1562
rect 9996 -1622 10006 -1562
rect 9606 -1732 10006 -1622
rect 10062 -1562 10462 -1552
rect 10062 -1622 10072 -1562
rect 10132 -1622 10392 -1562
rect 10452 -1622 10462 -1562
rect 10062 -1732 10462 -1622
rect 10520 -1562 10920 -1552
rect 10520 -1622 10530 -1562
rect 10590 -1622 10850 -1562
rect 10910 -1622 10920 -1562
rect 10520 -1732 10920 -1622
rect 10976 -1562 11376 -1552
rect 10976 -1622 10986 -1562
rect 11046 -1622 11306 -1562
rect 11366 -1622 11376 -1562
rect 10976 -1732 11376 -1622
rect 11432 -1562 11832 -1552
rect 11432 -1622 11442 -1562
rect 11502 -1622 11762 -1562
rect 11822 -1622 11832 -1562
rect 11432 -1732 11832 -1622
rect 11890 -1562 12290 -1552
rect 11890 -1622 11900 -1562
rect 11960 -1622 12220 -1562
rect 12280 -1622 12290 -1562
rect 11890 -1732 12290 -1622
rect 12346 -1562 12746 -1552
rect 12346 -1622 12356 -1562
rect 12416 -1622 12676 -1562
rect 12736 -1622 12746 -1562
rect 12346 -1732 12746 -1622
rect 12802 -1562 13202 -1552
rect 12802 -1622 12812 -1562
rect 12872 -1622 13132 -1562
rect 13192 -1622 13202 -1562
rect 12802 -1732 13202 -1622
rect 13260 -1562 13660 -1552
rect 13260 -1622 13270 -1562
rect 13330 -1622 13590 -1562
rect 13650 -1622 13660 -1562
rect 13260 -1732 13660 -1622
rect 13716 -1562 14116 -1552
rect 13716 -1622 13726 -1562
rect 13786 -1622 14046 -1562
rect 14106 -1622 14116 -1562
rect 13716 -1732 14116 -1622
rect 14172 -1562 14572 -1552
rect 14172 -1622 14182 -1562
rect 14242 -1622 14502 -1562
rect 14562 -1622 14572 -1562
rect 14172 -1732 14572 -1622
rect 14630 -1562 15030 -1552
rect 14630 -1622 14640 -1562
rect 14700 -1622 14960 -1562
rect 15020 -1622 15030 -1562
rect 14630 -1732 15030 -1622
rect 15086 -1562 15486 -1552
rect 15086 -1622 15096 -1562
rect 15156 -1622 15416 -1562
rect 15476 -1622 15486 -1562
rect 15086 -1732 15486 -1622
rect 456 -1802 15486 -1732
rect 456 -1912 856 -1802
rect 456 -1972 466 -1912
rect 526 -1972 786 -1912
rect 846 -1972 856 -1912
rect 456 -1982 856 -1972
rect 912 -1912 1312 -1802
rect 912 -1972 922 -1912
rect 982 -1972 1242 -1912
rect 1302 -1972 1312 -1912
rect 912 -1982 1312 -1972
rect 1370 -1912 1770 -1802
rect 1370 -1972 1380 -1912
rect 1440 -1972 1700 -1912
rect 1760 -1972 1770 -1912
rect 1370 -1982 1770 -1972
rect 1826 -1912 2226 -1802
rect 1826 -1972 1836 -1912
rect 1896 -1972 2156 -1912
rect 2216 -1972 2226 -1912
rect 1826 -1982 2226 -1972
rect 2282 -1912 2682 -1802
rect 2282 -1972 2292 -1912
rect 2352 -1972 2612 -1912
rect 2672 -1972 2682 -1912
rect 2282 -1982 2682 -1972
rect 2740 -1912 3140 -1802
rect 2740 -1972 2750 -1912
rect 2810 -1972 3070 -1912
rect 3130 -1972 3140 -1912
rect 2740 -1982 3140 -1972
rect 3196 -1912 3596 -1802
rect 3196 -1972 3206 -1912
rect 3266 -1972 3526 -1912
rect 3586 -1972 3596 -1912
rect 3196 -1982 3596 -1972
rect 3652 -1912 4052 -1802
rect 3652 -1972 3662 -1912
rect 3722 -1972 3982 -1912
rect 4042 -1972 4052 -1912
rect 3652 -1982 4052 -1972
rect 4110 -1912 4510 -1802
rect 4110 -1972 4120 -1912
rect 4180 -1972 4440 -1912
rect 4500 -1972 4510 -1912
rect 4110 -1982 4510 -1972
rect 4566 -1912 4966 -1802
rect 4566 -1972 4576 -1912
rect 4636 -1972 4896 -1912
rect 4956 -1972 4966 -1912
rect 4566 -1982 4966 -1972
rect 5022 -1912 5422 -1802
rect 5022 -1972 5032 -1912
rect 5092 -1972 5352 -1912
rect 5412 -1972 5422 -1912
rect 5022 -1982 5422 -1972
rect 5480 -1912 5880 -1802
rect 5480 -1972 5490 -1912
rect 5550 -1972 5810 -1912
rect 5870 -1972 5880 -1912
rect 5480 -1982 5880 -1972
rect 5936 -1912 6336 -1802
rect 5936 -1972 5946 -1912
rect 6006 -1972 6266 -1912
rect 6326 -1972 6336 -1912
rect 5936 -1982 6336 -1972
rect 6392 -1912 6792 -1802
rect 6392 -1972 6402 -1912
rect 6462 -1972 6722 -1912
rect 6782 -1972 6792 -1912
rect 6392 -1982 6792 -1972
rect 6850 -1912 7250 -1802
rect 6850 -1972 6860 -1912
rect 6920 -1972 7180 -1912
rect 7240 -1972 7250 -1912
rect 6850 -1982 7250 -1972
rect 7306 -1912 7706 -1802
rect 7306 -1972 7316 -1912
rect 7376 -1972 7636 -1912
rect 7696 -1972 7706 -1912
rect 7306 -1982 7706 -1972
rect 7762 -1912 8162 -1802
rect 7762 -1972 7772 -1912
rect 7832 -1972 8092 -1912
rect 8152 -1972 8162 -1912
rect 7762 -1982 8162 -1972
rect 8236 -1912 8636 -1802
rect 8236 -1972 8246 -1912
rect 8306 -1972 8566 -1912
rect 8626 -1972 8636 -1912
rect 8236 -1982 8636 -1972
rect 8692 -1912 9092 -1802
rect 8692 -1972 8702 -1912
rect 8762 -1972 9022 -1912
rect 9082 -1972 9092 -1912
rect 8692 -1982 9092 -1972
rect 9150 -1912 9550 -1802
rect 9150 -1972 9160 -1912
rect 9220 -1972 9480 -1912
rect 9540 -1972 9550 -1912
rect 9150 -1982 9550 -1972
rect 9606 -1912 10006 -1802
rect 9606 -1972 9616 -1912
rect 9676 -1972 9936 -1912
rect 9996 -1972 10006 -1912
rect 9606 -1982 10006 -1972
rect 10062 -1912 10462 -1802
rect 10062 -1972 10072 -1912
rect 10132 -1972 10392 -1912
rect 10452 -1972 10462 -1912
rect 10062 -1982 10462 -1972
rect 10520 -1912 10920 -1802
rect 10520 -1972 10530 -1912
rect 10590 -1972 10850 -1912
rect 10910 -1972 10920 -1912
rect 10520 -1982 10920 -1972
rect 10976 -1912 11376 -1802
rect 10976 -1972 10986 -1912
rect 11046 -1972 11306 -1912
rect 11366 -1972 11376 -1912
rect 10976 -1982 11376 -1972
rect 11432 -1912 11832 -1802
rect 11432 -1972 11442 -1912
rect 11502 -1972 11762 -1912
rect 11822 -1972 11832 -1912
rect 11432 -1982 11832 -1972
rect 11890 -1912 12290 -1802
rect 11890 -1972 11900 -1912
rect 11960 -1972 12220 -1912
rect 12280 -1972 12290 -1912
rect 11890 -1982 12290 -1972
rect 12346 -1912 12746 -1802
rect 12346 -1972 12356 -1912
rect 12416 -1972 12676 -1912
rect 12736 -1972 12746 -1912
rect 12346 -1982 12746 -1972
rect 12802 -1912 13202 -1802
rect 12802 -1972 12812 -1912
rect 12872 -1972 13132 -1912
rect 13192 -1972 13202 -1912
rect 12802 -1982 13202 -1972
rect 13260 -1912 13660 -1802
rect 13260 -1972 13270 -1912
rect 13330 -1972 13590 -1912
rect 13650 -1972 13660 -1912
rect 13260 -1982 13660 -1972
rect 13716 -1912 14116 -1802
rect 13716 -1972 13726 -1912
rect 13786 -1972 14046 -1912
rect 14106 -1972 14116 -1912
rect 13716 -1982 14116 -1972
rect 14172 -1912 14572 -1802
rect 14172 -1972 14182 -1912
rect 14242 -1972 14502 -1912
rect 14562 -1972 14572 -1912
rect 14172 -1982 14572 -1972
rect 14630 -1912 15030 -1802
rect 14630 -1972 14640 -1912
rect 14700 -1972 14960 -1912
rect 15020 -1972 15030 -1912
rect 14630 -1982 15030 -1972
rect 15086 -1912 15486 -1802
rect 15086 -1972 15096 -1912
rect 15156 -1972 15416 -1912
rect 15476 -1972 15486 -1912
rect 15086 -1982 15486 -1972
rect 66 -2054 80 -1982
rect 456 -2054 526 -1982
rect 912 -2054 983 -1982
rect 1370 -2054 1441 -1982
rect 1826 -2054 1897 -1982
rect 2282 -2054 2353 -1982
rect 2740 -2054 2811 -1982
rect 3196 -2054 3267 -1982
rect 3652 -2054 3723 -1982
rect 4110 -2054 4181 -1982
rect 4566 -2054 4637 -1982
rect 5022 -2054 5093 -1982
rect 5480 -2054 5551 -1982
rect 5936 -2054 6007 -1982
rect 6392 -2054 6463 -1982
rect 6850 -2054 6921 -1982
rect 7306 -2054 7377 -1982
rect 7762 -2054 7833 -1982
rect 8236 -2054 8307 -1982
rect 8692 -2054 8763 -1982
rect 9150 -2054 9221 -1982
rect 9606 -2054 9677 -1982
rect 10062 -2054 10133 -1982
rect 10520 -2054 10591 -1982
rect 10976 -2054 11047 -1982
rect 11432 -2054 11503 -1982
rect 11890 -2054 11961 -1982
rect 12346 -2054 12417 -1982
rect 12802 -2054 12873 -1982
rect 13260 -2054 13331 -1982
rect 13716 -2054 13787 -1982
rect 14172 -2054 14243 -1982
rect 14630 -2054 14701 -1982
rect 66 -2064 400 -2054
rect 0 -2124 10 -2064
rect 70 -2124 330 -2064
rect 390 -2124 400 -2064
rect 0 -2414 14 -2124
rect 66 -2414 400 -2124
rect 0 -2474 10 -2414
rect 70 -2474 330 -2414
rect 390 -2474 400 -2414
rect 0 -2556 14 -2474
rect 66 -2484 400 -2474
rect 456 -2064 856 -2054
rect 456 -2124 466 -2064
rect 526 -2124 786 -2064
rect 846 -2124 856 -2064
rect 456 -2234 856 -2124
rect 912 -2064 1312 -2054
rect 912 -2124 922 -2064
rect 982 -2124 1242 -2064
rect 1302 -2124 1312 -2064
rect 912 -2234 1312 -2124
rect 1370 -2064 1770 -2054
rect 1370 -2124 1380 -2064
rect 1440 -2124 1700 -2064
rect 1760 -2124 1770 -2064
rect 1370 -2234 1770 -2124
rect 1826 -2064 2226 -2054
rect 1826 -2124 1836 -2064
rect 1896 -2124 2156 -2064
rect 2216 -2124 2226 -2064
rect 1826 -2234 2226 -2124
rect 2282 -2064 2682 -2054
rect 2282 -2124 2292 -2064
rect 2352 -2124 2612 -2064
rect 2672 -2124 2682 -2064
rect 2282 -2234 2682 -2124
rect 2740 -2064 3140 -2054
rect 2740 -2124 2750 -2064
rect 2810 -2124 3070 -2064
rect 3130 -2124 3140 -2064
rect 2740 -2234 3140 -2124
rect 3196 -2064 3596 -2054
rect 3196 -2124 3206 -2064
rect 3266 -2124 3526 -2064
rect 3586 -2124 3596 -2064
rect 3196 -2234 3596 -2124
rect 3652 -2064 4052 -2054
rect 3652 -2124 3662 -2064
rect 3722 -2124 3982 -2064
rect 4042 -2124 4052 -2064
rect 3652 -2234 4052 -2124
rect 4110 -2064 4510 -2054
rect 4110 -2124 4120 -2064
rect 4180 -2124 4440 -2064
rect 4500 -2124 4510 -2064
rect 4110 -2234 4510 -2124
rect 4566 -2064 4966 -2054
rect 4566 -2124 4576 -2064
rect 4636 -2124 4896 -2064
rect 4956 -2124 4966 -2064
rect 4566 -2234 4966 -2124
rect 5022 -2064 5422 -2054
rect 5022 -2124 5032 -2064
rect 5092 -2124 5352 -2064
rect 5412 -2124 5422 -2064
rect 5022 -2234 5422 -2124
rect 5480 -2064 5880 -2054
rect 5480 -2124 5490 -2064
rect 5550 -2124 5810 -2064
rect 5870 -2124 5880 -2064
rect 5480 -2234 5880 -2124
rect 5936 -2064 6336 -2054
rect 5936 -2124 5946 -2064
rect 6006 -2124 6266 -2064
rect 6326 -2124 6336 -2064
rect 5936 -2234 6336 -2124
rect 6392 -2064 6792 -2054
rect 6392 -2124 6402 -2064
rect 6462 -2124 6722 -2064
rect 6782 -2124 6792 -2064
rect 6392 -2234 6792 -2124
rect 6850 -2064 7250 -2054
rect 6850 -2124 6860 -2064
rect 6920 -2124 7180 -2064
rect 7240 -2124 7250 -2064
rect 6850 -2234 7250 -2124
rect 7306 -2064 7706 -2054
rect 7306 -2124 7316 -2064
rect 7376 -2124 7636 -2064
rect 7696 -2124 7706 -2064
rect 7306 -2234 7706 -2124
rect 7762 -2064 8162 -2054
rect 7762 -2124 7772 -2064
rect 7832 -2124 8092 -2064
rect 8152 -2124 8162 -2064
rect 7762 -2234 8162 -2124
rect 8236 -2064 8636 -2054
rect 8236 -2124 8246 -2064
rect 8306 -2124 8566 -2064
rect 8626 -2124 8636 -2064
rect 8236 -2234 8636 -2124
rect 8692 -2064 9092 -2054
rect 8692 -2124 8702 -2064
rect 8762 -2124 9022 -2064
rect 9082 -2124 9092 -2064
rect 8692 -2234 9092 -2124
rect 9150 -2064 9550 -2054
rect 9150 -2124 9160 -2064
rect 9220 -2124 9480 -2064
rect 9540 -2124 9550 -2064
rect 9150 -2234 9550 -2124
rect 9606 -2064 10006 -2054
rect 9606 -2124 9616 -2064
rect 9676 -2124 9936 -2064
rect 9996 -2124 10006 -2064
rect 9606 -2234 10006 -2124
rect 10062 -2064 10462 -2054
rect 10062 -2124 10072 -2064
rect 10132 -2124 10392 -2064
rect 10452 -2124 10462 -2064
rect 10062 -2234 10462 -2124
rect 10520 -2064 10920 -2054
rect 10520 -2124 10530 -2064
rect 10590 -2124 10850 -2064
rect 10910 -2124 10920 -2064
rect 10520 -2234 10920 -2124
rect 10976 -2064 11376 -2054
rect 10976 -2124 10986 -2064
rect 11046 -2124 11306 -2064
rect 11366 -2124 11376 -2064
rect 10976 -2234 11376 -2124
rect 11432 -2064 11832 -2054
rect 11432 -2124 11442 -2064
rect 11502 -2124 11762 -2064
rect 11822 -2124 11832 -2064
rect 11432 -2234 11832 -2124
rect 11890 -2064 12290 -2054
rect 11890 -2124 11900 -2064
rect 11960 -2124 12220 -2064
rect 12280 -2124 12290 -2064
rect 11890 -2234 12290 -2124
rect 12346 -2064 12746 -2054
rect 12346 -2124 12356 -2064
rect 12416 -2124 12676 -2064
rect 12736 -2124 12746 -2064
rect 12346 -2234 12746 -2124
rect 12802 -2064 13202 -2054
rect 12802 -2124 12812 -2064
rect 12872 -2124 13132 -2064
rect 13192 -2124 13202 -2064
rect 12802 -2234 13202 -2124
rect 13260 -2064 13660 -2054
rect 13260 -2124 13270 -2064
rect 13330 -2124 13590 -2064
rect 13650 -2124 13660 -2064
rect 13260 -2234 13660 -2124
rect 13716 -2064 14116 -2054
rect 13716 -2124 13726 -2064
rect 13786 -2124 14046 -2064
rect 14106 -2124 14116 -2064
rect 13716 -2234 14116 -2124
rect 14172 -2064 14572 -2054
rect 14172 -2124 14182 -2064
rect 14242 -2124 14502 -2064
rect 14562 -2124 14572 -2064
rect 14172 -2234 14572 -2124
rect 14630 -2064 15030 -2054
rect 14630 -2124 14640 -2064
rect 14700 -2124 14960 -2064
rect 15020 -2124 15030 -2064
rect 14630 -2234 15030 -2124
rect 15086 -2064 15486 -2054
rect 15086 -2124 15096 -2064
rect 15156 -2124 15416 -2064
rect 15476 -2124 15486 -2064
rect 15086 -2234 15486 -2124
rect 456 -2304 15486 -2234
rect 456 -2414 856 -2304
rect 456 -2474 466 -2414
rect 526 -2474 786 -2414
rect 846 -2474 856 -2414
rect 456 -2484 856 -2474
rect 912 -2414 1312 -2304
rect 912 -2474 922 -2414
rect 982 -2474 1242 -2414
rect 1302 -2474 1312 -2414
rect 912 -2484 1312 -2474
rect 1370 -2414 1770 -2304
rect 1370 -2474 1380 -2414
rect 1440 -2474 1700 -2414
rect 1760 -2474 1770 -2414
rect 1370 -2484 1770 -2474
rect 1826 -2414 2226 -2304
rect 1826 -2474 1836 -2414
rect 1896 -2474 2156 -2414
rect 2216 -2474 2226 -2414
rect 1826 -2484 2226 -2474
rect 2282 -2414 2682 -2304
rect 2282 -2474 2292 -2414
rect 2352 -2474 2612 -2414
rect 2672 -2474 2682 -2414
rect 2282 -2484 2682 -2474
rect 2740 -2414 3140 -2304
rect 2740 -2474 2750 -2414
rect 2810 -2474 3070 -2414
rect 3130 -2474 3140 -2414
rect 2740 -2484 3140 -2474
rect 3196 -2414 3596 -2304
rect 3196 -2474 3206 -2414
rect 3266 -2474 3526 -2414
rect 3586 -2474 3596 -2414
rect 3196 -2484 3596 -2474
rect 3652 -2414 4052 -2304
rect 3652 -2474 3662 -2414
rect 3722 -2474 3982 -2414
rect 4042 -2474 4052 -2414
rect 3652 -2484 4052 -2474
rect 4110 -2414 4510 -2304
rect 4110 -2474 4120 -2414
rect 4180 -2474 4440 -2414
rect 4500 -2474 4510 -2414
rect 4110 -2484 4510 -2474
rect 4566 -2414 4966 -2304
rect 4566 -2474 4576 -2414
rect 4636 -2474 4896 -2414
rect 4956 -2474 4966 -2414
rect 4566 -2484 4966 -2474
rect 5022 -2414 5422 -2304
rect 5022 -2474 5032 -2414
rect 5092 -2474 5352 -2414
rect 5412 -2474 5422 -2414
rect 5022 -2484 5422 -2474
rect 5480 -2414 5880 -2304
rect 5480 -2474 5490 -2414
rect 5550 -2474 5810 -2414
rect 5870 -2474 5880 -2414
rect 5480 -2484 5880 -2474
rect 5936 -2414 6336 -2304
rect 5936 -2474 5946 -2414
rect 6006 -2474 6266 -2414
rect 6326 -2474 6336 -2414
rect 5936 -2484 6336 -2474
rect 6392 -2414 6792 -2304
rect 6392 -2474 6402 -2414
rect 6462 -2474 6722 -2414
rect 6782 -2474 6792 -2414
rect 6392 -2484 6792 -2474
rect 6850 -2414 7250 -2304
rect 6850 -2474 6860 -2414
rect 6920 -2474 7180 -2414
rect 7240 -2474 7250 -2414
rect 6850 -2484 7250 -2474
rect 7306 -2414 7706 -2304
rect 7306 -2474 7316 -2414
rect 7376 -2474 7636 -2414
rect 7696 -2474 7706 -2414
rect 7306 -2484 7706 -2474
rect 7762 -2414 8162 -2304
rect 7762 -2474 7772 -2414
rect 7832 -2474 8092 -2414
rect 8152 -2474 8162 -2414
rect 7762 -2484 8162 -2474
rect 8236 -2414 8636 -2304
rect 8236 -2474 8246 -2414
rect 8306 -2474 8566 -2414
rect 8626 -2474 8636 -2414
rect 8236 -2484 8636 -2474
rect 8692 -2414 9092 -2304
rect 8692 -2474 8702 -2414
rect 8762 -2474 9022 -2414
rect 9082 -2474 9092 -2414
rect 8692 -2484 9092 -2474
rect 9150 -2414 9550 -2304
rect 9150 -2474 9160 -2414
rect 9220 -2474 9480 -2414
rect 9540 -2474 9550 -2414
rect 9150 -2484 9550 -2474
rect 9606 -2414 10006 -2304
rect 9606 -2474 9616 -2414
rect 9676 -2474 9936 -2414
rect 9996 -2474 10006 -2414
rect 9606 -2484 10006 -2474
rect 10062 -2414 10462 -2304
rect 10062 -2474 10072 -2414
rect 10132 -2474 10392 -2414
rect 10452 -2474 10462 -2414
rect 10062 -2484 10462 -2474
rect 10520 -2414 10920 -2304
rect 10520 -2474 10530 -2414
rect 10590 -2474 10850 -2414
rect 10910 -2474 10920 -2414
rect 10520 -2484 10920 -2474
rect 10976 -2414 11376 -2304
rect 10976 -2474 10986 -2414
rect 11046 -2474 11306 -2414
rect 11366 -2474 11376 -2414
rect 10976 -2484 11376 -2474
rect 11432 -2414 11832 -2304
rect 11432 -2474 11442 -2414
rect 11502 -2474 11762 -2414
rect 11822 -2474 11832 -2414
rect 11432 -2484 11832 -2474
rect 11890 -2414 12290 -2304
rect 11890 -2474 11900 -2414
rect 11960 -2474 12220 -2414
rect 12280 -2474 12290 -2414
rect 11890 -2484 12290 -2474
rect 12346 -2414 12746 -2304
rect 12346 -2474 12356 -2414
rect 12416 -2474 12676 -2414
rect 12736 -2474 12746 -2414
rect 12346 -2484 12746 -2474
rect 12802 -2414 13202 -2304
rect 12802 -2474 12812 -2414
rect 12872 -2474 13132 -2414
rect 13192 -2474 13202 -2414
rect 12802 -2484 13202 -2474
rect 13260 -2414 13660 -2304
rect 13260 -2474 13270 -2414
rect 13330 -2474 13590 -2414
rect 13650 -2474 13660 -2414
rect 13260 -2484 13660 -2474
rect 13716 -2414 14116 -2304
rect 13716 -2474 13726 -2414
rect 13786 -2474 14046 -2414
rect 14106 -2474 14116 -2414
rect 13716 -2484 14116 -2474
rect 14172 -2414 14572 -2304
rect 14172 -2474 14182 -2414
rect 14242 -2474 14502 -2414
rect 14562 -2474 14572 -2414
rect 14172 -2484 14572 -2474
rect 14630 -2414 15030 -2304
rect 14630 -2474 14640 -2414
rect 14700 -2474 14960 -2414
rect 15020 -2474 15030 -2414
rect 14630 -2484 15030 -2474
rect 15086 -2414 15486 -2304
rect 15086 -2474 15096 -2414
rect 15156 -2474 15416 -2414
rect 15476 -2474 15486 -2414
rect 15086 -2484 15486 -2474
rect 66 -2546 80 -2484
rect 456 -2546 527 -2484
rect 912 -2546 983 -2484
rect 1370 -2546 1441 -2484
rect 1826 -2546 1897 -2484
rect 2282 -2546 2353 -2484
rect 2740 -2546 2810 -2484
rect 3196 -2546 3266 -2484
rect 3652 -2546 3722 -2484
rect 4110 -2546 4180 -2484
rect 4566 -2546 4636 -2484
rect 5022 -2546 5092 -2484
rect 5480 -2546 5550 -2484
rect 5936 -2546 6006 -2484
rect 6392 -2546 6462 -2484
rect 6850 -2546 6920 -2484
rect 7306 -2546 7376 -2484
rect 7762 -2546 7832 -2484
rect 8236 -2546 8306 -2484
rect 8692 -2546 8762 -2484
rect 9150 -2546 9220 -2484
rect 9606 -2546 9676 -2484
rect 10062 -2546 10132 -2484
rect 10520 -2546 10590 -2484
rect 10976 -2546 11046 -2484
rect 11432 -2546 11502 -2484
rect 11890 -2546 11960 -2484
rect 12346 -2546 12416 -2484
rect 12802 -2546 12872 -2484
rect 13260 -2546 13330 -2484
rect 13716 -2546 13786 -2484
rect 14172 -2546 14242 -2484
rect 14630 -2546 14700 -2484
rect 66 -2556 400 -2546
rect 0 -2616 10 -2556
rect 70 -2616 330 -2556
rect 390 -2616 400 -2556
rect 0 -2906 14 -2616
rect 66 -2906 400 -2616
rect 0 -2966 10 -2906
rect 70 -2966 330 -2906
rect 390 -2966 400 -2906
rect 0 -3552 14 -2966
rect 66 -2976 400 -2966
rect 456 -2556 856 -2546
rect 456 -2616 466 -2556
rect 526 -2616 786 -2556
rect 846 -2616 856 -2556
rect 456 -2726 856 -2616
rect 912 -2556 1312 -2546
rect 912 -2616 922 -2556
rect 982 -2616 1242 -2556
rect 1302 -2616 1312 -2556
rect 912 -2726 1312 -2616
rect 1370 -2556 1770 -2546
rect 1370 -2616 1380 -2556
rect 1440 -2616 1700 -2556
rect 1760 -2616 1770 -2556
rect 1370 -2726 1770 -2616
rect 1826 -2556 2226 -2546
rect 1826 -2616 1836 -2556
rect 1896 -2616 2156 -2556
rect 2216 -2616 2226 -2556
rect 1826 -2726 2226 -2616
rect 2282 -2556 2682 -2546
rect 2282 -2616 2292 -2556
rect 2352 -2616 2612 -2556
rect 2672 -2616 2682 -2556
rect 2282 -2726 2682 -2616
rect 2740 -2556 3140 -2546
rect 2740 -2616 2750 -2556
rect 2810 -2616 3070 -2556
rect 3130 -2616 3140 -2556
rect 2740 -2726 3140 -2616
rect 3196 -2556 3596 -2546
rect 3196 -2616 3206 -2556
rect 3266 -2616 3526 -2556
rect 3586 -2616 3596 -2556
rect 3196 -2726 3596 -2616
rect 3652 -2556 4052 -2546
rect 3652 -2616 3662 -2556
rect 3722 -2616 3982 -2556
rect 4042 -2616 4052 -2556
rect 3652 -2726 4052 -2616
rect 4110 -2556 4510 -2546
rect 4110 -2616 4120 -2556
rect 4180 -2616 4440 -2556
rect 4500 -2616 4510 -2556
rect 4110 -2726 4510 -2616
rect 4566 -2556 4966 -2546
rect 4566 -2616 4576 -2556
rect 4636 -2616 4896 -2556
rect 4956 -2616 4966 -2556
rect 4566 -2726 4966 -2616
rect 5022 -2556 5422 -2546
rect 5022 -2616 5032 -2556
rect 5092 -2616 5352 -2556
rect 5412 -2616 5422 -2556
rect 5022 -2726 5422 -2616
rect 5480 -2556 5880 -2546
rect 5480 -2616 5490 -2556
rect 5550 -2616 5810 -2556
rect 5870 -2616 5880 -2556
rect 5480 -2726 5880 -2616
rect 5936 -2556 6336 -2546
rect 5936 -2616 5946 -2556
rect 6006 -2616 6266 -2556
rect 6326 -2616 6336 -2556
rect 5936 -2726 6336 -2616
rect 6392 -2556 6792 -2546
rect 6392 -2616 6402 -2556
rect 6462 -2616 6722 -2556
rect 6782 -2616 6792 -2556
rect 6392 -2726 6792 -2616
rect 6850 -2556 7250 -2546
rect 6850 -2616 6860 -2556
rect 6920 -2616 7180 -2556
rect 7240 -2616 7250 -2556
rect 6850 -2726 7250 -2616
rect 7306 -2556 7706 -2546
rect 7306 -2616 7316 -2556
rect 7376 -2616 7636 -2556
rect 7696 -2616 7706 -2556
rect 7306 -2726 7706 -2616
rect 7762 -2556 8162 -2546
rect 7762 -2616 7772 -2556
rect 7832 -2616 8092 -2556
rect 8152 -2616 8162 -2556
rect 7762 -2726 8162 -2616
rect 8236 -2556 8636 -2546
rect 8236 -2616 8246 -2556
rect 8306 -2616 8566 -2556
rect 8626 -2616 8636 -2556
rect 8236 -2726 8636 -2616
rect 8692 -2556 9092 -2546
rect 8692 -2616 8702 -2556
rect 8762 -2616 9022 -2556
rect 9082 -2616 9092 -2556
rect 8692 -2726 9092 -2616
rect 9150 -2556 9550 -2546
rect 9150 -2616 9160 -2556
rect 9220 -2616 9480 -2556
rect 9540 -2616 9550 -2556
rect 9150 -2726 9550 -2616
rect 9606 -2556 10006 -2546
rect 9606 -2616 9616 -2556
rect 9676 -2616 9936 -2556
rect 9996 -2616 10006 -2556
rect 9606 -2726 10006 -2616
rect 10062 -2556 10462 -2546
rect 10062 -2616 10072 -2556
rect 10132 -2616 10392 -2556
rect 10452 -2616 10462 -2556
rect 10062 -2726 10462 -2616
rect 10520 -2556 10920 -2546
rect 10520 -2616 10530 -2556
rect 10590 -2616 10850 -2556
rect 10910 -2616 10920 -2556
rect 10520 -2726 10920 -2616
rect 10976 -2556 11376 -2546
rect 10976 -2616 10986 -2556
rect 11046 -2616 11306 -2556
rect 11366 -2616 11376 -2556
rect 10976 -2726 11376 -2616
rect 11432 -2556 11832 -2546
rect 11432 -2616 11442 -2556
rect 11502 -2616 11762 -2556
rect 11822 -2616 11832 -2556
rect 11432 -2726 11832 -2616
rect 11890 -2556 12290 -2546
rect 11890 -2616 11900 -2556
rect 11960 -2616 12220 -2556
rect 12280 -2616 12290 -2556
rect 11890 -2726 12290 -2616
rect 12346 -2556 12746 -2546
rect 12346 -2616 12356 -2556
rect 12416 -2616 12676 -2556
rect 12736 -2616 12746 -2556
rect 12346 -2726 12746 -2616
rect 12802 -2556 13202 -2546
rect 12802 -2616 12812 -2556
rect 12872 -2616 13132 -2556
rect 13192 -2616 13202 -2556
rect 12802 -2726 13202 -2616
rect 13260 -2556 13660 -2546
rect 13260 -2616 13270 -2556
rect 13330 -2616 13590 -2556
rect 13650 -2616 13660 -2556
rect 13260 -2726 13660 -2616
rect 13716 -2556 14116 -2546
rect 13716 -2616 13726 -2556
rect 13786 -2616 14046 -2556
rect 14106 -2616 14116 -2556
rect 13716 -2726 14116 -2616
rect 14172 -2556 14572 -2546
rect 14172 -2616 14182 -2556
rect 14242 -2616 14502 -2556
rect 14562 -2616 14572 -2556
rect 14172 -2726 14572 -2616
rect 14630 -2556 15030 -2546
rect 14630 -2616 14640 -2556
rect 14700 -2616 14960 -2556
rect 15020 -2616 15030 -2556
rect 14630 -2726 15030 -2616
rect 15086 -2556 15486 -2546
rect 15086 -2616 15096 -2556
rect 15156 -2616 15416 -2556
rect 15476 -2616 15486 -2556
rect 15086 -2726 15486 -2616
rect 456 -2796 15486 -2726
rect 456 -2906 856 -2796
rect 456 -2966 466 -2906
rect 526 -2966 786 -2906
rect 846 -2966 856 -2906
rect 456 -2976 856 -2966
rect 912 -2906 1312 -2796
rect 912 -2966 922 -2906
rect 982 -2966 1242 -2906
rect 1302 -2966 1312 -2906
rect 912 -2976 1312 -2966
rect 1370 -2906 1770 -2796
rect 1370 -2966 1380 -2906
rect 1440 -2966 1700 -2906
rect 1760 -2966 1770 -2906
rect 1370 -2976 1770 -2966
rect 1826 -2906 2226 -2796
rect 1826 -2966 1836 -2906
rect 1896 -2966 2156 -2906
rect 2216 -2966 2226 -2906
rect 1826 -2976 2226 -2966
rect 2282 -2906 2682 -2796
rect 2282 -2966 2292 -2906
rect 2352 -2966 2612 -2906
rect 2672 -2966 2682 -2906
rect 2282 -2976 2682 -2966
rect 2740 -2906 3140 -2796
rect 2740 -2966 2750 -2906
rect 2810 -2966 3070 -2906
rect 3130 -2966 3140 -2906
rect 2740 -2976 3140 -2966
rect 3196 -2906 3596 -2796
rect 3196 -2966 3206 -2906
rect 3266 -2966 3526 -2906
rect 3586 -2966 3596 -2906
rect 3196 -2976 3596 -2966
rect 3652 -2906 4052 -2796
rect 3652 -2966 3662 -2906
rect 3722 -2966 3982 -2906
rect 4042 -2966 4052 -2906
rect 3652 -2976 4052 -2966
rect 4110 -2906 4510 -2796
rect 4110 -2966 4120 -2906
rect 4180 -2966 4440 -2906
rect 4500 -2966 4510 -2906
rect 4110 -2976 4510 -2966
rect 4566 -2906 4966 -2796
rect 4566 -2966 4576 -2906
rect 4636 -2966 4896 -2906
rect 4956 -2966 4966 -2906
rect 4566 -2976 4966 -2966
rect 5022 -2906 5422 -2796
rect 5022 -2966 5032 -2906
rect 5092 -2966 5352 -2906
rect 5412 -2966 5422 -2906
rect 5022 -2976 5422 -2966
rect 5480 -2906 5880 -2796
rect 5480 -2966 5490 -2906
rect 5550 -2966 5810 -2906
rect 5870 -2966 5880 -2906
rect 5480 -2976 5880 -2966
rect 5936 -2906 6336 -2796
rect 5936 -2966 5946 -2906
rect 6006 -2966 6266 -2906
rect 6326 -2966 6336 -2906
rect 5936 -2976 6336 -2966
rect 6392 -2906 6792 -2796
rect 6392 -2966 6402 -2906
rect 6462 -2966 6722 -2906
rect 6782 -2966 6792 -2906
rect 6392 -2976 6792 -2966
rect 6850 -2906 7250 -2796
rect 6850 -2966 6860 -2906
rect 6920 -2966 7180 -2906
rect 7240 -2966 7250 -2906
rect 6850 -2976 7250 -2966
rect 7306 -2906 7706 -2796
rect 7306 -2966 7316 -2906
rect 7376 -2966 7636 -2906
rect 7696 -2966 7706 -2906
rect 7306 -2976 7706 -2966
rect 7762 -2906 8162 -2796
rect 7762 -2966 7772 -2906
rect 7832 -2966 8092 -2906
rect 8152 -2966 8162 -2906
rect 7762 -2976 8162 -2966
rect 8236 -2906 8636 -2796
rect 8236 -2966 8246 -2906
rect 8306 -2966 8566 -2906
rect 8626 -2966 8636 -2906
rect 8236 -2976 8636 -2966
rect 8692 -2906 9092 -2796
rect 8692 -2966 8702 -2906
rect 8762 -2966 9022 -2906
rect 9082 -2966 9092 -2906
rect 8692 -2976 9092 -2966
rect 9150 -2906 9550 -2796
rect 9150 -2966 9160 -2906
rect 9220 -2966 9480 -2906
rect 9540 -2966 9550 -2906
rect 9150 -2976 9550 -2966
rect 9606 -2906 10006 -2796
rect 9606 -2966 9616 -2906
rect 9676 -2966 9936 -2906
rect 9996 -2966 10006 -2906
rect 9606 -2976 10006 -2966
rect 10062 -2906 10462 -2796
rect 10062 -2966 10072 -2906
rect 10132 -2966 10392 -2906
rect 10452 -2966 10462 -2906
rect 10062 -2976 10462 -2966
rect 10520 -2906 10920 -2796
rect 10520 -2966 10530 -2906
rect 10590 -2966 10850 -2906
rect 10910 -2966 10920 -2906
rect 10520 -2976 10920 -2966
rect 10976 -2906 11376 -2796
rect 10976 -2966 10986 -2906
rect 11046 -2966 11306 -2906
rect 11366 -2966 11376 -2906
rect 10976 -2976 11376 -2966
rect 11432 -2906 11832 -2796
rect 11432 -2966 11442 -2906
rect 11502 -2966 11762 -2906
rect 11822 -2966 11832 -2906
rect 11432 -2976 11832 -2966
rect 11890 -2906 12290 -2796
rect 11890 -2966 11900 -2906
rect 11960 -2966 12220 -2906
rect 12280 -2966 12290 -2906
rect 11890 -2976 12290 -2966
rect 12346 -2906 12746 -2796
rect 12346 -2966 12356 -2906
rect 12416 -2966 12676 -2906
rect 12736 -2966 12746 -2906
rect 12346 -2976 12746 -2966
rect 12802 -2906 13202 -2796
rect 12802 -2966 12812 -2906
rect 12872 -2966 13132 -2906
rect 13192 -2966 13202 -2906
rect 12802 -2976 13202 -2966
rect 13260 -2906 13660 -2796
rect 13260 -2966 13270 -2906
rect 13330 -2966 13590 -2906
rect 13650 -2966 13660 -2906
rect 13260 -2976 13660 -2966
rect 13716 -2906 14116 -2796
rect 13716 -2966 13726 -2906
rect 13786 -2966 14046 -2906
rect 14106 -2966 14116 -2906
rect 13716 -2976 14116 -2966
rect 14172 -2906 14572 -2796
rect 14172 -2966 14182 -2906
rect 14242 -2966 14502 -2906
rect 14562 -2966 14572 -2906
rect 14172 -2976 14572 -2966
rect 14630 -2906 15030 -2796
rect 14630 -2966 14640 -2906
rect 14700 -2966 14960 -2906
rect 15020 -2966 15030 -2906
rect 14630 -2976 15030 -2966
rect 15086 -2906 15486 -2796
rect 15086 -2966 15096 -2906
rect 15156 -2966 15416 -2906
rect 15476 -2966 15486 -2906
rect 15086 -2976 15486 -2966
rect 66 -3542 80 -2976
rect 456 -3049 526 -2976
rect 912 -3040 982 -2976
rect 1370 -3040 1440 -2976
rect 1826 -3041 1896 -2976
rect 2282 -3041 2352 -2976
rect 2740 -3041 2810 -2976
rect 3196 -3041 3266 -2976
rect 3652 -3040 3722 -2976
rect 4110 -3041 4180 -2976
rect 4566 -3041 4636 -2976
rect 5022 -3040 5092 -2976
rect 5480 -3041 5550 -2976
rect 5936 -3041 6006 -2976
rect 6392 -3041 6462 -2976
rect 6850 -3041 6920 -2976
rect 7306 -3041 7376 -2976
rect 7762 -3041 7832 -2976
rect 8236 -3041 8306 -2976
rect 8692 -3041 8762 -2976
rect 9150 -3041 9220 -2976
rect 9606 -3041 9676 -2976
rect 10062 -3041 10132 -2976
rect 10520 -3041 10590 -2976
rect 10976 -3042 11047 -2976
rect 11432 -3043 11503 -2976
rect 11890 -3042 11961 -2976
rect 12346 -3043 12417 -2976
rect 12802 -3042 12873 -2976
rect 13260 -3043 13331 -2976
rect 13716 -3043 13787 -2976
rect 14172 -3045 14243 -2976
rect 14630 -3047 14701 -2976
rect 340 -3289 400 -3219
rect 456 -3289 15250 -3219
rect 456 -3542 526 -3470
rect 912 -3542 983 -3470
rect 1370 -3542 1441 -3470
rect 1826 -3542 1897 -3470
rect 2282 -3542 2353 -3470
rect 2740 -3542 2811 -3470
rect 3196 -3542 3267 -3470
rect 3652 -3542 3723 -3470
rect 4110 -3542 4181 -3470
rect 4566 -3542 4637 -3470
rect 5022 -3542 5093 -3470
rect 5480 -3542 5551 -3470
rect 5936 -3542 6007 -3470
rect 6392 -3542 6463 -3470
rect 6850 -3542 6921 -3470
rect 7306 -3542 7377 -3470
rect 7762 -3542 7833 -3470
rect 8236 -3542 8307 -3470
rect 8692 -3542 8763 -3470
rect 9150 -3542 9221 -3470
rect 9606 -3542 9677 -3470
rect 10062 -3542 10133 -3470
rect 10520 -3542 10591 -3470
rect 10976 -3542 11047 -3470
rect 11432 -3542 11503 -3470
rect 11890 -3542 11961 -3470
rect 12346 -3542 12417 -3470
rect 12802 -3542 12873 -3470
rect 13260 -3542 13331 -3470
rect 13716 -3542 13787 -3470
rect 14172 -3542 14243 -3470
rect 14630 -3542 14701 -3470
rect 66 -3552 400 -3542
rect 0 -3612 10 -3552
rect 70 -3612 330 -3552
rect 390 -3612 400 -3552
rect 0 -3902 14 -3612
rect 66 -3902 400 -3612
rect 0 -3962 10 -3902
rect 70 -3962 330 -3902
rect 390 -3962 400 -3902
rect 0 -4044 14 -3962
rect 66 -3972 400 -3962
rect 456 -3552 856 -3542
rect 456 -3612 466 -3552
rect 526 -3612 786 -3552
rect 846 -3612 856 -3552
rect 456 -3722 856 -3612
rect 912 -3552 1312 -3542
rect 912 -3612 922 -3552
rect 982 -3612 1242 -3552
rect 1302 -3612 1312 -3552
rect 912 -3722 1312 -3612
rect 1370 -3552 1770 -3542
rect 1370 -3612 1380 -3552
rect 1440 -3612 1700 -3552
rect 1760 -3612 1770 -3552
rect 1370 -3722 1770 -3612
rect 1826 -3552 2226 -3542
rect 1826 -3612 1836 -3552
rect 1896 -3612 2156 -3552
rect 2216 -3612 2226 -3552
rect 1826 -3722 2226 -3612
rect 2282 -3552 2682 -3542
rect 2282 -3612 2292 -3552
rect 2352 -3612 2612 -3552
rect 2672 -3612 2682 -3552
rect 2282 -3722 2682 -3612
rect 2740 -3552 3140 -3542
rect 2740 -3612 2750 -3552
rect 2810 -3612 3070 -3552
rect 3130 -3612 3140 -3552
rect 2740 -3722 3140 -3612
rect 3196 -3552 3596 -3542
rect 3196 -3612 3206 -3552
rect 3266 -3612 3526 -3552
rect 3586 -3612 3596 -3552
rect 3196 -3722 3596 -3612
rect 3652 -3552 4052 -3542
rect 3652 -3612 3662 -3552
rect 3722 -3612 3982 -3552
rect 4042 -3612 4052 -3552
rect 3652 -3722 4052 -3612
rect 4110 -3552 4510 -3542
rect 4110 -3612 4120 -3552
rect 4180 -3612 4440 -3552
rect 4500 -3612 4510 -3552
rect 4110 -3722 4510 -3612
rect 4566 -3552 4966 -3542
rect 4566 -3612 4576 -3552
rect 4636 -3612 4896 -3552
rect 4956 -3612 4966 -3552
rect 4566 -3722 4966 -3612
rect 5022 -3552 5422 -3542
rect 5022 -3612 5032 -3552
rect 5092 -3612 5352 -3552
rect 5412 -3612 5422 -3552
rect 5022 -3722 5422 -3612
rect 5480 -3552 5880 -3542
rect 5480 -3612 5490 -3552
rect 5550 -3612 5810 -3552
rect 5870 -3612 5880 -3552
rect 5480 -3722 5880 -3612
rect 5936 -3552 6336 -3542
rect 5936 -3612 5946 -3552
rect 6006 -3612 6266 -3552
rect 6326 -3612 6336 -3552
rect 5936 -3722 6336 -3612
rect 6392 -3552 6792 -3542
rect 6392 -3612 6402 -3552
rect 6462 -3612 6722 -3552
rect 6782 -3612 6792 -3552
rect 6392 -3722 6792 -3612
rect 6850 -3552 7250 -3542
rect 6850 -3612 6860 -3552
rect 6920 -3612 7180 -3552
rect 7240 -3612 7250 -3552
rect 6850 -3722 7250 -3612
rect 7306 -3552 7706 -3542
rect 7306 -3612 7316 -3552
rect 7376 -3612 7636 -3552
rect 7696 -3612 7706 -3552
rect 7306 -3722 7706 -3612
rect 7762 -3552 8162 -3542
rect 7762 -3612 7772 -3552
rect 7832 -3612 8092 -3552
rect 8152 -3612 8162 -3552
rect 7762 -3722 8162 -3612
rect 8236 -3552 8636 -3542
rect 8236 -3612 8246 -3552
rect 8306 -3612 8566 -3552
rect 8626 -3612 8636 -3552
rect 8236 -3722 8636 -3612
rect 8692 -3552 9092 -3542
rect 8692 -3612 8702 -3552
rect 8762 -3612 9022 -3552
rect 9082 -3612 9092 -3552
rect 8692 -3722 9092 -3612
rect 9150 -3552 9550 -3542
rect 9150 -3612 9160 -3552
rect 9220 -3612 9480 -3552
rect 9540 -3612 9550 -3552
rect 9150 -3722 9550 -3612
rect 9606 -3552 10006 -3542
rect 9606 -3612 9616 -3552
rect 9676 -3612 9936 -3552
rect 9996 -3612 10006 -3552
rect 9606 -3722 10006 -3612
rect 10062 -3552 10462 -3542
rect 10062 -3612 10072 -3552
rect 10132 -3612 10392 -3552
rect 10452 -3612 10462 -3552
rect 10062 -3722 10462 -3612
rect 10520 -3552 10920 -3542
rect 10520 -3612 10530 -3552
rect 10590 -3612 10850 -3552
rect 10910 -3612 10920 -3552
rect 10520 -3722 10920 -3612
rect 10976 -3552 11376 -3542
rect 10976 -3612 10986 -3552
rect 11046 -3612 11306 -3552
rect 11366 -3612 11376 -3552
rect 10976 -3722 11376 -3612
rect 11432 -3552 11832 -3542
rect 11432 -3612 11442 -3552
rect 11502 -3612 11762 -3552
rect 11822 -3612 11832 -3552
rect 11432 -3722 11832 -3612
rect 11890 -3552 12290 -3542
rect 11890 -3612 11900 -3552
rect 11960 -3612 12220 -3552
rect 12280 -3612 12290 -3552
rect 11890 -3722 12290 -3612
rect 12346 -3552 12746 -3542
rect 12346 -3612 12356 -3552
rect 12416 -3612 12676 -3552
rect 12736 -3612 12746 -3552
rect 12346 -3722 12746 -3612
rect 12802 -3552 13202 -3542
rect 12802 -3612 12812 -3552
rect 12872 -3612 13132 -3552
rect 13192 -3612 13202 -3552
rect 12802 -3722 13202 -3612
rect 13260 -3552 13660 -3542
rect 13260 -3612 13270 -3552
rect 13330 -3612 13590 -3552
rect 13650 -3612 13660 -3552
rect 13260 -3722 13660 -3612
rect 13716 -3552 14116 -3542
rect 13716 -3612 13726 -3552
rect 13786 -3612 14046 -3552
rect 14106 -3612 14116 -3552
rect 13716 -3722 14116 -3612
rect 14172 -3552 14572 -3542
rect 14172 -3612 14182 -3552
rect 14242 -3612 14502 -3552
rect 14562 -3612 14572 -3552
rect 14172 -3722 14572 -3612
rect 14630 -3552 15030 -3542
rect 14630 -3612 14640 -3552
rect 14700 -3612 14960 -3552
rect 15020 -3612 15030 -3552
rect 14630 -3722 15030 -3612
rect 15086 -3552 15486 -3542
rect 15086 -3612 15096 -3552
rect 15156 -3612 15416 -3552
rect 15476 -3612 15486 -3552
rect 15086 -3722 15486 -3612
rect 456 -3792 15486 -3722
rect 456 -3902 856 -3792
rect 456 -3962 466 -3902
rect 526 -3962 786 -3902
rect 846 -3962 856 -3902
rect 456 -3972 856 -3962
rect 912 -3902 1312 -3792
rect 912 -3962 922 -3902
rect 982 -3962 1242 -3902
rect 1302 -3962 1312 -3902
rect 912 -3972 1312 -3962
rect 1370 -3902 1770 -3792
rect 1370 -3962 1380 -3902
rect 1440 -3962 1700 -3902
rect 1760 -3962 1770 -3902
rect 1370 -3972 1770 -3962
rect 1826 -3902 2226 -3792
rect 1826 -3962 1836 -3902
rect 1896 -3962 2156 -3902
rect 2216 -3962 2226 -3902
rect 1826 -3972 2226 -3962
rect 2282 -3902 2682 -3792
rect 2282 -3962 2292 -3902
rect 2352 -3962 2612 -3902
rect 2672 -3962 2682 -3902
rect 2282 -3972 2682 -3962
rect 2740 -3902 3140 -3792
rect 2740 -3962 2750 -3902
rect 2810 -3962 3070 -3902
rect 3130 -3962 3140 -3902
rect 2740 -3972 3140 -3962
rect 3196 -3902 3596 -3792
rect 3196 -3962 3206 -3902
rect 3266 -3962 3526 -3902
rect 3586 -3962 3596 -3902
rect 3196 -3972 3596 -3962
rect 3652 -3902 4052 -3792
rect 3652 -3962 3662 -3902
rect 3722 -3962 3982 -3902
rect 4042 -3962 4052 -3902
rect 3652 -3972 4052 -3962
rect 4110 -3902 4510 -3792
rect 4110 -3962 4120 -3902
rect 4180 -3962 4440 -3902
rect 4500 -3962 4510 -3902
rect 4110 -3972 4510 -3962
rect 4566 -3902 4966 -3792
rect 4566 -3962 4576 -3902
rect 4636 -3962 4896 -3902
rect 4956 -3962 4966 -3902
rect 4566 -3972 4966 -3962
rect 5022 -3902 5422 -3792
rect 5022 -3962 5032 -3902
rect 5092 -3962 5352 -3902
rect 5412 -3962 5422 -3902
rect 5022 -3972 5422 -3962
rect 5480 -3902 5880 -3792
rect 5480 -3962 5490 -3902
rect 5550 -3962 5810 -3902
rect 5870 -3962 5880 -3902
rect 5480 -3972 5880 -3962
rect 5936 -3902 6336 -3792
rect 5936 -3962 5946 -3902
rect 6006 -3962 6266 -3902
rect 6326 -3962 6336 -3902
rect 5936 -3972 6336 -3962
rect 6392 -3902 6792 -3792
rect 6392 -3962 6402 -3902
rect 6462 -3962 6722 -3902
rect 6782 -3962 6792 -3902
rect 6392 -3972 6792 -3962
rect 6850 -3902 7250 -3792
rect 6850 -3962 6860 -3902
rect 6920 -3962 7180 -3902
rect 7240 -3962 7250 -3902
rect 6850 -3972 7250 -3962
rect 7306 -3902 7706 -3792
rect 7306 -3962 7316 -3902
rect 7376 -3962 7636 -3902
rect 7696 -3962 7706 -3902
rect 7306 -3972 7706 -3962
rect 7762 -3902 8162 -3792
rect 7762 -3962 7772 -3902
rect 7832 -3962 8092 -3902
rect 8152 -3962 8162 -3902
rect 7762 -3972 8162 -3962
rect 8236 -3902 8636 -3792
rect 8236 -3962 8246 -3902
rect 8306 -3962 8566 -3902
rect 8626 -3962 8636 -3902
rect 8236 -3972 8636 -3962
rect 8692 -3902 9092 -3792
rect 8692 -3962 8702 -3902
rect 8762 -3962 9022 -3902
rect 9082 -3962 9092 -3902
rect 8692 -3972 9092 -3962
rect 9150 -3902 9550 -3792
rect 9150 -3962 9160 -3902
rect 9220 -3962 9480 -3902
rect 9540 -3962 9550 -3902
rect 9150 -3972 9550 -3962
rect 9606 -3902 10006 -3792
rect 9606 -3962 9616 -3902
rect 9676 -3962 9936 -3902
rect 9996 -3962 10006 -3902
rect 9606 -3972 10006 -3962
rect 10062 -3902 10462 -3792
rect 10062 -3962 10072 -3902
rect 10132 -3962 10392 -3902
rect 10452 -3962 10462 -3902
rect 10062 -3972 10462 -3962
rect 10520 -3902 10920 -3792
rect 10520 -3962 10530 -3902
rect 10590 -3962 10850 -3902
rect 10910 -3962 10920 -3902
rect 10520 -3972 10920 -3962
rect 10976 -3902 11376 -3792
rect 10976 -3962 10986 -3902
rect 11046 -3962 11306 -3902
rect 11366 -3962 11376 -3902
rect 10976 -3972 11376 -3962
rect 11432 -3902 11832 -3792
rect 11432 -3962 11442 -3902
rect 11502 -3962 11762 -3902
rect 11822 -3962 11832 -3902
rect 11432 -3972 11832 -3962
rect 11890 -3902 12290 -3792
rect 11890 -3962 11900 -3902
rect 11960 -3962 12220 -3902
rect 12280 -3962 12290 -3902
rect 11890 -3972 12290 -3962
rect 12346 -3902 12746 -3792
rect 12346 -3962 12356 -3902
rect 12416 -3962 12676 -3902
rect 12736 -3962 12746 -3902
rect 12346 -3972 12746 -3962
rect 12802 -3902 13202 -3792
rect 12802 -3962 12812 -3902
rect 12872 -3962 13132 -3902
rect 13192 -3962 13202 -3902
rect 12802 -3972 13202 -3962
rect 13260 -3902 13660 -3792
rect 13260 -3962 13270 -3902
rect 13330 -3962 13590 -3902
rect 13650 -3962 13660 -3902
rect 13260 -3972 13660 -3962
rect 13716 -3902 14116 -3792
rect 13716 -3962 13726 -3902
rect 13786 -3962 14046 -3902
rect 14106 -3962 14116 -3902
rect 13716 -3972 14116 -3962
rect 14172 -3902 14572 -3792
rect 14172 -3962 14182 -3902
rect 14242 -3962 14502 -3902
rect 14562 -3962 14572 -3902
rect 14172 -3972 14572 -3962
rect 14630 -3902 15030 -3792
rect 14630 -3962 14640 -3902
rect 14700 -3962 14960 -3902
rect 15020 -3962 15030 -3902
rect 14630 -3972 15030 -3962
rect 15086 -3902 15486 -3792
rect 15086 -3962 15096 -3902
rect 15156 -3962 15416 -3902
rect 15476 -3962 15486 -3902
rect 15086 -3972 15486 -3962
rect 66 -4034 80 -3972
rect 456 -4034 527 -3972
rect 912 -4034 983 -3972
rect 1370 -4034 1441 -3972
rect 1826 -4034 1897 -3972
rect 2282 -4034 2353 -3972
rect 2740 -4034 2810 -3972
rect 3196 -4034 3266 -3972
rect 3652 -4034 3722 -3972
rect 4110 -4034 4180 -3972
rect 4566 -4034 4636 -3972
rect 5022 -4034 5092 -3972
rect 5480 -4034 5550 -3972
rect 5936 -4034 6006 -3972
rect 6392 -4034 6462 -3972
rect 6850 -4034 6920 -3972
rect 7306 -4034 7376 -3972
rect 7762 -4034 7832 -3972
rect 8236 -4034 8306 -3972
rect 8692 -4034 8762 -3972
rect 9150 -4034 9220 -3972
rect 9606 -4034 9676 -3972
rect 10062 -4034 10132 -3972
rect 10520 -4034 10590 -3972
rect 10976 -4034 11046 -3972
rect 11432 -4034 11502 -3972
rect 11890 -4034 11960 -3972
rect 12346 -4034 12416 -3972
rect 12802 -4034 12872 -3972
rect 13260 -4034 13330 -3972
rect 13716 -4034 13786 -3972
rect 14172 -4034 14242 -3972
rect 14630 -4034 14700 -3972
rect 66 -4044 400 -4034
rect 0 -4104 10 -4044
rect 70 -4104 330 -4044
rect 390 -4104 400 -4044
rect 0 -4394 14 -4104
rect 66 -4394 400 -4104
rect 0 -4454 10 -4394
rect 70 -4454 330 -4394
rect 390 -4454 400 -4394
rect 0 -4560 14 -4454
rect 66 -4464 400 -4454
rect 456 -4044 856 -4034
rect 456 -4104 466 -4044
rect 526 -4104 786 -4044
rect 846 -4104 856 -4044
rect 456 -4214 856 -4104
rect 912 -4044 1312 -4034
rect 912 -4104 922 -4044
rect 982 -4104 1242 -4044
rect 1302 -4104 1312 -4044
rect 912 -4214 1312 -4104
rect 1370 -4044 1770 -4034
rect 1370 -4104 1380 -4044
rect 1440 -4104 1700 -4044
rect 1760 -4104 1770 -4044
rect 1370 -4214 1770 -4104
rect 1826 -4044 2226 -4034
rect 1826 -4104 1836 -4044
rect 1896 -4104 2156 -4044
rect 2216 -4104 2226 -4044
rect 1826 -4214 2226 -4104
rect 2282 -4044 2682 -4034
rect 2282 -4104 2292 -4044
rect 2352 -4104 2612 -4044
rect 2672 -4104 2682 -4044
rect 2282 -4214 2682 -4104
rect 2740 -4044 3140 -4034
rect 2740 -4104 2750 -4044
rect 2810 -4104 3070 -4044
rect 3130 -4104 3140 -4044
rect 2740 -4214 3140 -4104
rect 3196 -4044 3596 -4034
rect 3196 -4104 3206 -4044
rect 3266 -4104 3526 -4044
rect 3586 -4104 3596 -4044
rect 3196 -4214 3596 -4104
rect 3652 -4044 4052 -4034
rect 3652 -4104 3662 -4044
rect 3722 -4104 3982 -4044
rect 4042 -4104 4052 -4044
rect 3652 -4214 4052 -4104
rect 4110 -4044 4510 -4034
rect 4110 -4104 4120 -4044
rect 4180 -4104 4440 -4044
rect 4500 -4104 4510 -4044
rect 4110 -4214 4510 -4104
rect 4566 -4044 4966 -4034
rect 4566 -4104 4576 -4044
rect 4636 -4104 4896 -4044
rect 4956 -4104 4966 -4044
rect 4566 -4214 4966 -4104
rect 5022 -4044 5422 -4034
rect 5022 -4104 5032 -4044
rect 5092 -4104 5352 -4044
rect 5412 -4104 5422 -4044
rect 5022 -4214 5422 -4104
rect 5480 -4044 5880 -4034
rect 5480 -4104 5490 -4044
rect 5550 -4104 5810 -4044
rect 5870 -4104 5880 -4044
rect 5480 -4214 5880 -4104
rect 5936 -4044 6336 -4034
rect 5936 -4104 5946 -4044
rect 6006 -4104 6266 -4044
rect 6326 -4104 6336 -4044
rect 5936 -4214 6336 -4104
rect 6392 -4044 6792 -4034
rect 6392 -4104 6402 -4044
rect 6462 -4104 6722 -4044
rect 6782 -4104 6792 -4044
rect 6392 -4214 6792 -4104
rect 6850 -4044 7250 -4034
rect 6850 -4104 6860 -4044
rect 6920 -4104 7180 -4044
rect 7240 -4104 7250 -4044
rect 6850 -4214 7250 -4104
rect 7306 -4044 7706 -4034
rect 7306 -4104 7316 -4044
rect 7376 -4104 7636 -4044
rect 7696 -4104 7706 -4044
rect 7306 -4214 7706 -4104
rect 7762 -4044 8162 -4034
rect 7762 -4104 7772 -4044
rect 7832 -4104 8092 -4044
rect 8152 -4104 8162 -4044
rect 7762 -4214 8162 -4104
rect 8236 -4044 8636 -4034
rect 8236 -4104 8246 -4044
rect 8306 -4104 8566 -4044
rect 8626 -4104 8636 -4044
rect 8236 -4214 8636 -4104
rect 8692 -4044 9092 -4034
rect 8692 -4104 8702 -4044
rect 8762 -4104 9022 -4044
rect 9082 -4104 9092 -4044
rect 8692 -4214 9092 -4104
rect 9150 -4044 9550 -4034
rect 9150 -4104 9160 -4044
rect 9220 -4104 9480 -4044
rect 9540 -4104 9550 -4044
rect 9150 -4214 9550 -4104
rect 9606 -4044 10006 -4034
rect 9606 -4104 9616 -4044
rect 9676 -4104 9936 -4044
rect 9996 -4104 10006 -4044
rect 9606 -4214 10006 -4104
rect 10062 -4044 10462 -4034
rect 10062 -4104 10072 -4044
rect 10132 -4104 10392 -4044
rect 10452 -4104 10462 -4044
rect 10062 -4214 10462 -4104
rect 10520 -4044 10920 -4034
rect 10520 -4104 10530 -4044
rect 10590 -4104 10850 -4044
rect 10910 -4104 10920 -4044
rect 10520 -4214 10920 -4104
rect 10976 -4044 11376 -4034
rect 10976 -4104 10986 -4044
rect 11046 -4104 11306 -4044
rect 11366 -4104 11376 -4044
rect 10976 -4214 11376 -4104
rect 11432 -4044 11832 -4034
rect 11432 -4104 11442 -4044
rect 11502 -4104 11762 -4044
rect 11822 -4104 11832 -4044
rect 11432 -4214 11832 -4104
rect 11890 -4044 12290 -4034
rect 11890 -4104 11900 -4044
rect 11960 -4104 12220 -4044
rect 12280 -4104 12290 -4044
rect 11890 -4214 12290 -4104
rect 12346 -4044 12746 -4034
rect 12346 -4104 12356 -4044
rect 12416 -4104 12676 -4044
rect 12736 -4104 12746 -4044
rect 12346 -4214 12746 -4104
rect 12802 -4044 13202 -4034
rect 12802 -4104 12812 -4044
rect 12872 -4104 13132 -4044
rect 13192 -4104 13202 -4044
rect 12802 -4214 13202 -4104
rect 13260 -4044 13660 -4034
rect 13260 -4104 13270 -4044
rect 13330 -4104 13590 -4044
rect 13650 -4104 13660 -4044
rect 13260 -4214 13660 -4104
rect 13716 -4044 14116 -4034
rect 13716 -4104 13726 -4044
rect 13786 -4104 14046 -4044
rect 14106 -4104 14116 -4044
rect 13716 -4214 14116 -4104
rect 14172 -4044 14572 -4034
rect 14172 -4104 14182 -4044
rect 14242 -4104 14502 -4044
rect 14562 -4104 14572 -4044
rect 14172 -4214 14572 -4104
rect 14630 -4044 15030 -4034
rect 14630 -4104 14640 -4044
rect 14700 -4104 14960 -4044
rect 15020 -4104 15030 -4044
rect 14630 -4214 15030 -4104
rect 15086 -4044 15486 -4034
rect 15086 -4104 15096 -4044
rect 15156 -4104 15416 -4044
rect 15476 -4104 15486 -4044
rect 15086 -4214 15486 -4104
rect 456 -4284 15486 -4214
rect 456 -4394 856 -4284
rect 456 -4454 466 -4394
rect 526 -4454 786 -4394
rect 846 -4454 856 -4394
rect 456 -4464 856 -4454
rect 912 -4394 1312 -4284
rect 912 -4454 922 -4394
rect 982 -4454 1242 -4394
rect 1302 -4454 1312 -4394
rect 912 -4464 1312 -4454
rect 1370 -4394 1770 -4284
rect 1370 -4454 1380 -4394
rect 1440 -4454 1700 -4394
rect 1760 -4454 1770 -4394
rect 1370 -4464 1770 -4454
rect 1826 -4394 2226 -4284
rect 1826 -4454 1836 -4394
rect 1896 -4454 2156 -4394
rect 2216 -4454 2226 -4394
rect 1826 -4464 2226 -4454
rect 2282 -4394 2682 -4284
rect 2282 -4454 2292 -4394
rect 2352 -4454 2612 -4394
rect 2672 -4454 2682 -4394
rect 2282 -4464 2682 -4454
rect 2740 -4394 3140 -4284
rect 2740 -4454 2750 -4394
rect 2810 -4454 3070 -4394
rect 3130 -4454 3140 -4394
rect 2740 -4464 3140 -4454
rect 3196 -4394 3596 -4284
rect 3196 -4454 3206 -4394
rect 3266 -4454 3526 -4394
rect 3586 -4454 3596 -4394
rect 3196 -4464 3596 -4454
rect 3652 -4394 4052 -4284
rect 3652 -4454 3662 -4394
rect 3722 -4454 3982 -4394
rect 4042 -4454 4052 -4394
rect 3652 -4464 4052 -4454
rect 4110 -4394 4510 -4284
rect 4110 -4454 4120 -4394
rect 4180 -4454 4440 -4394
rect 4500 -4454 4510 -4394
rect 4110 -4464 4510 -4454
rect 4566 -4394 4966 -4284
rect 4566 -4454 4576 -4394
rect 4636 -4454 4896 -4394
rect 4956 -4454 4966 -4394
rect 4566 -4464 4966 -4454
rect 5022 -4394 5422 -4284
rect 5022 -4454 5032 -4394
rect 5092 -4454 5352 -4394
rect 5412 -4454 5422 -4394
rect 5022 -4464 5422 -4454
rect 5480 -4394 5880 -4284
rect 5480 -4454 5490 -4394
rect 5550 -4454 5810 -4394
rect 5870 -4454 5880 -4394
rect 5480 -4464 5880 -4454
rect 5936 -4394 6336 -4284
rect 5936 -4454 5946 -4394
rect 6006 -4454 6266 -4394
rect 6326 -4454 6336 -4394
rect 5936 -4464 6336 -4454
rect 6392 -4394 6792 -4284
rect 6392 -4454 6402 -4394
rect 6462 -4454 6722 -4394
rect 6782 -4454 6792 -4394
rect 6392 -4464 6792 -4454
rect 6850 -4394 7250 -4284
rect 6850 -4454 6860 -4394
rect 6920 -4454 7180 -4394
rect 7240 -4454 7250 -4394
rect 6850 -4464 7250 -4454
rect 7306 -4394 7706 -4284
rect 7306 -4454 7316 -4394
rect 7376 -4454 7636 -4394
rect 7696 -4454 7706 -4394
rect 7306 -4464 7706 -4454
rect 7762 -4394 8162 -4284
rect 7762 -4454 7772 -4394
rect 7832 -4454 8092 -4394
rect 8152 -4454 8162 -4394
rect 7762 -4464 8162 -4454
rect 8236 -4394 8636 -4284
rect 8236 -4454 8246 -4394
rect 8306 -4454 8566 -4394
rect 8626 -4454 8636 -4394
rect 8236 -4464 8636 -4454
rect 8692 -4394 9092 -4284
rect 8692 -4454 8702 -4394
rect 8762 -4454 9022 -4394
rect 9082 -4454 9092 -4394
rect 8692 -4464 9092 -4454
rect 9150 -4394 9550 -4284
rect 9150 -4454 9160 -4394
rect 9220 -4454 9480 -4394
rect 9540 -4454 9550 -4394
rect 9150 -4464 9550 -4454
rect 9606 -4394 10006 -4284
rect 9606 -4454 9616 -4394
rect 9676 -4454 9936 -4394
rect 9996 -4454 10006 -4394
rect 9606 -4464 10006 -4454
rect 10062 -4394 10462 -4284
rect 10062 -4454 10072 -4394
rect 10132 -4454 10392 -4394
rect 10452 -4454 10462 -4394
rect 10062 -4464 10462 -4454
rect 10520 -4394 10920 -4284
rect 10520 -4454 10530 -4394
rect 10590 -4454 10850 -4394
rect 10910 -4454 10920 -4394
rect 10520 -4464 10920 -4454
rect 10976 -4394 11376 -4284
rect 10976 -4454 10986 -4394
rect 11046 -4454 11306 -4394
rect 11366 -4454 11376 -4394
rect 10976 -4464 11376 -4454
rect 11432 -4394 11832 -4284
rect 11432 -4454 11442 -4394
rect 11502 -4454 11762 -4394
rect 11822 -4454 11832 -4394
rect 11432 -4464 11832 -4454
rect 11890 -4394 12290 -4284
rect 11890 -4454 11900 -4394
rect 11960 -4454 12220 -4394
rect 12280 -4454 12290 -4394
rect 11890 -4464 12290 -4454
rect 12346 -4394 12746 -4284
rect 12346 -4454 12356 -4394
rect 12416 -4454 12676 -4394
rect 12736 -4454 12746 -4394
rect 12346 -4464 12746 -4454
rect 12802 -4394 13202 -4284
rect 12802 -4454 12812 -4394
rect 12872 -4454 13132 -4394
rect 13192 -4454 13202 -4394
rect 12802 -4464 13202 -4454
rect 13260 -4394 13660 -4284
rect 13260 -4454 13270 -4394
rect 13330 -4454 13590 -4394
rect 13650 -4454 13660 -4394
rect 13260 -4464 13660 -4454
rect 13716 -4394 14116 -4284
rect 13716 -4454 13726 -4394
rect 13786 -4454 14046 -4394
rect 14106 -4454 14116 -4394
rect 13716 -4464 14116 -4454
rect 14172 -4394 14572 -4284
rect 14172 -4454 14182 -4394
rect 14242 -4454 14502 -4394
rect 14562 -4454 14572 -4394
rect 14172 -4464 14572 -4454
rect 14630 -4394 15030 -4284
rect 14630 -4454 14640 -4394
rect 14700 -4454 14960 -4394
rect 15020 -4454 15030 -4394
rect 14630 -4464 15030 -4454
rect 15086 -4394 15486 -4284
rect 15086 -4454 15096 -4394
rect 15156 -4454 15416 -4394
rect 15476 -4454 15486 -4394
rect 15086 -4464 15486 -4454
rect 66 -4550 80 -4464
rect 456 -4550 526 -4464
rect 912 -4550 982 -4464
rect 1370 -4550 1440 -4464
rect 1826 -4550 1896 -4464
rect 2282 -4550 2352 -4464
rect 2740 -4550 2810 -4464
rect 3196 -4550 3266 -4464
rect 3652 -4550 3722 -4464
rect 4110 -4550 4180 -4464
rect 4566 -4550 4636 -4464
rect 5022 -4550 5092 -4464
rect 5480 -4550 5550 -4464
rect 5936 -4550 6006 -4464
rect 6392 -4550 6462 -4464
rect 6850 -4550 6920 -4464
rect 7306 -4550 7376 -4464
rect 7762 -4550 7832 -4464
rect 8236 -4550 8306 -4464
rect 8692 -4550 8762 -4464
rect 9150 -4550 9220 -4464
rect 9606 -4550 9676 -4464
rect 10062 -4550 10132 -4464
rect 10520 -4550 10590 -4464
rect 10976 -4550 11046 -4464
rect 11432 -4550 11502 -4464
rect 11890 -4550 11960 -4464
rect 12346 -4550 12416 -4464
rect 12802 -4550 12872 -4464
rect 13260 -4550 13330 -4464
rect 13716 -4550 13786 -4464
rect 14172 -4550 14242 -4464
rect 14630 -4550 14700 -4464
rect 66 -4560 400 -4550
rect 0 -4620 10 -4560
rect 70 -4620 330 -4560
rect 390 -4620 400 -4560
rect 0 -4910 14 -4620
rect 66 -4910 400 -4620
rect 0 -4970 10 -4910
rect 70 -4970 330 -4910
rect 390 -4970 400 -4910
rect 0 -5062 14 -4970
rect 66 -4980 400 -4970
rect 456 -4560 856 -4550
rect 456 -4620 466 -4560
rect 526 -4620 786 -4560
rect 846 -4620 856 -4560
rect 456 -4730 856 -4620
rect 912 -4560 1312 -4550
rect 912 -4620 922 -4560
rect 982 -4620 1242 -4560
rect 1302 -4620 1312 -4560
rect 912 -4730 1312 -4620
rect 1370 -4560 1770 -4550
rect 1370 -4620 1380 -4560
rect 1440 -4620 1700 -4560
rect 1760 -4620 1770 -4560
rect 1370 -4730 1770 -4620
rect 1826 -4560 2226 -4550
rect 1826 -4620 1836 -4560
rect 1896 -4620 2156 -4560
rect 2216 -4620 2226 -4560
rect 1826 -4730 2226 -4620
rect 2282 -4560 2682 -4550
rect 2282 -4620 2292 -4560
rect 2352 -4620 2612 -4560
rect 2672 -4620 2682 -4560
rect 2282 -4730 2682 -4620
rect 2740 -4560 3140 -4550
rect 2740 -4620 2750 -4560
rect 2810 -4620 3070 -4560
rect 3130 -4620 3140 -4560
rect 2740 -4730 3140 -4620
rect 3196 -4560 3596 -4550
rect 3196 -4620 3206 -4560
rect 3266 -4620 3526 -4560
rect 3586 -4620 3596 -4560
rect 3196 -4730 3596 -4620
rect 3652 -4560 4052 -4550
rect 3652 -4620 3662 -4560
rect 3722 -4620 3982 -4560
rect 4042 -4620 4052 -4560
rect 3652 -4730 4052 -4620
rect 4110 -4560 4510 -4550
rect 4110 -4620 4120 -4560
rect 4180 -4620 4440 -4560
rect 4500 -4620 4510 -4560
rect 4110 -4730 4510 -4620
rect 4566 -4560 4966 -4550
rect 4566 -4620 4576 -4560
rect 4636 -4620 4896 -4560
rect 4956 -4620 4966 -4560
rect 4566 -4730 4966 -4620
rect 5022 -4560 5422 -4550
rect 5022 -4620 5032 -4560
rect 5092 -4620 5352 -4560
rect 5412 -4620 5422 -4560
rect 5022 -4730 5422 -4620
rect 5480 -4560 5880 -4550
rect 5480 -4620 5490 -4560
rect 5550 -4620 5810 -4560
rect 5870 -4620 5880 -4560
rect 5480 -4730 5880 -4620
rect 5936 -4560 6336 -4550
rect 5936 -4620 5946 -4560
rect 6006 -4620 6266 -4560
rect 6326 -4620 6336 -4560
rect 5936 -4730 6336 -4620
rect 6392 -4560 6792 -4550
rect 6392 -4620 6402 -4560
rect 6462 -4620 6722 -4560
rect 6782 -4620 6792 -4560
rect 6392 -4730 6792 -4620
rect 6850 -4560 7250 -4550
rect 6850 -4620 6860 -4560
rect 6920 -4620 7180 -4560
rect 7240 -4620 7250 -4560
rect 6850 -4730 7250 -4620
rect 7306 -4560 7706 -4550
rect 7306 -4620 7316 -4560
rect 7376 -4620 7636 -4560
rect 7696 -4620 7706 -4560
rect 7306 -4730 7706 -4620
rect 7762 -4560 8162 -4550
rect 7762 -4620 7772 -4560
rect 7832 -4620 8092 -4560
rect 8152 -4620 8162 -4560
rect 7762 -4730 8162 -4620
rect 8236 -4560 8636 -4550
rect 8236 -4620 8246 -4560
rect 8306 -4620 8566 -4560
rect 8626 -4620 8636 -4560
rect 8236 -4730 8636 -4620
rect 8692 -4560 9092 -4550
rect 8692 -4620 8702 -4560
rect 8762 -4620 9022 -4560
rect 9082 -4620 9092 -4560
rect 8692 -4730 9092 -4620
rect 9150 -4560 9550 -4550
rect 9150 -4620 9160 -4560
rect 9220 -4620 9480 -4560
rect 9540 -4620 9550 -4560
rect 9150 -4730 9550 -4620
rect 9606 -4560 10006 -4550
rect 9606 -4620 9616 -4560
rect 9676 -4620 9936 -4560
rect 9996 -4620 10006 -4560
rect 9606 -4730 10006 -4620
rect 10062 -4560 10462 -4550
rect 10062 -4620 10072 -4560
rect 10132 -4620 10392 -4560
rect 10452 -4620 10462 -4560
rect 10062 -4730 10462 -4620
rect 10520 -4560 10920 -4550
rect 10520 -4620 10530 -4560
rect 10590 -4620 10850 -4560
rect 10910 -4620 10920 -4560
rect 10520 -4730 10920 -4620
rect 10976 -4560 11376 -4550
rect 10976 -4620 10986 -4560
rect 11046 -4620 11306 -4560
rect 11366 -4620 11376 -4560
rect 10976 -4730 11376 -4620
rect 11432 -4560 11832 -4550
rect 11432 -4620 11442 -4560
rect 11502 -4620 11762 -4560
rect 11822 -4620 11832 -4560
rect 11432 -4730 11832 -4620
rect 11890 -4560 12290 -4550
rect 11890 -4620 11900 -4560
rect 11960 -4620 12220 -4560
rect 12280 -4620 12290 -4560
rect 11890 -4730 12290 -4620
rect 12346 -4560 12746 -4550
rect 12346 -4620 12356 -4560
rect 12416 -4620 12676 -4560
rect 12736 -4620 12746 -4560
rect 12346 -4730 12746 -4620
rect 12802 -4560 13202 -4550
rect 12802 -4620 12812 -4560
rect 12872 -4620 13132 -4560
rect 13192 -4620 13202 -4560
rect 12802 -4730 13202 -4620
rect 13260 -4560 13660 -4550
rect 13260 -4620 13270 -4560
rect 13330 -4620 13590 -4560
rect 13650 -4620 13660 -4560
rect 13260 -4730 13660 -4620
rect 13716 -4560 14116 -4550
rect 13716 -4620 13726 -4560
rect 13786 -4620 14046 -4560
rect 14106 -4620 14116 -4560
rect 13716 -4730 14116 -4620
rect 14172 -4560 14572 -4550
rect 14172 -4620 14182 -4560
rect 14242 -4620 14502 -4560
rect 14562 -4620 14572 -4560
rect 14172 -4730 14572 -4620
rect 14630 -4560 15030 -4550
rect 14630 -4620 14640 -4560
rect 14700 -4620 14960 -4560
rect 15020 -4620 15030 -4560
rect 14630 -4730 15030 -4620
rect 15086 -4560 15486 -4550
rect 15086 -4620 15096 -4560
rect 15156 -4620 15416 -4560
rect 15476 -4620 15486 -4560
rect 15086 -4730 15486 -4620
rect 456 -4800 15486 -4730
rect 456 -4910 856 -4800
rect 456 -4970 466 -4910
rect 526 -4970 786 -4910
rect 846 -4970 856 -4910
rect 456 -4980 856 -4970
rect 912 -4910 1312 -4800
rect 912 -4970 922 -4910
rect 982 -4970 1242 -4910
rect 1302 -4970 1312 -4910
rect 912 -4980 1312 -4970
rect 1370 -4910 1770 -4800
rect 1370 -4970 1380 -4910
rect 1440 -4970 1700 -4910
rect 1760 -4970 1770 -4910
rect 1370 -4980 1770 -4970
rect 1826 -4910 2226 -4800
rect 1826 -4970 1836 -4910
rect 1896 -4970 2156 -4910
rect 2216 -4970 2226 -4910
rect 1826 -4980 2226 -4970
rect 2282 -4910 2682 -4800
rect 2282 -4970 2292 -4910
rect 2352 -4970 2612 -4910
rect 2672 -4970 2682 -4910
rect 2282 -4980 2682 -4970
rect 2740 -4910 3140 -4800
rect 2740 -4970 2750 -4910
rect 2810 -4970 3070 -4910
rect 3130 -4970 3140 -4910
rect 2740 -4980 3140 -4970
rect 3196 -4910 3596 -4800
rect 3196 -4970 3206 -4910
rect 3266 -4970 3526 -4910
rect 3586 -4970 3596 -4910
rect 3196 -4980 3596 -4970
rect 3652 -4910 4052 -4800
rect 3652 -4970 3662 -4910
rect 3722 -4970 3982 -4910
rect 4042 -4970 4052 -4910
rect 3652 -4980 4052 -4970
rect 4110 -4910 4510 -4800
rect 4110 -4970 4120 -4910
rect 4180 -4970 4440 -4910
rect 4500 -4970 4510 -4910
rect 4110 -4980 4510 -4970
rect 4566 -4910 4966 -4800
rect 4566 -4970 4576 -4910
rect 4636 -4970 4896 -4910
rect 4956 -4970 4966 -4910
rect 4566 -4980 4966 -4970
rect 5022 -4910 5422 -4800
rect 5022 -4970 5032 -4910
rect 5092 -4970 5352 -4910
rect 5412 -4970 5422 -4910
rect 5022 -4980 5422 -4970
rect 5480 -4910 5880 -4800
rect 5480 -4970 5490 -4910
rect 5550 -4970 5810 -4910
rect 5870 -4970 5880 -4910
rect 5480 -4980 5880 -4970
rect 5936 -4910 6336 -4800
rect 5936 -4970 5946 -4910
rect 6006 -4970 6266 -4910
rect 6326 -4970 6336 -4910
rect 5936 -4980 6336 -4970
rect 6392 -4910 6792 -4800
rect 6392 -4970 6402 -4910
rect 6462 -4970 6722 -4910
rect 6782 -4970 6792 -4910
rect 6392 -4980 6792 -4970
rect 6850 -4910 7250 -4800
rect 6850 -4970 6860 -4910
rect 6920 -4970 7180 -4910
rect 7240 -4970 7250 -4910
rect 6850 -4980 7250 -4970
rect 7306 -4910 7706 -4800
rect 7306 -4970 7316 -4910
rect 7376 -4970 7636 -4910
rect 7696 -4970 7706 -4910
rect 7306 -4980 7706 -4970
rect 7762 -4910 8162 -4800
rect 7762 -4970 7772 -4910
rect 7832 -4970 8092 -4910
rect 8152 -4970 8162 -4910
rect 7762 -4980 8162 -4970
rect 8236 -4910 8636 -4800
rect 8236 -4970 8246 -4910
rect 8306 -4970 8566 -4910
rect 8626 -4970 8636 -4910
rect 8236 -4980 8636 -4970
rect 8692 -4910 9092 -4800
rect 8692 -4970 8702 -4910
rect 8762 -4970 9022 -4910
rect 9082 -4970 9092 -4910
rect 8692 -4980 9092 -4970
rect 9150 -4910 9550 -4800
rect 9150 -4970 9160 -4910
rect 9220 -4970 9480 -4910
rect 9540 -4970 9550 -4910
rect 9150 -4980 9550 -4970
rect 9606 -4910 10006 -4800
rect 9606 -4970 9616 -4910
rect 9676 -4970 9936 -4910
rect 9996 -4970 10006 -4910
rect 9606 -4980 10006 -4970
rect 10062 -4910 10462 -4800
rect 10062 -4970 10072 -4910
rect 10132 -4970 10392 -4910
rect 10452 -4970 10462 -4910
rect 10062 -4980 10462 -4970
rect 10520 -4910 10920 -4800
rect 10520 -4970 10530 -4910
rect 10590 -4970 10850 -4910
rect 10910 -4970 10920 -4910
rect 10520 -4980 10920 -4970
rect 10976 -4910 11376 -4800
rect 10976 -4970 10986 -4910
rect 11046 -4970 11306 -4910
rect 11366 -4970 11376 -4910
rect 10976 -4980 11376 -4970
rect 11432 -4910 11832 -4800
rect 11432 -4970 11442 -4910
rect 11502 -4970 11762 -4910
rect 11822 -4970 11832 -4910
rect 11432 -4980 11832 -4970
rect 11890 -4910 12290 -4800
rect 11890 -4970 11900 -4910
rect 11960 -4970 12220 -4910
rect 12280 -4970 12290 -4910
rect 11890 -4980 12290 -4970
rect 12346 -4910 12746 -4800
rect 12346 -4970 12356 -4910
rect 12416 -4970 12676 -4910
rect 12736 -4970 12746 -4910
rect 12346 -4980 12746 -4970
rect 12802 -4910 13202 -4800
rect 12802 -4970 12812 -4910
rect 12872 -4970 13132 -4910
rect 13192 -4970 13202 -4910
rect 12802 -4980 13202 -4970
rect 13260 -4910 13660 -4800
rect 13260 -4970 13270 -4910
rect 13330 -4970 13590 -4910
rect 13650 -4970 13660 -4910
rect 13260 -4980 13660 -4970
rect 13716 -4910 14116 -4800
rect 13716 -4970 13726 -4910
rect 13786 -4970 14046 -4910
rect 14106 -4970 14116 -4910
rect 13716 -4980 14116 -4970
rect 14172 -4910 14572 -4800
rect 14172 -4970 14182 -4910
rect 14242 -4970 14502 -4910
rect 14562 -4970 14572 -4910
rect 14172 -4980 14572 -4970
rect 14630 -4910 15030 -4800
rect 14630 -4970 14640 -4910
rect 14700 -4970 14960 -4910
rect 15020 -4970 15030 -4910
rect 14630 -4980 15030 -4970
rect 15086 -4910 15486 -4800
rect 15086 -4970 15096 -4910
rect 15156 -4970 15416 -4910
rect 15476 -4970 15486 -4910
rect 15086 -4980 15486 -4970
rect 66 -5052 80 -4980
rect 456 -5052 526 -4980
rect 912 -5052 983 -4980
rect 1370 -5052 1441 -4980
rect 1826 -5052 1897 -4980
rect 2282 -5052 2353 -4980
rect 2740 -5052 2811 -4980
rect 3196 -5052 3267 -4980
rect 3652 -5052 3723 -4980
rect 4110 -5052 4181 -4980
rect 4566 -5052 4637 -4980
rect 5022 -5052 5093 -4980
rect 5480 -5052 5551 -4980
rect 5936 -5052 6007 -4980
rect 6392 -5052 6463 -4980
rect 6850 -5052 6921 -4980
rect 7306 -5052 7377 -4980
rect 7762 -5052 7833 -4980
rect 8236 -5052 8307 -4980
rect 8692 -5052 8763 -4980
rect 9150 -5052 9221 -4980
rect 9606 -5052 9677 -4980
rect 10062 -5052 10133 -4980
rect 10520 -5052 10591 -4980
rect 10976 -5052 11047 -4980
rect 11432 -5052 11503 -4980
rect 11890 -5052 11961 -4980
rect 12346 -5052 12417 -4980
rect 12802 -5052 12873 -4980
rect 13260 -5052 13331 -4980
rect 13716 -5052 13787 -4980
rect 14172 -5052 14243 -4980
rect 14630 -5052 14701 -4980
rect 66 -5062 400 -5052
rect 0 -5122 10 -5062
rect 70 -5122 330 -5062
rect 390 -5122 400 -5062
rect 0 -5412 14 -5122
rect 66 -5412 400 -5122
rect 0 -5472 10 -5412
rect 70 -5472 330 -5412
rect 390 -5472 400 -5412
rect 0 -5554 14 -5472
rect 66 -5482 400 -5472
rect 456 -5062 856 -5052
rect 456 -5122 466 -5062
rect 526 -5122 786 -5062
rect 846 -5122 856 -5062
rect 456 -5232 856 -5122
rect 912 -5062 1312 -5052
rect 912 -5122 922 -5062
rect 982 -5122 1242 -5062
rect 1302 -5122 1312 -5062
rect 912 -5232 1312 -5122
rect 1370 -5062 1770 -5052
rect 1370 -5122 1380 -5062
rect 1440 -5122 1700 -5062
rect 1760 -5122 1770 -5062
rect 1370 -5232 1770 -5122
rect 1826 -5062 2226 -5052
rect 1826 -5122 1836 -5062
rect 1896 -5122 2156 -5062
rect 2216 -5122 2226 -5062
rect 1826 -5232 2226 -5122
rect 2282 -5062 2682 -5052
rect 2282 -5122 2292 -5062
rect 2352 -5122 2612 -5062
rect 2672 -5122 2682 -5062
rect 2282 -5232 2682 -5122
rect 456 -5233 2682 -5232
rect 2740 -5062 3140 -5052
rect 2740 -5122 2750 -5062
rect 2810 -5122 3070 -5062
rect 3130 -5122 3140 -5062
rect 2740 -5232 3140 -5122
rect 3196 -5062 3596 -5052
rect 3196 -5122 3206 -5062
rect 3266 -5122 3526 -5062
rect 3586 -5122 3596 -5062
rect 3196 -5232 3596 -5122
rect 3652 -5062 4052 -5052
rect 3652 -5122 3662 -5062
rect 3722 -5122 3982 -5062
rect 4042 -5122 4052 -5062
rect 3652 -5232 4052 -5122
rect 4110 -5062 4510 -5052
rect 4110 -5122 4120 -5062
rect 4180 -5122 4440 -5062
rect 4500 -5122 4510 -5062
rect 4110 -5232 4510 -5122
rect 4566 -5062 4966 -5052
rect 4566 -5122 4576 -5062
rect 4636 -5122 4896 -5062
rect 4956 -5122 4966 -5062
rect 4566 -5232 4966 -5122
rect 5022 -5062 5422 -5052
rect 5022 -5122 5032 -5062
rect 5092 -5122 5352 -5062
rect 5412 -5122 5422 -5062
rect 5022 -5232 5422 -5122
rect 5480 -5062 5880 -5052
rect 5480 -5122 5490 -5062
rect 5550 -5122 5810 -5062
rect 5870 -5122 5880 -5062
rect 5480 -5232 5880 -5122
rect 5936 -5062 6336 -5052
rect 5936 -5122 5946 -5062
rect 6006 -5122 6266 -5062
rect 6326 -5122 6336 -5062
rect 5936 -5232 6336 -5122
rect 6392 -5062 6792 -5052
rect 6392 -5122 6402 -5062
rect 6462 -5122 6722 -5062
rect 6782 -5122 6792 -5062
rect 6392 -5232 6792 -5122
rect 6850 -5062 7250 -5052
rect 6850 -5122 6860 -5062
rect 6920 -5122 7180 -5062
rect 7240 -5122 7250 -5062
rect 6850 -5232 7250 -5122
rect 7306 -5062 7706 -5052
rect 7306 -5122 7316 -5062
rect 7376 -5122 7636 -5062
rect 7696 -5122 7706 -5062
rect 7306 -5232 7706 -5122
rect 7762 -5062 8162 -5052
rect 7762 -5122 7772 -5062
rect 7832 -5122 8092 -5062
rect 8152 -5122 8162 -5062
rect 7762 -5232 8162 -5122
rect 8236 -5062 8636 -5052
rect 8236 -5122 8246 -5062
rect 8306 -5122 8566 -5062
rect 8626 -5122 8636 -5062
rect 8236 -5232 8636 -5122
rect 8692 -5062 9092 -5052
rect 8692 -5122 8702 -5062
rect 8762 -5122 9022 -5062
rect 9082 -5122 9092 -5062
rect 8692 -5232 9092 -5122
rect 9150 -5062 9550 -5052
rect 9150 -5122 9160 -5062
rect 9220 -5122 9480 -5062
rect 9540 -5122 9550 -5062
rect 9150 -5232 9550 -5122
rect 9606 -5062 10006 -5052
rect 9606 -5122 9616 -5062
rect 9676 -5122 9936 -5062
rect 9996 -5122 10006 -5062
rect 9606 -5232 10006 -5122
rect 10062 -5062 10462 -5052
rect 10062 -5122 10072 -5062
rect 10132 -5122 10392 -5062
rect 10452 -5122 10462 -5062
rect 10062 -5232 10462 -5122
rect 2740 -5233 10462 -5232
rect 10520 -5062 10920 -5052
rect 10520 -5122 10530 -5062
rect 10590 -5122 10850 -5062
rect 10910 -5122 10920 -5062
rect 10520 -5232 10920 -5122
rect 10976 -5062 11376 -5052
rect 10976 -5122 10986 -5062
rect 11046 -5122 11306 -5062
rect 11366 -5122 11376 -5062
rect 10976 -5232 11376 -5122
rect 11432 -5062 11832 -5052
rect 11432 -5122 11442 -5062
rect 11502 -5122 11762 -5062
rect 11822 -5122 11832 -5062
rect 11432 -5232 11832 -5122
rect 11890 -5062 12290 -5052
rect 11890 -5122 11900 -5062
rect 11960 -5122 12220 -5062
rect 12280 -5122 12290 -5062
rect 11890 -5232 12290 -5122
rect 12346 -5062 12746 -5052
rect 12346 -5122 12356 -5062
rect 12416 -5122 12676 -5062
rect 12736 -5122 12746 -5062
rect 12346 -5232 12746 -5122
rect 12802 -5062 13202 -5052
rect 12802 -5122 12812 -5062
rect 12872 -5122 13132 -5062
rect 13192 -5122 13202 -5062
rect 12802 -5232 13202 -5122
rect 13260 -5062 13660 -5052
rect 13260 -5122 13270 -5062
rect 13330 -5122 13590 -5062
rect 13650 -5122 13660 -5062
rect 13260 -5232 13660 -5122
rect 13716 -5062 14116 -5052
rect 13716 -5122 13726 -5062
rect 13786 -5122 14046 -5062
rect 14106 -5122 14116 -5062
rect 13716 -5232 14116 -5122
rect 14172 -5062 14572 -5052
rect 14172 -5122 14182 -5062
rect 14242 -5122 14502 -5062
rect 14562 -5122 14572 -5062
rect 14172 -5232 14572 -5122
rect 14630 -5062 15030 -5052
rect 14630 -5122 14640 -5062
rect 14700 -5122 14960 -5062
rect 15020 -5122 15030 -5062
rect 14630 -5232 15030 -5122
rect 15086 -5062 15486 -5052
rect 15086 -5122 15096 -5062
rect 15156 -5122 15416 -5062
rect 15476 -5122 15486 -5062
rect 15086 -5232 15486 -5122
rect 10520 -5233 15486 -5232
rect 456 -5303 15486 -5233
rect 456 -5412 856 -5303
rect 456 -5472 466 -5412
rect 526 -5472 786 -5412
rect 846 -5472 856 -5412
rect 456 -5482 856 -5472
rect 912 -5412 1312 -5303
rect 912 -5472 922 -5412
rect 982 -5472 1242 -5412
rect 1302 -5472 1312 -5412
rect 912 -5482 1312 -5472
rect 1370 -5412 1770 -5303
rect 1370 -5472 1380 -5412
rect 1440 -5472 1700 -5412
rect 1760 -5472 1770 -5412
rect 1370 -5482 1770 -5472
rect 1826 -5412 2226 -5303
rect 1826 -5472 1836 -5412
rect 1896 -5472 2156 -5412
rect 2216 -5472 2226 -5412
rect 1826 -5482 2226 -5472
rect 2282 -5412 2682 -5303
rect 2282 -5472 2292 -5412
rect 2352 -5472 2612 -5412
rect 2672 -5472 2682 -5412
rect 2282 -5482 2682 -5472
rect 2740 -5412 3140 -5303
rect 2740 -5472 2750 -5412
rect 2810 -5472 3070 -5412
rect 3130 -5472 3140 -5412
rect 2740 -5482 3140 -5472
rect 3196 -5412 3596 -5303
rect 3196 -5472 3206 -5412
rect 3266 -5472 3526 -5412
rect 3586 -5472 3596 -5412
rect 3196 -5482 3596 -5472
rect 3652 -5412 4052 -5303
rect 3652 -5472 3662 -5412
rect 3722 -5472 3982 -5412
rect 4042 -5472 4052 -5412
rect 3652 -5482 4052 -5472
rect 4110 -5412 4510 -5303
rect 4110 -5472 4120 -5412
rect 4180 -5472 4440 -5412
rect 4500 -5472 4510 -5412
rect 4110 -5482 4510 -5472
rect 4566 -5412 4966 -5303
rect 4566 -5472 4576 -5412
rect 4636 -5472 4896 -5412
rect 4956 -5472 4966 -5412
rect 4566 -5482 4966 -5472
rect 5022 -5412 5422 -5303
rect 5022 -5472 5032 -5412
rect 5092 -5472 5352 -5412
rect 5412 -5472 5422 -5412
rect 5022 -5482 5422 -5472
rect 5480 -5412 5880 -5303
rect 5480 -5472 5490 -5412
rect 5550 -5472 5810 -5412
rect 5870 -5472 5880 -5412
rect 5480 -5482 5880 -5472
rect 5936 -5412 6336 -5303
rect 5936 -5472 5946 -5412
rect 6006 -5472 6266 -5412
rect 6326 -5472 6336 -5412
rect 5936 -5482 6336 -5472
rect 6392 -5412 6792 -5303
rect 6392 -5472 6402 -5412
rect 6462 -5472 6722 -5412
rect 6782 -5472 6792 -5412
rect 6392 -5482 6792 -5472
rect 6850 -5412 7250 -5303
rect 6850 -5472 6860 -5412
rect 6920 -5472 7180 -5412
rect 7240 -5472 7250 -5412
rect 6850 -5482 7250 -5472
rect 7306 -5412 7706 -5303
rect 7306 -5472 7316 -5412
rect 7376 -5472 7636 -5412
rect 7696 -5472 7706 -5412
rect 7306 -5482 7706 -5472
rect 7762 -5412 8162 -5303
rect 7762 -5472 7772 -5412
rect 7832 -5472 8092 -5412
rect 8152 -5472 8162 -5412
rect 7762 -5482 8162 -5472
rect 8236 -5412 8636 -5303
rect 8236 -5472 8246 -5412
rect 8306 -5472 8566 -5412
rect 8626 -5472 8636 -5412
rect 8236 -5482 8636 -5472
rect 8692 -5412 9092 -5303
rect 8692 -5472 8702 -5412
rect 8762 -5472 9022 -5412
rect 9082 -5472 9092 -5412
rect 8692 -5482 9092 -5472
rect 9150 -5412 9550 -5303
rect 9150 -5472 9160 -5412
rect 9220 -5472 9480 -5412
rect 9540 -5472 9550 -5412
rect 9150 -5482 9550 -5472
rect 9606 -5412 10006 -5303
rect 9606 -5472 9616 -5412
rect 9676 -5472 9936 -5412
rect 9996 -5472 10006 -5412
rect 9606 -5482 10006 -5472
rect 10062 -5412 10462 -5303
rect 10062 -5472 10072 -5412
rect 10132 -5472 10392 -5412
rect 10452 -5472 10462 -5412
rect 10062 -5482 10462 -5472
rect 10520 -5412 10920 -5303
rect 10520 -5472 10530 -5412
rect 10590 -5472 10850 -5412
rect 10910 -5472 10920 -5412
rect 10520 -5482 10920 -5472
rect 10976 -5412 11376 -5303
rect 10976 -5472 10986 -5412
rect 11046 -5472 11306 -5412
rect 11366 -5472 11376 -5412
rect 10976 -5482 11376 -5472
rect 11432 -5412 11832 -5303
rect 11432 -5472 11442 -5412
rect 11502 -5472 11762 -5412
rect 11822 -5472 11832 -5412
rect 11432 -5482 11832 -5472
rect 11890 -5412 12290 -5303
rect 11890 -5472 11900 -5412
rect 11960 -5472 12220 -5412
rect 12280 -5472 12290 -5412
rect 11890 -5482 12290 -5472
rect 12346 -5412 12746 -5303
rect 12346 -5472 12356 -5412
rect 12416 -5472 12676 -5412
rect 12736 -5472 12746 -5412
rect 12346 -5482 12746 -5472
rect 12802 -5412 13202 -5303
rect 12802 -5472 12812 -5412
rect 12872 -5472 13132 -5412
rect 13192 -5472 13202 -5412
rect 12802 -5482 13202 -5472
rect 13260 -5412 13660 -5303
rect 13260 -5472 13270 -5412
rect 13330 -5472 13590 -5412
rect 13650 -5472 13660 -5412
rect 13260 -5482 13660 -5472
rect 13716 -5412 14116 -5303
rect 13716 -5472 13726 -5412
rect 13786 -5472 14046 -5412
rect 14106 -5472 14116 -5412
rect 13716 -5482 14116 -5472
rect 14172 -5412 14572 -5303
rect 14172 -5472 14182 -5412
rect 14242 -5472 14502 -5412
rect 14562 -5472 14572 -5412
rect 14172 -5482 14572 -5472
rect 14630 -5412 15030 -5303
rect 14630 -5472 14640 -5412
rect 14700 -5472 14960 -5412
rect 15020 -5472 15030 -5412
rect 14630 -5482 15030 -5472
rect 15086 -5412 15486 -5303
rect 15086 -5472 15096 -5412
rect 15156 -5472 15416 -5412
rect 15476 -5472 15486 -5412
rect 15086 -5482 15486 -5472
rect 66 -5544 80 -5482
rect 456 -5544 527 -5482
rect 912 -5544 983 -5482
rect 1370 -5544 1441 -5482
rect 1826 -5544 1897 -5482
rect 2282 -5544 2353 -5482
rect 2740 -5544 2810 -5482
rect 3196 -5544 3266 -5482
rect 3652 -5544 3722 -5482
rect 66 -5554 400 -5544
rect 0 -5614 10 -5554
rect 70 -5614 330 -5554
rect 390 -5614 400 -5554
rect 0 -5904 14 -5614
rect 66 -5904 400 -5614
rect 0 -5964 10 -5904
rect 70 -5964 330 -5904
rect 390 -5964 400 -5904
rect 0 -6051 14 -5964
rect 66 -5974 400 -5964
rect 456 -5554 856 -5544
rect 456 -5614 466 -5554
rect 526 -5614 786 -5554
rect 846 -5614 856 -5554
rect 456 -5724 856 -5614
rect 912 -5554 1312 -5544
rect 912 -5614 922 -5554
rect 982 -5614 1242 -5554
rect 1302 -5614 1312 -5554
rect 912 -5724 1312 -5614
rect 1370 -5554 1770 -5544
rect 1370 -5614 1380 -5554
rect 1440 -5614 1700 -5554
rect 1760 -5614 1770 -5554
rect 1370 -5724 1770 -5614
rect 1826 -5554 2226 -5544
rect 1826 -5614 1836 -5554
rect 1896 -5614 2156 -5554
rect 2216 -5614 2226 -5554
rect 1826 -5724 2226 -5614
rect 2282 -5554 2682 -5544
rect 2282 -5614 2292 -5554
rect 2352 -5614 2612 -5554
rect 2672 -5614 2682 -5554
rect 2282 -5724 2682 -5614
rect 456 -5725 2682 -5724
rect 2740 -5554 3140 -5544
rect 2740 -5614 2750 -5554
rect 2810 -5614 3070 -5554
rect 3130 -5614 3140 -5554
rect 2740 -5724 3140 -5614
rect 3196 -5554 3596 -5544
rect 3196 -5614 3206 -5554
rect 3266 -5614 3526 -5554
rect 3586 -5614 3596 -5554
rect 3196 -5724 3596 -5614
rect 3652 -5554 4052 -5544
rect 3652 -5614 3662 -5554
rect 3722 -5614 3982 -5554
rect 4042 -5614 4052 -5554
rect 3652 -5724 4052 -5614
rect 4110 -5554 4510 -5544
rect 4110 -5614 4120 -5554
rect 4180 -5614 4440 -5554
rect 4500 -5614 4510 -5554
rect 4110 -5724 4510 -5614
rect 4566 -5554 4966 -5544
rect 4566 -5614 4576 -5554
rect 4636 -5614 4896 -5554
rect 4956 -5614 4966 -5554
rect 4566 -5724 4966 -5614
rect 5022 -5554 5422 -5544
rect 5022 -5614 5032 -5554
rect 5092 -5614 5352 -5554
rect 5412 -5614 5422 -5554
rect 5022 -5724 5422 -5614
rect 5480 -5554 5880 -5544
rect 5480 -5614 5490 -5554
rect 5550 -5614 5810 -5554
rect 5870 -5614 5880 -5554
rect 5480 -5724 5880 -5614
rect 5936 -5554 6336 -5544
rect 5936 -5614 5946 -5554
rect 6006 -5614 6266 -5554
rect 6326 -5614 6336 -5554
rect 5936 -5724 6336 -5614
rect 6392 -5554 6792 -5544
rect 6392 -5614 6402 -5554
rect 6462 -5614 6722 -5554
rect 6782 -5614 6792 -5554
rect 6392 -5724 6792 -5614
rect 6850 -5554 7250 -5544
rect 6850 -5614 6860 -5554
rect 6920 -5614 7180 -5554
rect 7240 -5614 7250 -5554
rect 6850 -5724 7250 -5614
rect 7306 -5554 7706 -5544
rect 7306 -5614 7316 -5554
rect 7376 -5614 7636 -5554
rect 7696 -5614 7706 -5554
rect 7306 -5724 7706 -5614
rect 7762 -5554 8162 -5544
rect 7762 -5614 7772 -5554
rect 7832 -5614 8092 -5554
rect 8152 -5614 8162 -5554
rect 7762 -5724 8162 -5614
rect 8236 -5554 8636 -5544
rect 8236 -5614 8246 -5554
rect 8306 -5614 8566 -5554
rect 8626 -5614 8636 -5554
rect 8236 -5724 8636 -5614
rect 8692 -5554 9092 -5544
rect 8692 -5614 8702 -5554
rect 8762 -5614 9022 -5554
rect 9082 -5614 9092 -5554
rect 8692 -5724 9092 -5614
rect 9150 -5554 9550 -5544
rect 9150 -5614 9160 -5554
rect 9220 -5614 9480 -5554
rect 9540 -5614 9550 -5554
rect 9150 -5724 9550 -5614
rect 9606 -5554 10006 -5544
rect 9606 -5614 9616 -5554
rect 9676 -5614 9936 -5554
rect 9996 -5614 10006 -5554
rect 9606 -5724 10006 -5614
rect 10062 -5554 10462 -5544
rect 10062 -5614 10072 -5554
rect 10132 -5614 10392 -5554
rect 10452 -5614 10462 -5554
rect 10062 -5724 10462 -5614
rect 2740 -5725 4053 -5724
rect 456 -5795 4053 -5725
rect 4110 -5725 10462 -5724
rect 10520 -5554 10920 -5544
rect 10520 -5614 10530 -5554
rect 10590 -5614 10850 -5554
rect 10910 -5614 10920 -5554
rect 10520 -5724 10920 -5614
rect 10976 -5554 11376 -5544
rect 10976 -5614 10986 -5554
rect 11046 -5614 11306 -5554
rect 11366 -5614 11376 -5554
rect 10976 -5724 11376 -5614
rect 11432 -5554 11832 -5544
rect 11432 -5614 11442 -5554
rect 11502 -5614 11762 -5554
rect 11822 -5614 11832 -5554
rect 11432 -5724 11832 -5614
rect 11890 -5554 12290 -5544
rect 11890 -5614 11900 -5554
rect 11960 -5614 12220 -5554
rect 12280 -5614 12290 -5554
rect 11890 -5724 12290 -5614
rect 12346 -5554 12746 -5544
rect 12346 -5614 12356 -5554
rect 12416 -5614 12676 -5554
rect 12736 -5614 12746 -5554
rect 12346 -5724 12746 -5614
rect 12802 -5554 13202 -5544
rect 12802 -5614 12812 -5554
rect 12872 -5614 13132 -5554
rect 13192 -5614 13202 -5554
rect 12802 -5724 13202 -5614
rect 13260 -5554 13660 -5544
rect 13260 -5614 13270 -5554
rect 13330 -5614 13590 -5554
rect 13650 -5614 13660 -5554
rect 13260 -5724 13660 -5614
rect 13716 -5554 14116 -5544
rect 13716 -5614 13726 -5554
rect 13786 -5614 14046 -5554
rect 14106 -5614 14116 -5554
rect 13716 -5724 14116 -5614
rect 14172 -5554 14572 -5544
rect 14172 -5614 14182 -5554
rect 14242 -5614 14502 -5554
rect 14562 -5614 14572 -5554
rect 14172 -5724 14572 -5614
rect 14630 -5554 15030 -5544
rect 14630 -5614 14640 -5554
rect 14700 -5614 14960 -5554
rect 15020 -5614 15030 -5554
rect 14630 -5724 15030 -5614
rect 15086 -5554 15486 -5544
rect 15086 -5614 15096 -5554
rect 15156 -5614 15416 -5554
rect 15476 -5614 15486 -5554
rect 15086 -5724 15486 -5614
rect 10520 -5725 15486 -5724
rect 4110 -5795 15486 -5725
rect 456 -5904 856 -5795
rect 456 -5964 466 -5904
rect 526 -5964 786 -5904
rect 846 -5964 856 -5904
rect 456 -5974 856 -5964
rect 912 -5904 1312 -5795
rect 912 -5964 922 -5904
rect 982 -5964 1242 -5904
rect 1302 -5964 1312 -5904
rect 912 -5974 1312 -5964
rect 1370 -5904 1770 -5795
rect 1370 -5964 1380 -5904
rect 1440 -5964 1700 -5904
rect 1760 -5964 1770 -5904
rect 1370 -5974 1770 -5964
rect 1826 -5904 2226 -5795
rect 1826 -5964 1836 -5904
rect 1896 -5964 2156 -5904
rect 2216 -5964 2226 -5904
rect 1826 -5974 2226 -5964
rect 2282 -5904 2682 -5795
rect 2282 -5964 2292 -5904
rect 2352 -5964 2612 -5904
rect 2672 -5964 2682 -5904
rect 2282 -5974 2682 -5964
rect 2740 -5904 3140 -5795
rect 2740 -5964 2750 -5904
rect 2810 -5964 3070 -5904
rect 3130 -5964 3140 -5904
rect 2740 -5974 3140 -5964
rect 3196 -5904 3596 -5795
rect 3196 -5964 3206 -5904
rect 3266 -5964 3526 -5904
rect 3586 -5964 3596 -5904
rect 3196 -5974 3596 -5964
rect 3652 -5904 4052 -5795
rect 3652 -5964 3662 -5904
rect 3722 -5964 3982 -5904
rect 4042 -5964 4052 -5904
rect 3652 -5974 4052 -5964
rect 4110 -5904 4510 -5795
rect 4110 -5964 4120 -5904
rect 4180 -5964 4440 -5904
rect 4500 -5964 4510 -5904
rect 4110 -5974 4510 -5964
rect 4566 -5904 4966 -5795
rect 4566 -5964 4576 -5904
rect 4636 -5964 4896 -5904
rect 4956 -5964 4966 -5904
rect 4566 -5974 4966 -5964
rect 5022 -5904 5422 -5795
rect 5022 -5964 5032 -5904
rect 5092 -5964 5352 -5904
rect 5412 -5964 5422 -5904
rect 5022 -5974 5422 -5964
rect 5480 -5904 5880 -5795
rect 5480 -5964 5490 -5904
rect 5550 -5964 5810 -5904
rect 5870 -5964 5880 -5904
rect 5480 -5974 5880 -5964
rect 5936 -5904 6336 -5795
rect 5936 -5964 5946 -5904
rect 6006 -5964 6266 -5904
rect 6326 -5964 6336 -5904
rect 5936 -5974 6336 -5964
rect 6392 -5904 6792 -5795
rect 6392 -5964 6402 -5904
rect 6462 -5964 6722 -5904
rect 6782 -5964 6792 -5904
rect 6392 -5974 6792 -5964
rect 6850 -5904 7250 -5795
rect 6850 -5964 6860 -5904
rect 6920 -5964 7180 -5904
rect 7240 -5964 7250 -5904
rect 6850 -5974 7250 -5964
rect 7306 -5904 7706 -5795
rect 7306 -5964 7316 -5904
rect 7376 -5964 7636 -5904
rect 7696 -5964 7706 -5904
rect 7306 -5974 7706 -5964
rect 7762 -5904 8162 -5795
rect 7762 -5964 7772 -5904
rect 7832 -5964 8092 -5904
rect 8152 -5964 8162 -5904
rect 7762 -5974 8162 -5964
rect 8236 -5904 8636 -5795
rect 8236 -5964 8246 -5904
rect 8306 -5964 8566 -5904
rect 8626 -5964 8636 -5904
rect 8236 -5974 8636 -5964
rect 8692 -5904 9092 -5795
rect 8692 -5964 8702 -5904
rect 8762 -5964 9022 -5904
rect 9082 -5964 9092 -5904
rect 8692 -5974 9092 -5964
rect 9150 -5904 9550 -5795
rect 9150 -5964 9160 -5904
rect 9220 -5964 9480 -5904
rect 9540 -5964 9550 -5904
rect 9150 -5974 9550 -5964
rect 9606 -5904 10006 -5795
rect 9606 -5964 9616 -5904
rect 9676 -5964 9936 -5904
rect 9996 -5964 10006 -5904
rect 9606 -5974 10006 -5964
rect 10062 -5904 10462 -5795
rect 10062 -5964 10072 -5904
rect 10132 -5964 10392 -5904
rect 10452 -5964 10462 -5904
rect 10062 -5974 10462 -5964
rect 10520 -5904 10920 -5795
rect 10520 -5964 10530 -5904
rect 10590 -5964 10850 -5904
rect 10910 -5964 10920 -5904
rect 10520 -5974 10920 -5964
rect 10976 -5904 11376 -5795
rect 10976 -5964 10986 -5904
rect 11046 -5964 11306 -5904
rect 11366 -5964 11376 -5904
rect 10976 -5974 11376 -5964
rect 11432 -5904 11832 -5795
rect 11432 -5964 11442 -5904
rect 11502 -5964 11762 -5904
rect 11822 -5964 11832 -5904
rect 11432 -5974 11832 -5964
rect 11890 -5904 12290 -5795
rect 11890 -5964 11900 -5904
rect 11960 -5964 12220 -5904
rect 12280 -5964 12290 -5904
rect 11890 -5974 12290 -5964
rect 12346 -5904 12746 -5795
rect 12346 -5964 12356 -5904
rect 12416 -5964 12676 -5904
rect 12736 -5964 12746 -5904
rect 12346 -5974 12746 -5964
rect 12802 -5904 13202 -5795
rect 12802 -5964 12812 -5904
rect 12872 -5964 13132 -5904
rect 13192 -5964 13202 -5904
rect 12802 -5974 13202 -5964
rect 13260 -5904 13660 -5795
rect 13260 -5964 13270 -5904
rect 13330 -5964 13590 -5904
rect 13650 -5964 13660 -5904
rect 13260 -5974 13660 -5964
rect 13716 -5904 14116 -5795
rect 13716 -5964 13726 -5904
rect 13786 -5964 14046 -5904
rect 14106 -5964 14116 -5904
rect 13716 -5974 14116 -5964
rect 14172 -5904 14572 -5795
rect 14172 -5964 14182 -5904
rect 14242 -5964 14502 -5904
rect 14562 -5964 14572 -5904
rect 14172 -5974 14572 -5964
rect 14630 -5904 15030 -5795
rect 14630 -5964 14640 -5904
rect 14700 -5964 14960 -5904
rect 15020 -5964 15030 -5904
rect 14630 -5974 15030 -5964
rect 15086 -5904 15486 -5795
rect 15086 -5964 15096 -5904
rect 15156 -5964 15416 -5904
rect 15476 -5964 15486 -5904
rect 15086 -5974 15486 -5964
rect 66 -6041 80 -5974
rect 456 -5975 527 -5974
rect 457 -6041 527 -5975
rect 913 -6041 984 -5974
rect 1371 -6041 1442 -5974
rect 1827 -6041 1898 -5974
rect 2283 -6041 2354 -5974
rect 2741 -6041 2812 -5974
rect 3197 -6041 3268 -5974
rect 3653 -6041 3724 -5974
rect 4111 -6041 4182 -5974
rect 4567 -6041 4638 -5974
rect 5023 -6041 5094 -5974
rect 5481 -6041 5552 -5974
rect 5937 -6041 6008 -5974
rect 6393 -6041 6464 -5974
rect 6851 -6041 6922 -5974
rect 7307 -6041 7378 -5974
rect 7763 -6041 7834 -5974
rect 8237 -6041 8308 -5974
rect 8693 -6041 8764 -5974
rect 9151 -6041 9222 -5974
rect 9607 -6041 9678 -5974
rect 10063 -6041 10134 -5974
rect 10521 -6041 10592 -5974
rect 10977 -6041 11048 -5974
rect 11433 -6041 11504 -5974
rect 11891 -6041 11962 -5974
rect 12347 -6041 12418 -5974
rect 12803 -6041 12874 -5974
rect 13261 -6041 13332 -5974
rect 13717 -6041 13788 -5974
rect 14173 -6041 14244 -5974
rect 14631 -6041 14702 -5974
rect 66 -6051 400 -6041
rect 0 -6111 11 -6051
rect 71 -6111 331 -6051
rect 391 -6111 400 -6051
rect 0 -6401 14 -6111
rect 66 -6401 400 -6111
rect 0 -6461 11 -6401
rect 71 -6461 331 -6401
rect 391 -6461 400 -6401
rect 0 -6543 14 -6461
rect 66 -6471 400 -6461
rect 457 -6051 857 -6041
rect 457 -6111 467 -6051
rect 527 -6111 787 -6051
rect 847 -6111 857 -6051
rect 457 -6219 857 -6111
rect 913 -6051 1313 -6041
rect 913 -6111 923 -6051
rect 983 -6111 1243 -6051
rect 1303 -6111 1313 -6051
rect 913 -6219 1313 -6111
rect 1371 -6051 1771 -6041
rect 1371 -6111 1381 -6051
rect 1441 -6111 1701 -6051
rect 1761 -6111 1771 -6051
rect 1371 -6219 1771 -6111
rect 1827 -6051 2227 -6041
rect 1827 -6111 1837 -6051
rect 1897 -6111 2157 -6051
rect 2217 -6111 2227 -6051
rect 1827 -6219 2227 -6111
rect 2283 -6051 2683 -6041
rect 2283 -6111 2293 -6051
rect 2353 -6111 2613 -6051
rect 2673 -6111 2683 -6051
rect 2283 -6219 2683 -6111
rect 2741 -6051 3141 -6041
rect 2741 -6111 2751 -6051
rect 2811 -6111 3071 -6051
rect 3131 -6111 3141 -6051
rect 2741 -6219 3141 -6111
rect 3197 -6051 3597 -6041
rect 3197 -6111 3207 -6051
rect 3267 -6111 3527 -6051
rect 3587 -6111 3597 -6051
rect 3197 -6219 3597 -6111
rect 3653 -6051 4053 -6041
rect 3653 -6111 3663 -6051
rect 3723 -6111 3983 -6051
rect 4043 -6111 4053 -6051
rect 3653 -6219 4053 -6111
rect 4111 -6051 4511 -6041
rect 4111 -6111 4121 -6051
rect 4181 -6111 4441 -6051
rect 4501 -6111 4511 -6051
rect 4111 -6219 4511 -6111
rect 4567 -6051 4967 -6041
rect 4567 -6111 4577 -6051
rect 4637 -6111 4897 -6051
rect 4957 -6111 4967 -6051
rect 4567 -6219 4967 -6111
rect 5023 -6051 5423 -6041
rect 5023 -6111 5033 -6051
rect 5093 -6111 5353 -6051
rect 5413 -6111 5423 -6051
rect 5023 -6219 5423 -6111
rect 5481 -6051 5881 -6041
rect 5481 -6111 5491 -6051
rect 5551 -6111 5811 -6051
rect 5871 -6111 5881 -6051
rect 5481 -6219 5881 -6111
rect 5937 -6051 6337 -6041
rect 5937 -6111 5947 -6051
rect 6007 -6111 6267 -6051
rect 6327 -6111 6337 -6051
rect 5937 -6219 6337 -6111
rect 6393 -6051 6793 -6041
rect 6393 -6111 6403 -6051
rect 6463 -6111 6723 -6051
rect 6783 -6111 6793 -6051
rect 6393 -6219 6793 -6111
rect 6851 -6051 7251 -6041
rect 6851 -6111 6861 -6051
rect 6921 -6111 7181 -6051
rect 7241 -6111 7251 -6051
rect 6851 -6219 7251 -6111
rect 7307 -6051 7707 -6041
rect 7307 -6111 7317 -6051
rect 7377 -6111 7637 -6051
rect 7697 -6111 7707 -6051
rect 7307 -6219 7707 -6111
rect 7763 -6051 8163 -6041
rect 7763 -6111 7773 -6051
rect 7833 -6111 8093 -6051
rect 8153 -6111 8163 -6051
rect 7763 -6219 8163 -6111
rect 8237 -6051 8637 -6041
rect 8237 -6111 8247 -6051
rect 8307 -6111 8567 -6051
rect 8627 -6111 8637 -6051
rect 8237 -6219 8637 -6111
rect 8693 -6051 9093 -6041
rect 8693 -6111 8703 -6051
rect 8763 -6111 9023 -6051
rect 9083 -6111 9093 -6051
rect 8693 -6219 9093 -6111
rect 9151 -6051 9551 -6041
rect 9151 -6111 9161 -6051
rect 9221 -6111 9481 -6051
rect 9541 -6111 9551 -6051
rect 9151 -6219 9551 -6111
rect 9607 -6051 10007 -6041
rect 9607 -6111 9617 -6051
rect 9677 -6111 9937 -6051
rect 9997 -6111 10007 -6051
rect 9607 -6219 10007 -6111
rect 10063 -6051 10463 -6041
rect 10063 -6111 10073 -6051
rect 10133 -6111 10393 -6051
rect 10453 -6111 10463 -6051
rect 10063 -6219 10463 -6111
rect 10521 -6051 10921 -6041
rect 10521 -6111 10531 -6051
rect 10591 -6111 10851 -6051
rect 10911 -6111 10921 -6051
rect 10521 -6219 10921 -6111
rect 10977 -6051 11377 -6041
rect 10977 -6111 10987 -6051
rect 11047 -6111 11307 -6051
rect 11367 -6111 11377 -6051
rect 10977 -6219 11377 -6111
rect 11433 -6051 11833 -6041
rect 11433 -6111 11443 -6051
rect 11503 -6111 11763 -6051
rect 11823 -6111 11833 -6051
rect 11433 -6219 11833 -6111
rect 11891 -6051 12291 -6041
rect 11891 -6111 11901 -6051
rect 11961 -6111 12221 -6051
rect 12281 -6111 12291 -6051
rect 11891 -6219 12291 -6111
rect 12347 -6051 12747 -6041
rect 12347 -6111 12357 -6051
rect 12417 -6111 12677 -6051
rect 12737 -6111 12747 -6051
rect 12347 -6219 12747 -6111
rect 12803 -6051 13203 -6041
rect 12803 -6111 12813 -6051
rect 12873 -6111 13133 -6051
rect 13193 -6111 13203 -6051
rect 12803 -6219 13203 -6111
rect 13261 -6051 13661 -6041
rect 13261 -6111 13271 -6051
rect 13331 -6111 13591 -6051
rect 13651 -6111 13661 -6051
rect 13261 -6219 13661 -6111
rect 13717 -6051 14117 -6041
rect 13717 -6111 13727 -6051
rect 13787 -6111 14047 -6051
rect 14107 -6111 14117 -6051
rect 13717 -6219 14117 -6111
rect 14173 -6051 14573 -6041
rect 14173 -6111 14183 -6051
rect 14243 -6111 14503 -6051
rect 14563 -6111 14573 -6051
rect 14173 -6219 14573 -6111
rect 14631 -6051 15031 -6041
rect 14631 -6111 14641 -6051
rect 14701 -6111 14961 -6051
rect 15021 -6111 15031 -6051
rect 14631 -6219 15031 -6111
rect 15087 -6051 15487 -6041
rect 15087 -6111 15097 -6051
rect 15157 -6111 15417 -6051
rect 15477 -6111 15487 -6051
rect 15087 -6219 15487 -6111
rect 457 -6289 4053 -6219
rect 457 -6291 2683 -6289
rect 457 -6401 857 -6291
rect 457 -6461 467 -6401
rect 527 -6461 787 -6401
rect 847 -6461 857 -6401
rect 457 -6471 857 -6461
rect 913 -6401 1313 -6291
rect 913 -6461 923 -6401
rect 983 -6461 1243 -6401
rect 1303 -6461 1313 -6401
rect 913 -6471 1313 -6461
rect 1371 -6401 1771 -6291
rect 1371 -6461 1381 -6401
rect 1441 -6461 1701 -6401
rect 1761 -6461 1771 -6401
rect 1371 -6471 1771 -6461
rect 1827 -6401 2227 -6291
rect 1827 -6461 1837 -6401
rect 1897 -6461 2157 -6401
rect 2217 -6461 2227 -6401
rect 1827 -6471 2227 -6461
rect 2283 -6401 2683 -6291
rect 2283 -6461 2293 -6401
rect 2353 -6461 2613 -6401
rect 2673 -6461 2683 -6401
rect 2283 -6471 2683 -6461
rect 2741 -6291 4053 -6289
rect 4110 -6289 15487 -6219
rect 4110 -6291 10463 -6289
rect 2741 -6401 3141 -6291
rect 2741 -6461 2751 -6401
rect 2811 -6461 3071 -6401
rect 3131 -6461 3141 -6401
rect 2741 -6471 3141 -6461
rect 3197 -6401 3597 -6291
rect 3197 -6461 3207 -6401
rect 3267 -6461 3527 -6401
rect 3587 -6461 3597 -6401
rect 3197 -6471 3597 -6461
rect 3653 -6401 4053 -6291
rect 3653 -6461 3663 -6401
rect 3723 -6461 3983 -6401
rect 4043 -6461 4053 -6401
rect 3653 -6471 4053 -6461
rect 4111 -6401 4511 -6291
rect 4111 -6461 4121 -6401
rect 4181 -6461 4441 -6401
rect 4501 -6461 4511 -6401
rect 4111 -6471 4511 -6461
rect 4567 -6401 4967 -6291
rect 4567 -6461 4577 -6401
rect 4637 -6461 4897 -6401
rect 4957 -6461 4967 -6401
rect 4567 -6471 4967 -6461
rect 5023 -6401 5423 -6291
rect 5023 -6461 5033 -6401
rect 5093 -6461 5353 -6401
rect 5413 -6461 5423 -6401
rect 5023 -6471 5423 -6461
rect 5481 -6401 5881 -6291
rect 5481 -6461 5491 -6401
rect 5551 -6461 5811 -6401
rect 5871 -6461 5881 -6401
rect 5481 -6471 5881 -6461
rect 5937 -6401 6337 -6291
rect 5937 -6461 5947 -6401
rect 6007 -6461 6267 -6401
rect 6327 -6461 6337 -6401
rect 5937 -6471 6337 -6461
rect 6393 -6401 6793 -6291
rect 6393 -6461 6403 -6401
rect 6463 -6461 6723 -6401
rect 6783 -6461 6793 -6401
rect 6393 -6471 6793 -6461
rect 6851 -6401 7251 -6291
rect 6851 -6461 6861 -6401
rect 6921 -6461 7181 -6401
rect 7241 -6461 7251 -6401
rect 6851 -6471 7251 -6461
rect 7307 -6401 7707 -6291
rect 7307 -6461 7317 -6401
rect 7377 -6461 7637 -6401
rect 7697 -6461 7707 -6401
rect 7307 -6471 7707 -6461
rect 7763 -6401 8163 -6291
rect 7763 -6461 7773 -6401
rect 7833 -6461 8093 -6401
rect 8153 -6461 8163 -6401
rect 7763 -6471 8163 -6461
rect 8237 -6401 8637 -6291
rect 8237 -6461 8247 -6401
rect 8307 -6461 8567 -6401
rect 8627 -6461 8637 -6401
rect 8237 -6471 8637 -6461
rect 8693 -6401 9093 -6291
rect 8693 -6461 8703 -6401
rect 8763 -6461 9023 -6401
rect 9083 -6461 9093 -6401
rect 8693 -6471 9093 -6461
rect 9151 -6401 9551 -6291
rect 9151 -6461 9161 -6401
rect 9221 -6461 9481 -6401
rect 9541 -6461 9551 -6401
rect 9151 -6471 9551 -6461
rect 9607 -6401 10007 -6291
rect 9607 -6461 9617 -6401
rect 9677 -6461 9937 -6401
rect 9997 -6461 10007 -6401
rect 9607 -6471 10007 -6461
rect 10063 -6401 10463 -6291
rect 10063 -6461 10073 -6401
rect 10133 -6461 10393 -6401
rect 10453 -6461 10463 -6401
rect 10063 -6471 10463 -6461
rect 10521 -6291 15487 -6289
rect 10521 -6401 10921 -6291
rect 10521 -6461 10531 -6401
rect 10591 -6461 10851 -6401
rect 10911 -6461 10921 -6401
rect 10521 -6471 10921 -6461
rect 10977 -6401 11377 -6291
rect 10977 -6461 10987 -6401
rect 11047 -6461 11307 -6401
rect 11367 -6461 11377 -6401
rect 10977 -6471 11377 -6461
rect 11433 -6401 11833 -6291
rect 11433 -6461 11443 -6401
rect 11503 -6461 11763 -6401
rect 11823 -6461 11833 -6401
rect 11433 -6471 11833 -6461
rect 11891 -6401 12291 -6291
rect 11891 -6461 11901 -6401
rect 11961 -6461 12221 -6401
rect 12281 -6461 12291 -6401
rect 11891 -6471 12291 -6461
rect 12347 -6401 12747 -6291
rect 12347 -6461 12357 -6401
rect 12417 -6461 12677 -6401
rect 12737 -6461 12747 -6401
rect 12347 -6471 12747 -6461
rect 12803 -6401 13203 -6291
rect 12803 -6461 12813 -6401
rect 12873 -6461 13133 -6401
rect 13193 -6461 13203 -6401
rect 12803 -6471 13203 -6461
rect 13261 -6401 13661 -6291
rect 13261 -6461 13271 -6401
rect 13331 -6461 13591 -6401
rect 13651 -6461 13661 -6401
rect 13261 -6471 13661 -6461
rect 13717 -6401 14117 -6291
rect 13717 -6461 13727 -6401
rect 13787 -6461 14047 -6401
rect 14107 -6461 14117 -6401
rect 13717 -6471 14117 -6461
rect 14173 -6401 14573 -6291
rect 14173 -6461 14183 -6401
rect 14243 -6461 14503 -6401
rect 14563 -6461 14573 -6401
rect 14173 -6471 14573 -6461
rect 14631 -6401 15031 -6291
rect 14631 -6461 14641 -6401
rect 14701 -6461 14961 -6401
rect 15021 -6461 15031 -6401
rect 14631 -6471 15031 -6461
rect 15087 -6401 15487 -6291
rect 15087 -6461 15097 -6401
rect 15157 -6461 15417 -6401
rect 15477 -6461 15487 -6401
rect 15087 -6471 15487 -6461
rect 66 -6533 80 -6471
rect 457 -6533 528 -6471
rect 913 -6533 984 -6471
rect 1371 -6533 1442 -6471
rect 1827 -6533 1898 -6471
rect 2283 -6533 2354 -6471
rect 2741 -6533 2811 -6471
rect 3197 -6533 3267 -6471
rect 3653 -6533 3723 -6471
rect 4111 -6533 4181 -6471
rect 4567 -6533 4637 -6471
rect 5023 -6533 5093 -6471
rect 5481 -6533 5551 -6471
rect 5937 -6533 6007 -6471
rect 6393 -6533 6463 -6471
rect 6851 -6533 6921 -6471
rect 7307 -6533 7377 -6471
rect 7763 -6533 7833 -6471
rect 8237 -6533 8307 -6471
rect 8693 -6533 8763 -6471
rect 9151 -6533 9221 -6471
rect 9607 -6533 9677 -6471
rect 10063 -6533 10133 -6471
rect 10521 -6533 10591 -6471
rect 10977 -6533 11047 -6471
rect 11433 -6533 11503 -6471
rect 11891 -6533 11961 -6471
rect 12347 -6533 12417 -6471
rect 12803 -6533 12873 -6471
rect 13261 -6533 13331 -6471
rect 13717 -6533 13787 -6471
rect 14173 -6533 14243 -6471
rect 14631 -6533 14701 -6471
rect 66 -6543 400 -6533
rect 0 -6603 11 -6543
rect 71 -6603 331 -6543
rect 391 -6603 400 -6543
rect 0 -6893 14 -6603
rect 66 -6893 400 -6603
rect 0 -6953 11 -6893
rect 71 -6953 331 -6893
rect 391 -6953 400 -6893
rect 0 -7059 14 -6953
rect 66 -6963 400 -6953
rect 457 -6543 857 -6533
rect 457 -6603 467 -6543
rect 527 -6603 787 -6543
rect 847 -6603 857 -6543
rect 457 -6712 857 -6603
rect 913 -6543 1313 -6533
rect 913 -6603 923 -6543
rect 983 -6603 1243 -6543
rect 1303 -6603 1313 -6543
rect 913 -6712 1313 -6603
rect 1371 -6543 1771 -6533
rect 1371 -6603 1381 -6543
rect 1441 -6603 1701 -6543
rect 1761 -6603 1771 -6543
rect 1371 -6712 1771 -6603
rect 1827 -6543 2227 -6533
rect 1827 -6603 1837 -6543
rect 1897 -6603 2157 -6543
rect 2217 -6603 2227 -6543
rect 1827 -6712 2227 -6603
rect 2283 -6543 2683 -6533
rect 2283 -6603 2293 -6543
rect 2353 -6603 2613 -6543
rect 2673 -6603 2683 -6543
rect 2283 -6712 2683 -6603
rect 2741 -6543 3141 -6533
rect 2741 -6603 2751 -6543
rect 2811 -6603 3071 -6543
rect 3131 -6603 3141 -6543
rect 2741 -6712 3141 -6603
rect 3197 -6543 3597 -6533
rect 3197 -6603 3207 -6543
rect 3267 -6603 3527 -6543
rect 3587 -6603 3597 -6543
rect 3197 -6712 3597 -6603
rect 3653 -6543 4053 -6533
rect 3653 -6603 3663 -6543
rect 3723 -6603 3983 -6543
rect 4043 -6603 4053 -6543
rect 3653 -6712 4053 -6603
rect 4111 -6543 4511 -6533
rect 4111 -6603 4121 -6543
rect 4181 -6603 4441 -6543
rect 4501 -6603 4511 -6543
rect 4111 -6712 4511 -6603
rect 4567 -6543 4967 -6533
rect 4567 -6603 4577 -6543
rect 4637 -6603 4897 -6543
rect 4957 -6603 4967 -6543
rect 4567 -6712 4967 -6603
rect 5023 -6543 5423 -6533
rect 5023 -6603 5033 -6543
rect 5093 -6603 5353 -6543
rect 5413 -6603 5423 -6543
rect 5023 -6712 5423 -6603
rect 5481 -6543 5881 -6533
rect 5481 -6603 5491 -6543
rect 5551 -6603 5811 -6543
rect 5871 -6603 5881 -6543
rect 5481 -6712 5881 -6603
rect 5937 -6543 6337 -6533
rect 5937 -6603 5947 -6543
rect 6007 -6603 6267 -6543
rect 6327 -6603 6337 -6543
rect 5937 -6712 6337 -6603
rect 6393 -6543 6793 -6533
rect 6393 -6603 6403 -6543
rect 6463 -6603 6723 -6543
rect 6783 -6603 6793 -6543
rect 6393 -6712 6793 -6603
rect 6851 -6543 7251 -6533
rect 6851 -6603 6861 -6543
rect 6921 -6603 7181 -6543
rect 7241 -6603 7251 -6543
rect 6851 -6712 7251 -6603
rect 7307 -6543 7707 -6533
rect 7307 -6603 7317 -6543
rect 7377 -6603 7637 -6543
rect 7697 -6603 7707 -6543
rect 7307 -6712 7707 -6603
rect 7763 -6543 8163 -6533
rect 7763 -6603 7773 -6543
rect 7833 -6603 8093 -6543
rect 8153 -6603 8163 -6543
rect 7763 -6712 8163 -6603
rect 8237 -6543 8637 -6533
rect 8237 -6603 8247 -6543
rect 8307 -6603 8567 -6543
rect 8627 -6603 8637 -6543
rect 8237 -6712 8637 -6603
rect 8693 -6543 9093 -6533
rect 8693 -6603 8703 -6543
rect 8763 -6603 9023 -6543
rect 9083 -6603 9093 -6543
rect 8693 -6712 9093 -6603
rect 9151 -6543 9551 -6533
rect 9151 -6603 9161 -6543
rect 9221 -6603 9481 -6543
rect 9541 -6603 9551 -6543
rect 9151 -6712 9551 -6603
rect 9607 -6543 10007 -6533
rect 9607 -6603 9617 -6543
rect 9677 -6603 9937 -6543
rect 9997 -6603 10007 -6543
rect 9607 -6712 10007 -6603
rect 10063 -6543 10463 -6533
rect 10063 -6603 10073 -6543
rect 10133 -6603 10393 -6543
rect 10453 -6603 10463 -6543
rect 10063 -6712 10463 -6603
rect 10521 -6543 10921 -6533
rect 10521 -6603 10531 -6543
rect 10591 -6603 10851 -6543
rect 10911 -6603 10921 -6543
rect 10521 -6712 10921 -6603
rect 10977 -6543 11377 -6533
rect 10977 -6603 10987 -6543
rect 11047 -6603 11307 -6543
rect 11367 -6603 11377 -6543
rect 10977 -6712 11377 -6603
rect 11433 -6543 11833 -6533
rect 11433 -6603 11443 -6543
rect 11503 -6603 11763 -6543
rect 11823 -6603 11833 -6543
rect 11433 -6712 11833 -6603
rect 11891 -6543 12291 -6533
rect 11891 -6603 11901 -6543
rect 11961 -6603 12221 -6543
rect 12281 -6603 12291 -6543
rect 11891 -6712 12291 -6603
rect 12347 -6543 12747 -6533
rect 12347 -6603 12357 -6543
rect 12417 -6603 12677 -6543
rect 12737 -6603 12747 -6543
rect 12347 -6712 12747 -6603
rect 12803 -6543 13203 -6533
rect 12803 -6603 12813 -6543
rect 12873 -6603 13133 -6543
rect 13193 -6603 13203 -6543
rect 12803 -6712 13203 -6603
rect 13261 -6543 13661 -6533
rect 13261 -6603 13271 -6543
rect 13331 -6603 13591 -6543
rect 13651 -6603 13661 -6543
rect 13261 -6712 13661 -6603
rect 13717 -6543 14117 -6533
rect 13717 -6603 13727 -6543
rect 13787 -6603 14047 -6543
rect 14107 -6603 14117 -6543
rect 13717 -6712 14117 -6603
rect 14173 -6543 14573 -6533
rect 14173 -6603 14183 -6543
rect 14243 -6603 14503 -6543
rect 14563 -6603 14573 -6543
rect 14173 -6712 14573 -6603
rect 14631 -6543 15031 -6533
rect 14631 -6603 14641 -6543
rect 14701 -6603 14961 -6543
rect 15021 -6603 15031 -6543
rect 14631 -6712 15031 -6603
rect 15087 -6543 15487 -6533
rect 15087 -6603 15097 -6543
rect 15157 -6603 15417 -6543
rect 15477 -6603 15487 -6543
rect 15087 -6712 15487 -6603
rect 457 -6782 4053 -6712
rect 457 -6783 2683 -6782
rect 457 -6893 857 -6783
rect 457 -6953 467 -6893
rect 527 -6953 787 -6893
rect 847 -6953 857 -6893
rect 457 -6963 857 -6953
rect 913 -6893 1313 -6783
rect 913 -6953 923 -6893
rect 983 -6953 1243 -6893
rect 1303 -6953 1313 -6893
rect 913 -6963 1313 -6953
rect 1371 -6893 1771 -6783
rect 1371 -6953 1381 -6893
rect 1441 -6953 1701 -6893
rect 1761 -6953 1771 -6893
rect 1371 -6963 1771 -6953
rect 1827 -6893 2227 -6783
rect 1827 -6953 1837 -6893
rect 1897 -6953 2157 -6893
rect 2217 -6953 2227 -6893
rect 1827 -6963 2227 -6953
rect 2283 -6893 2683 -6783
rect 2283 -6953 2293 -6893
rect 2353 -6953 2613 -6893
rect 2673 -6953 2683 -6893
rect 2283 -6963 2683 -6953
rect 2741 -6783 4053 -6782
rect 4110 -6782 15487 -6712
rect 4110 -6783 10463 -6782
rect 2741 -6893 3141 -6783
rect 2741 -6953 2751 -6893
rect 2811 -6953 3071 -6893
rect 3131 -6953 3141 -6893
rect 2741 -6963 3141 -6953
rect 3197 -6893 3597 -6783
rect 3197 -6953 3207 -6893
rect 3267 -6953 3527 -6893
rect 3587 -6953 3597 -6893
rect 3197 -6963 3597 -6953
rect 3653 -6893 4053 -6783
rect 3653 -6953 3663 -6893
rect 3723 -6953 3983 -6893
rect 4043 -6953 4053 -6893
rect 3653 -6963 4053 -6953
rect 4111 -6893 4511 -6783
rect 4111 -6953 4121 -6893
rect 4181 -6953 4441 -6893
rect 4501 -6953 4511 -6893
rect 4111 -6963 4511 -6953
rect 4567 -6893 4967 -6783
rect 4567 -6953 4577 -6893
rect 4637 -6953 4897 -6893
rect 4957 -6953 4967 -6893
rect 4567 -6963 4967 -6953
rect 5023 -6893 5423 -6783
rect 5023 -6953 5033 -6893
rect 5093 -6953 5353 -6893
rect 5413 -6953 5423 -6893
rect 5023 -6963 5423 -6953
rect 5481 -6893 5881 -6783
rect 5481 -6953 5491 -6893
rect 5551 -6953 5811 -6893
rect 5871 -6953 5881 -6893
rect 5481 -6963 5881 -6953
rect 5937 -6893 6337 -6783
rect 5937 -6953 5947 -6893
rect 6007 -6953 6267 -6893
rect 6327 -6953 6337 -6893
rect 5937 -6963 6337 -6953
rect 6393 -6893 6793 -6783
rect 6393 -6953 6403 -6893
rect 6463 -6953 6723 -6893
rect 6783 -6953 6793 -6893
rect 6393 -6963 6793 -6953
rect 6851 -6893 7251 -6783
rect 6851 -6953 6861 -6893
rect 6921 -6953 7181 -6893
rect 7241 -6953 7251 -6893
rect 6851 -6963 7251 -6953
rect 7307 -6893 7707 -6783
rect 7307 -6953 7317 -6893
rect 7377 -6953 7637 -6893
rect 7697 -6953 7707 -6893
rect 7307 -6963 7707 -6953
rect 7763 -6893 8163 -6783
rect 7763 -6953 7773 -6893
rect 7833 -6953 8093 -6893
rect 8153 -6953 8163 -6893
rect 7763 -6963 8163 -6953
rect 8237 -6893 8637 -6783
rect 8237 -6953 8247 -6893
rect 8307 -6953 8567 -6893
rect 8627 -6953 8637 -6893
rect 8237 -6963 8637 -6953
rect 8693 -6893 9093 -6783
rect 8693 -6953 8703 -6893
rect 8763 -6953 9023 -6893
rect 9083 -6953 9093 -6893
rect 8693 -6963 9093 -6953
rect 9151 -6893 9551 -6783
rect 9151 -6953 9161 -6893
rect 9221 -6953 9481 -6893
rect 9541 -6953 9551 -6893
rect 9151 -6963 9551 -6953
rect 9607 -6893 10007 -6783
rect 9607 -6953 9617 -6893
rect 9677 -6953 9937 -6893
rect 9997 -6953 10007 -6893
rect 9607 -6963 10007 -6953
rect 10063 -6893 10463 -6783
rect 10063 -6953 10073 -6893
rect 10133 -6953 10393 -6893
rect 10453 -6953 10463 -6893
rect 10063 -6963 10463 -6953
rect 10521 -6783 15487 -6782
rect 10521 -6893 10921 -6783
rect 10521 -6953 10531 -6893
rect 10591 -6953 10851 -6893
rect 10911 -6953 10921 -6893
rect 10521 -6963 10921 -6953
rect 10977 -6893 11377 -6783
rect 10977 -6953 10987 -6893
rect 11047 -6953 11307 -6893
rect 11367 -6953 11377 -6893
rect 10977 -6963 11377 -6953
rect 11433 -6893 11833 -6783
rect 11433 -6953 11443 -6893
rect 11503 -6953 11763 -6893
rect 11823 -6953 11833 -6893
rect 11433 -6963 11833 -6953
rect 11891 -6893 12291 -6783
rect 11891 -6953 11901 -6893
rect 11961 -6953 12221 -6893
rect 12281 -6953 12291 -6893
rect 11891 -6963 12291 -6953
rect 12347 -6893 12747 -6783
rect 12347 -6953 12357 -6893
rect 12417 -6953 12677 -6893
rect 12737 -6953 12747 -6893
rect 12347 -6963 12747 -6953
rect 12803 -6893 13203 -6783
rect 12803 -6953 12813 -6893
rect 12873 -6953 13133 -6893
rect 13193 -6953 13203 -6893
rect 12803 -6963 13203 -6953
rect 13261 -6893 13661 -6783
rect 13261 -6953 13271 -6893
rect 13331 -6953 13591 -6893
rect 13651 -6953 13661 -6893
rect 13261 -6963 13661 -6953
rect 13717 -6893 14117 -6783
rect 13717 -6953 13727 -6893
rect 13787 -6953 14047 -6893
rect 14107 -6953 14117 -6893
rect 13717 -6963 14117 -6953
rect 14173 -6893 14573 -6783
rect 14173 -6953 14183 -6893
rect 14243 -6953 14503 -6893
rect 14563 -6953 14573 -6893
rect 14173 -6963 14573 -6953
rect 14631 -6893 15031 -6783
rect 14631 -6953 14641 -6893
rect 14701 -6953 14961 -6893
rect 15021 -6953 15031 -6893
rect 14631 -6963 15031 -6953
rect 15087 -6893 15487 -6783
rect 15087 -6953 15097 -6893
rect 15157 -6953 15417 -6893
rect 15477 -6953 15487 -6893
rect 15087 -6963 15487 -6953
rect 66 -7049 80 -6963
rect 457 -7049 527 -6963
rect 913 -7049 983 -6963
rect 1371 -7049 1441 -6963
rect 1827 -7049 1897 -6963
rect 2283 -7049 2353 -6963
rect 2741 -7049 2811 -6963
rect 3197 -7049 3267 -6963
rect 3653 -7049 3723 -6963
rect 4111 -7049 4181 -6963
rect 4567 -7049 4637 -6963
rect 5023 -7049 5093 -6963
rect 5481 -7049 5551 -6963
rect 5937 -7049 6007 -6963
rect 6393 -7049 6463 -6963
rect 6851 -7049 6921 -6963
rect 7307 -7049 7377 -6963
rect 7763 -7049 7833 -6963
rect 8237 -7049 8307 -6963
rect 8693 -7049 8763 -6963
rect 9151 -7049 9221 -6963
rect 9607 -7049 9677 -6963
rect 10063 -7049 10133 -6963
rect 10521 -7049 10591 -6963
rect 10977 -7049 11047 -6963
rect 11433 -7049 11503 -6963
rect 11891 -7049 11961 -6963
rect 12347 -7049 12417 -6963
rect 12803 -7049 12873 -6963
rect 13261 -7049 13331 -6963
rect 13717 -7049 13787 -6963
rect 14173 -7049 14243 -6963
rect 14631 -7049 14701 -6963
rect 66 -7059 400 -7049
rect 0 -7119 11 -7059
rect 71 -7119 331 -7059
rect 391 -7119 400 -7059
rect 0 -7409 14 -7119
rect 66 -7409 400 -7119
rect 0 -7469 11 -7409
rect 71 -7469 331 -7409
rect 391 -7469 400 -7409
rect 0 -7561 14 -7469
rect 66 -7479 400 -7469
rect 457 -7059 857 -7049
rect 457 -7119 467 -7059
rect 527 -7119 787 -7059
rect 847 -7119 857 -7059
rect 457 -7229 857 -7119
rect 913 -7059 1313 -7049
rect 913 -7119 923 -7059
rect 983 -7119 1243 -7059
rect 1303 -7119 1313 -7059
rect 913 -7229 1313 -7119
rect 1371 -7059 1771 -7049
rect 1371 -7119 1381 -7059
rect 1441 -7119 1701 -7059
rect 1761 -7119 1771 -7059
rect 1371 -7229 1771 -7119
rect 1827 -7059 2227 -7049
rect 1827 -7119 1837 -7059
rect 1897 -7119 2157 -7059
rect 2217 -7119 2227 -7059
rect 1827 -7229 2227 -7119
rect 2283 -7059 2683 -7049
rect 2283 -7119 2293 -7059
rect 2353 -7119 2613 -7059
rect 2673 -7119 2683 -7059
rect 2283 -7229 2683 -7119
rect 457 -7232 2683 -7229
rect 2741 -7059 3141 -7049
rect 2741 -7119 2751 -7059
rect 2811 -7119 3071 -7059
rect 3131 -7119 3141 -7059
rect 2741 -7229 3141 -7119
rect 3197 -7059 3597 -7049
rect 3197 -7119 3207 -7059
rect 3267 -7119 3527 -7059
rect 3587 -7119 3597 -7059
rect 3197 -7229 3597 -7119
rect 3653 -7059 4053 -7049
rect 3653 -7119 3663 -7059
rect 3723 -7119 3983 -7059
rect 4043 -7119 4053 -7059
rect 3653 -7229 4053 -7119
rect 2741 -7232 4053 -7229
rect 457 -7302 4053 -7232
rect 457 -7409 857 -7302
rect 457 -7469 467 -7409
rect 527 -7469 787 -7409
rect 847 -7469 857 -7409
rect 457 -7479 857 -7469
rect 913 -7409 1313 -7302
rect 913 -7469 923 -7409
rect 983 -7469 1243 -7409
rect 1303 -7469 1313 -7409
rect 913 -7479 1313 -7469
rect 1371 -7409 1771 -7302
rect 1371 -7469 1381 -7409
rect 1441 -7469 1701 -7409
rect 1761 -7469 1771 -7409
rect 1371 -7479 1771 -7469
rect 1827 -7409 2227 -7302
rect 1827 -7469 1837 -7409
rect 1897 -7469 2157 -7409
rect 2217 -7469 2227 -7409
rect 1827 -7479 2227 -7469
rect 2283 -7409 2683 -7302
rect 2283 -7469 2293 -7409
rect 2353 -7469 2613 -7409
rect 2673 -7469 2683 -7409
rect 2283 -7479 2683 -7469
rect 2741 -7409 3141 -7302
rect 2741 -7469 2751 -7409
rect 2811 -7469 3071 -7409
rect 3131 -7469 3141 -7409
rect 2741 -7479 3141 -7469
rect 3197 -7409 3597 -7302
rect 3197 -7469 3207 -7409
rect 3267 -7469 3527 -7409
rect 3587 -7469 3597 -7409
rect 3197 -7479 3597 -7469
rect 3653 -7409 4053 -7302
rect 3653 -7469 3663 -7409
rect 3723 -7469 3983 -7409
rect 4043 -7469 4053 -7409
rect 3653 -7479 4053 -7469
rect 4111 -7059 4511 -7049
rect 4111 -7119 4121 -7059
rect 4181 -7119 4441 -7059
rect 4501 -7119 4511 -7059
rect 4111 -7229 4511 -7119
rect 4567 -7059 4967 -7049
rect 4567 -7119 4577 -7059
rect 4637 -7119 4897 -7059
rect 4957 -7119 4967 -7059
rect 4567 -7229 4967 -7119
rect 5023 -7059 5423 -7049
rect 5023 -7119 5033 -7059
rect 5093 -7119 5353 -7059
rect 5413 -7119 5423 -7059
rect 5023 -7229 5423 -7119
rect 5481 -7059 5881 -7049
rect 5481 -7119 5491 -7059
rect 5551 -7119 5811 -7059
rect 5871 -7119 5881 -7059
rect 5481 -7229 5881 -7119
rect 5937 -7059 6337 -7049
rect 5937 -7119 5947 -7059
rect 6007 -7119 6267 -7059
rect 6327 -7119 6337 -7059
rect 5937 -7229 6337 -7119
rect 6393 -7059 6793 -7049
rect 6393 -7119 6403 -7059
rect 6463 -7119 6723 -7059
rect 6783 -7119 6793 -7059
rect 6393 -7229 6793 -7119
rect 6851 -7059 7251 -7049
rect 6851 -7119 6861 -7059
rect 6921 -7119 7181 -7059
rect 7241 -7119 7251 -7059
rect 6851 -7229 7251 -7119
rect 7307 -7059 7707 -7049
rect 7307 -7119 7317 -7059
rect 7377 -7119 7637 -7059
rect 7697 -7119 7707 -7059
rect 7307 -7229 7707 -7119
rect 7763 -7059 8163 -7049
rect 7763 -7119 7773 -7059
rect 7833 -7119 8093 -7059
rect 8153 -7119 8163 -7059
rect 7763 -7229 8163 -7119
rect 8237 -7059 8637 -7049
rect 8237 -7119 8247 -7059
rect 8307 -7119 8567 -7059
rect 8627 -7119 8637 -7059
rect 8237 -7229 8637 -7119
rect 8693 -7059 9093 -7049
rect 8693 -7119 8703 -7059
rect 8763 -7119 9023 -7059
rect 9083 -7119 9093 -7059
rect 8693 -7229 9093 -7119
rect 9151 -7059 9551 -7049
rect 9151 -7119 9161 -7059
rect 9221 -7119 9481 -7059
rect 9541 -7119 9551 -7059
rect 9151 -7229 9551 -7119
rect 9607 -7059 10007 -7049
rect 9607 -7119 9617 -7059
rect 9677 -7119 9937 -7059
rect 9997 -7119 10007 -7059
rect 9607 -7229 10007 -7119
rect 10063 -7059 10463 -7049
rect 10063 -7119 10073 -7059
rect 10133 -7119 10393 -7059
rect 10453 -7119 10463 -7059
rect 10063 -7229 10463 -7119
rect 4111 -7232 10463 -7229
rect 10521 -7059 10921 -7049
rect 10521 -7119 10531 -7059
rect 10591 -7119 10851 -7059
rect 10911 -7119 10921 -7059
rect 10521 -7229 10921 -7119
rect 10977 -7059 11377 -7049
rect 10977 -7119 10987 -7059
rect 11047 -7119 11307 -7059
rect 11367 -7119 11377 -7059
rect 10977 -7229 11377 -7119
rect 11433 -7059 11833 -7049
rect 11433 -7119 11443 -7059
rect 11503 -7119 11763 -7059
rect 11823 -7119 11833 -7059
rect 11433 -7229 11833 -7119
rect 11891 -7059 12291 -7049
rect 11891 -7119 11901 -7059
rect 11961 -7119 12221 -7059
rect 12281 -7119 12291 -7059
rect 11891 -7229 12291 -7119
rect 12347 -7059 12747 -7049
rect 12347 -7119 12357 -7059
rect 12417 -7119 12677 -7059
rect 12737 -7119 12747 -7059
rect 12347 -7229 12747 -7119
rect 12803 -7059 13203 -7049
rect 12803 -7119 12813 -7059
rect 12873 -7119 13133 -7059
rect 13193 -7119 13203 -7059
rect 12803 -7229 13203 -7119
rect 13261 -7059 13661 -7049
rect 13261 -7119 13271 -7059
rect 13331 -7119 13591 -7059
rect 13651 -7119 13661 -7059
rect 13261 -7229 13661 -7119
rect 13717 -7059 14117 -7049
rect 13717 -7119 13727 -7059
rect 13787 -7119 14047 -7059
rect 14107 -7119 14117 -7059
rect 13717 -7229 14117 -7119
rect 14173 -7059 14573 -7049
rect 14173 -7119 14183 -7059
rect 14243 -7119 14503 -7059
rect 14563 -7119 14573 -7059
rect 14173 -7229 14573 -7119
rect 14631 -7059 15031 -7049
rect 14631 -7119 14641 -7059
rect 14701 -7119 14961 -7059
rect 15021 -7119 15031 -7059
rect 14631 -7229 15031 -7119
rect 15087 -7059 15487 -7049
rect 15087 -7119 15097 -7059
rect 15157 -7119 15417 -7059
rect 15477 -7119 15487 -7059
rect 15087 -7229 15487 -7119
rect 10521 -7232 15487 -7229
rect 4111 -7302 15487 -7232
rect 4111 -7409 4511 -7302
rect 4111 -7469 4121 -7409
rect 4181 -7469 4441 -7409
rect 4501 -7469 4511 -7409
rect 4111 -7479 4511 -7469
rect 4567 -7409 4967 -7302
rect 4567 -7469 4577 -7409
rect 4637 -7469 4897 -7409
rect 4957 -7469 4967 -7409
rect 4567 -7479 4967 -7469
rect 5023 -7409 5423 -7302
rect 5023 -7469 5033 -7409
rect 5093 -7469 5353 -7409
rect 5413 -7469 5423 -7409
rect 5023 -7479 5423 -7469
rect 5481 -7409 5881 -7302
rect 5481 -7469 5491 -7409
rect 5551 -7469 5811 -7409
rect 5871 -7469 5881 -7409
rect 5481 -7479 5881 -7469
rect 5937 -7409 6337 -7302
rect 5937 -7469 5947 -7409
rect 6007 -7469 6267 -7409
rect 6327 -7469 6337 -7409
rect 5937 -7479 6337 -7469
rect 6393 -7409 6793 -7302
rect 6393 -7469 6403 -7409
rect 6463 -7469 6723 -7409
rect 6783 -7469 6793 -7409
rect 6393 -7479 6793 -7469
rect 6851 -7409 7251 -7302
rect 6851 -7469 6861 -7409
rect 6921 -7469 7181 -7409
rect 7241 -7469 7251 -7409
rect 6851 -7479 7251 -7469
rect 7307 -7409 7707 -7302
rect 7307 -7469 7317 -7409
rect 7377 -7469 7637 -7409
rect 7697 -7469 7707 -7409
rect 7307 -7479 7707 -7469
rect 7763 -7409 8163 -7302
rect 7763 -7469 7773 -7409
rect 7833 -7469 8093 -7409
rect 8153 -7469 8163 -7409
rect 7763 -7479 8163 -7469
rect 8237 -7409 8637 -7302
rect 8237 -7469 8247 -7409
rect 8307 -7469 8567 -7409
rect 8627 -7469 8637 -7409
rect 8237 -7479 8637 -7469
rect 8693 -7409 9093 -7302
rect 8693 -7469 8703 -7409
rect 8763 -7469 9023 -7409
rect 9083 -7469 9093 -7409
rect 8693 -7479 9093 -7469
rect 9151 -7409 9551 -7302
rect 9151 -7469 9161 -7409
rect 9221 -7469 9481 -7409
rect 9541 -7469 9551 -7409
rect 9151 -7479 9551 -7469
rect 9607 -7409 10007 -7302
rect 9607 -7469 9617 -7409
rect 9677 -7469 9937 -7409
rect 9997 -7469 10007 -7409
rect 9607 -7479 10007 -7469
rect 10063 -7409 10463 -7302
rect 10063 -7469 10073 -7409
rect 10133 -7469 10393 -7409
rect 10453 -7469 10463 -7409
rect 10063 -7479 10463 -7469
rect 10521 -7409 10921 -7302
rect 10521 -7469 10531 -7409
rect 10591 -7469 10851 -7409
rect 10911 -7469 10921 -7409
rect 10521 -7479 10921 -7469
rect 10977 -7409 11377 -7302
rect 10977 -7469 10987 -7409
rect 11047 -7469 11307 -7409
rect 11367 -7469 11377 -7409
rect 10977 -7479 11377 -7469
rect 11433 -7409 11833 -7302
rect 11433 -7469 11443 -7409
rect 11503 -7469 11763 -7409
rect 11823 -7469 11833 -7409
rect 11433 -7479 11833 -7469
rect 11891 -7409 12291 -7302
rect 11891 -7469 11901 -7409
rect 11961 -7469 12221 -7409
rect 12281 -7469 12291 -7409
rect 11891 -7479 12291 -7469
rect 12347 -7409 12747 -7302
rect 12347 -7469 12357 -7409
rect 12417 -7469 12677 -7409
rect 12737 -7469 12747 -7409
rect 12347 -7479 12747 -7469
rect 12803 -7409 13203 -7302
rect 12803 -7469 12813 -7409
rect 12873 -7469 13133 -7409
rect 13193 -7469 13203 -7409
rect 12803 -7479 13203 -7469
rect 13261 -7409 13661 -7302
rect 13261 -7469 13271 -7409
rect 13331 -7469 13591 -7409
rect 13651 -7469 13661 -7409
rect 13261 -7479 13661 -7469
rect 13717 -7409 14117 -7302
rect 13717 -7469 13727 -7409
rect 13787 -7469 14047 -7409
rect 14107 -7469 14117 -7409
rect 13717 -7479 14117 -7469
rect 14173 -7409 14573 -7302
rect 14173 -7469 14183 -7409
rect 14243 -7469 14503 -7409
rect 14563 -7469 14573 -7409
rect 14173 -7479 14573 -7469
rect 14631 -7409 15031 -7302
rect 14631 -7469 14641 -7409
rect 14701 -7469 14961 -7409
rect 15021 -7469 15031 -7409
rect 14631 -7479 15031 -7469
rect 15087 -7409 15487 -7302
rect 15087 -7469 15097 -7409
rect 15157 -7469 15417 -7409
rect 15477 -7469 15487 -7409
rect 15087 -7479 15487 -7469
rect 66 -7551 80 -7479
rect 457 -7551 527 -7479
rect 913 -7551 984 -7479
rect 1371 -7551 1442 -7479
rect 1827 -7551 1898 -7479
rect 2283 -7551 2354 -7479
rect 2741 -7551 2812 -7479
rect 3197 -7551 3268 -7479
rect 3653 -7551 3724 -7479
rect 4111 -7551 4182 -7479
rect 4567 -7551 4638 -7479
rect 5023 -7551 5094 -7479
rect 5481 -7551 5552 -7479
rect 5937 -7551 6008 -7479
rect 6393 -7551 6464 -7479
rect 6851 -7551 6922 -7479
rect 7307 -7551 7378 -7479
rect 7763 -7551 7834 -7479
rect 8237 -7551 8308 -7479
rect 8693 -7551 8764 -7479
rect 9151 -7551 9222 -7479
rect 9607 -7551 9678 -7479
rect 10063 -7551 10134 -7479
rect 10521 -7551 10592 -7479
rect 10977 -7551 11048 -7479
rect 11433 -7551 11504 -7479
rect 11891 -7551 11962 -7479
rect 12347 -7551 12418 -7479
rect 12803 -7551 12874 -7479
rect 13261 -7551 13332 -7479
rect 13717 -7551 13788 -7479
rect 14173 -7551 14244 -7479
rect 14631 -7551 14702 -7479
rect 66 -7561 400 -7551
rect 0 -7621 11 -7561
rect 71 -7621 331 -7561
rect 391 -7621 400 -7561
rect 0 -7911 14 -7621
rect 66 -7911 400 -7621
rect 0 -7971 11 -7911
rect 71 -7971 331 -7911
rect 391 -7971 400 -7911
rect 0 -8053 14 -7971
rect 66 -7981 400 -7971
rect 457 -7561 857 -7551
rect 457 -7621 467 -7561
rect 527 -7621 787 -7561
rect 847 -7621 857 -7561
rect 457 -7731 857 -7621
rect 913 -7561 1313 -7551
rect 913 -7621 923 -7561
rect 983 -7621 1243 -7561
rect 1303 -7621 1313 -7561
rect 913 -7731 1313 -7621
rect 1371 -7561 1771 -7551
rect 1371 -7621 1381 -7561
rect 1441 -7621 1701 -7561
rect 1761 -7621 1771 -7561
rect 1371 -7731 1771 -7621
rect 1827 -7561 2227 -7551
rect 1827 -7621 1837 -7561
rect 1897 -7621 2157 -7561
rect 2217 -7621 2227 -7561
rect 1827 -7731 2227 -7621
rect 2283 -7561 2683 -7551
rect 2283 -7621 2293 -7561
rect 2353 -7621 2613 -7561
rect 2673 -7621 2683 -7561
rect 2283 -7731 2683 -7621
rect 457 -7732 2683 -7731
rect 2741 -7561 3141 -7551
rect 2741 -7621 2751 -7561
rect 2811 -7621 3071 -7561
rect 3131 -7621 3141 -7561
rect 2741 -7731 3141 -7621
rect 3197 -7561 3597 -7551
rect 3197 -7621 3207 -7561
rect 3267 -7621 3527 -7561
rect 3587 -7621 3597 -7561
rect 3197 -7731 3597 -7621
rect 3653 -7561 4053 -7551
rect 3653 -7621 3663 -7561
rect 3723 -7621 3983 -7561
rect 4043 -7621 4053 -7561
rect 3653 -7731 4053 -7621
rect 2741 -7732 4053 -7731
rect 457 -7802 4053 -7732
rect 457 -7911 857 -7802
rect 457 -7971 467 -7911
rect 527 -7971 787 -7911
rect 847 -7971 857 -7911
rect 457 -7981 857 -7971
rect 913 -7911 1313 -7802
rect 913 -7971 923 -7911
rect 983 -7971 1243 -7911
rect 1303 -7971 1313 -7911
rect 913 -7981 1313 -7971
rect 1371 -7911 1771 -7802
rect 1371 -7971 1381 -7911
rect 1441 -7971 1701 -7911
rect 1761 -7971 1771 -7911
rect 1371 -7981 1771 -7971
rect 1827 -7911 2227 -7802
rect 1827 -7971 1837 -7911
rect 1897 -7971 2157 -7911
rect 2217 -7971 2227 -7911
rect 1827 -7981 2227 -7971
rect 2283 -7911 2683 -7802
rect 2283 -7971 2293 -7911
rect 2353 -7971 2613 -7911
rect 2673 -7971 2683 -7911
rect 2283 -7981 2683 -7971
rect 2741 -7911 3141 -7802
rect 2741 -7971 2751 -7911
rect 2811 -7971 3071 -7911
rect 3131 -7971 3141 -7911
rect 2741 -7981 3141 -7971
rect 3197 -7911 3597 -7802
rect 3197 -7971 3207 -7911
rect 3267 -7971 3527 -7911
rect 3587 -7971 3597 -7911
rect 3197 -7981 3597 -7971
rect 3653 -7911 4053 -7802
rect 3653 -7971 3663 -7911
rect 3723 -7971 3983 -7911
rect 4043 -7971 4053 -7911
rect 3653 -7981 4053 -7971
rect 4111 -7561 4511 -7551
rect 4111 -7621 4121 -7561
rect 4181 -7621 4441 -7561
rect 4501 -7621 4511 -7561
rect 4111 -7731 4511 -7621
rect 4567 -7561 4967 -7551
rect 4567 -7621 4577 -7561
rect 4637 -7621 4897 -7561
rect 4957 -7621 4967 -7561
rect 4567 -7731 4967 -7621
rect 5023 -7561 5423 -7551
rect 5023 -7621 5033 -7561
rect 5093 -7621 5353 -7561
rect 5413 -7621 5423 -7561
rect 5023 -7731 5423 -7621
rect 5481 -7561 5881 -7551
rect 5481 -7621 5491 -7561
rect 5551 -7621 5811 -7561
rect 5871 -7621 5881 -7561
rect 5481 -7731 5881 -7621
rect 5937 -7561 6337 -7551
rect 5937 -7621 5947 -7561
rect 6007 -7621 6267 -7561
rect 6327 -7621 6337 -7561
rect 5937 -7731 6337 -7621
rect 6393 -7561 6793 -7551
rect 6393 -7621 6403 -7561
rect 6463 -7621 6723 -7561
rect 6783 -7621 6793 -7561
rect 6393 -7731 6793 -7621
rect 6851 -7561 7251 -7551
rect 6851 -7621 6861 -7561
rect 6921 -7621 7181 -7561
rect 7241 -7621 7251 -7561
rect 6851 -7731 7251 -7621
rect 7307 -7561 7707 -7551
rect 7307 -7621 7317 -7561
rect 7377 -7621 7637 -7561
rect 7697 -7621 7707 -7561
rect 7307 -7731 7707 -7621
rect 7763 -7561 8163 -7551
rect 7763 -7621 7773 -7561
rect 7833 -7621 8093 -7561
rect 8153 -7621 8163 -7561
rect 7763 -7731 8163 -7621
rect 8237 -7561 8637 -7551
rect 8237 -7621 8247 -7561
rect 8307 -7621 8567 -7561
rect 8627 -7621 8637 -7561
rect 8237 -7731 8637 -7621
rect 8693 -7561 9093 -7551
rect 8693 -7621 8703 -7561
rect 8763 -7621 9023 -7561
rect 9083 -7621 9093 -7561
rect 8693 -7731 9093 -7621
rect 9151 -7561 9551 -7551
rect 9151 -7621 9161 -7561
rect 9221 -7621 9481 -7561
rect 9541 -7621 9551 -7561
rect 9151 -7731 9551 -7621
rect 9607 -7561 10007 -7551
rect 9607 -7621 9617 -7561
rect 9677 -7621 9937 -7561
rect 9997 -7621 10007 -7561
rect 9607 -7731 10007 -7621
rect 10063 -7561 10463 -7551
rect 10063 -7621 10073 -7561
rect 10133 -7621 10393 -7561
rect 10453 -7621 10463 -7561
rect 10063 -7731 10463 -7621
rect 4111 -7732 10463 -7731
rect 10521 -7561 10921 -7551
rect 10521 -7621 10531 -7561
rect 10591 -7621 10851 -7561
rect 10911 -7621 10921 -7561
rect 10521 -7731 10921 -7621
rect 10977 -7561 11377 -7551
rect 10977 -7621 10987 -7561
rect 11047 -7621 11307 -7561
rect 11367 -7621 11377 -7561
rect 10977 -7731 11377 -7621
rect 11433 -7561 11833 -7551
rect 11433 -7621 11443 -7561
rect 11503 -7621 11763 -7561
rect 11823 -7621 11833 -7561
rect 11433 -7731 11833 -7621
rect 11891 -7561 12291 -7551
rect 11891 -7621 11901 -7561
rect 11961 -7621 12221 -7561
rect 12281 -7621 12291 -7561
rect 11891 -7731 12291 -7621
rect 12347 -7561 12747 -7551
rect 12347 -7621 12357 -7561
rect 12417 -7621 12677 -7561
rect 12737 -7621 12747 -7561
rect 12347 -7731 12747 -7621
rect 12803 -7561 13203 -7551
rect 12803 -7621 12813 -7561
rect 12873 -7621 13133 -7561
rect 13193 -7621 13203 -7561
rect 12803 -7731 13203 -7621
rect 13261 -7561 13661 -7551
rect 13261 -7621 13271 -7561
rect 13331 -7621 13591 -7561
rect 13651 -7621 13661 -7561
rect 13261 -7731 13661 -7621
rect 13717 -7561 14117 -7551
rect 13717 -7621 13727 -7561
rect 13787 -7621 14047 -7561
rect 14107 -7621 14117 -7561
rect 13717 -7731 14117 -7621
rect 14173 -7561 14573 -7551
rect 14173 -7621 14183 -7561
rect 14243 -7621 14503 -7561
rect 14563 -7621 14573 -7561
rect 14173 -7731 14573 -7621
rect 14631 -7561 15031 -7551
rect 14631 -7621 14641 -7561
rect 14701 -7621 14961 -7561
rect 15021 -7621 15031 -7561
rect 14631 -7731 15031 -7621
rect 15087 -7561 15487 -7551
rect 15087 -7621 15097 -7561
rect 15157 -7621 15417 -7561
rect 15477 -7621 15487 -7561
rect 15087 -7731 15487 -7621
rect 10521 -7732 15487 -7731
rect 4111 -7802 15487 -7732
rect 4111 -7911 4511 -7802
rect 4111 -7971 4121 -7911
rect 4181 -7971 4441 -7911
rect 4501 -7971 4511 -7911
rect 4111 -7981 4511 -7971
rect 4567 -7911 4967 -7802
rect 4567 -7971 4577 -7911
rect 4637 -7971 4897 -7911
rect 4957 -7971 4967 -7911
rect 4567 -7981 4967 -7971
rect 5023 -7911 5423 -7802
rect 5023 -7971 5033 -7911
rect 5093 -7971 5353 -7911
rect 5413 -7971 5423 -7911
rect 5023 -7981 5423 -7971
rect 5481 -7911 5881 -7802
rect 5481 -7971 5491 -7911
rect 5551 -7971 5811 -7911
rect 5871 -7971 5881 -7911
rect 5481 -7981 5881 -7971
rect 5937 -7911 6337 -7802
rect 5937 -7971 5947 -7911
rect 6007 -7971 6267 -7911
rect 6327 -7971 6337 -7911
rect 5937 -7981 6337 -7971
rect 6393 -7911 6793 -7802
rect 6393 -7971 6403 -7911
rect 6463 -7971 6723 -7911
rect 6783 -7971 6793 -7911
rect 6393 -7981 6793 -7971
rect 6851 -7911 7251 -7802
rect 6851 -7971 6861 -7911
rect 6921 -7971 7181 -7911
rect 7241 -7971 7251 -7911
rect 6851 -7981 7251 -7971
rect 7307 -7911 7707 -7802
rect 7307 -7971 7317 -7911
rect 7377 -7971 7637 -7911
rect 7697 -7971 7707 -7911
rect 7307 -7981 7707 -7971
rect 7763 -7911 8163 -7802
rect 7763 -7971 7773 -7911
rect 7833 -7971 8093 -7911
rect 8153 -7971 8163 -7911
rect 7763 -7981 8163 -7971
rect 8237 -7911 8637 -7802
rect 8237 -7971 8247 -7911
rect 8307 -7971 8567 -7911
rect 8627 -7971 8637 -7911
rect 8237 -7981 8637 -7971
rect 8693 -7911 9093 -7802
rect 8693 -7971 8703 -7911
rect 8763 -7971 9023 -7911
rect 9083 -7971 9093 -7911
rect 8693 -7981 9093 -7971
rect 9151 -7911 9551 -7802
rect 9151 -7971 9161 -7911
rect 9221 -7971 9481 -7911
rect 9541 -7971 9551 -7911
rect 9151 -7981 9551 -7971
rect 9607 -7911 10007 -7802
rect 9607 -7971 9617 -7911
rect 9677 -7971 9937 -7911
rect 9997 -7971 10007 -7911
rect 9607 -7981 10007 -7971
rect 10063 -7911 10463 -7802
rect 10063 -7971 10073 -7911
rect 10133 -7971 10393 -7911
rect 10453 -7971 10463 -7911
rect 10063 -7981 10463 -7971
rect 10521 -7911 10921 -7802
rect 10521 -7971 10531 -7911
rect 10591 -7971 10851 -7911
rect 10911 -7971 10921 -7911
rect 10521 -7981 10921 -7971
rect 10977 -7911 11377 -7802
rect 10977 -7971 10987 -7911
rect 11047 -7971 11307 -7911
rect 11367 -7971 11377 -7911
rect 10977 -7981 11377 -7971
rect 11433 -7911 11833 -7802
rect 11433 -7971 11443 -7911
rect 11503 -7971 11763 -7911
rect 11823 -7971 11833 -7911
rect 11433 -7981 11833 -7971
rect 11891 -7911 12291 -7802
rect 11891 -7971 11901 -7911
rect 11961 -7971 12221 -7911
rect 12281 -7971 12291 -7911
rect 11891 -7981 12291 -7971
rect 12347 -7911 12747 -7802
rect 12347 -7971 12357 -7911
rect 12417 -7971 12677 -7911
rect 12737 -7971 12747 -7911
rect 12347 -7981 12747 -7971
rect 12803 -7911 13203 -7802
rect 12803 -7971 12813 -7911
rect 12873 -7971 13133 -7911
rect 13193 -7971 13203 -7911
rect 12803 -7981 13203 -7971
rect 13261 -7911 13661 -7802
rect 13261 -7971 13271 -7911
rect 13331 -7971 13591 -7911
rect 13651 -7971 13661 -7911
rect 13261 -7981 13661 -7971
rect 13717 -7911 14117 -7802
rect 13717 -7971 13727 -7911
rect 13787 -7971 14047 -7911
rect 14107 -7971 14117 -7911
rect 13717 -7981 14117 -7971
rect 14173 -7911 14573 -7802
rect 14173 -7971 14183 -7911
rect 14243 -7971 14503 -7911
rect 14563 -7971 14573 -7911
rect 14173 -7981 14573 -7971
rect 14631 -7911 15031 -7802
rect 14631 -7971 14641 -7911
rect 14701 -7971 14961 -7911
rect 15021 -7971 15031 -7911
rect 14631 -7981 15031 -7971
rect 15087 -7911 15487 -7802
rect 15087 -7971 15097 -7911
rect 15157 -7971 15417 -7911
rect 15477 -7971 15487 -7911
rect 15087 -7981 15487 -7971
rect 66 -8043 80 -7981
rect 457 -8043 528 -7981
rect 913 -8043 984 -7981
rect 1371 -8043 1442 -7981
rect 1827 -8043 1898 -7981
rect 2283 -8043 2354 -7981
rect 2741 -8043 2811 -7981
rect 3197 -8043 3267 -7981
rect 3653 -8043 3723 -7981
rect 4111 -8043 4181 -7981
rect 4567 -8043 4637 -7981
rect 5023 -8043 5093 -7981
rect 5481 -8043 5551 -7981
rect 5937 -8043 6007 -7981
rect 6393 -8043 6463 -7981
rect 6851 -8043 6921 -7981
rect 7307 -8043 7377 -7981
rect 7763 -8043 7833 -7981
rect 8237 -8043 8307 -7981
rect 8693 -8043 8763 -7981
rect 9151 -8043 9221 -7981
rect 9607 -8043 9677 -7981
rect 10063 -8043 10133 -7981
rect 10521 -8043 10591 -7981
rect 10977 -8043 11047 -7981
rect 11433 -8043 11503 -7981
rect 11891 -8043 11961 -7981
rect 12347 -8043 12417 -7981
rect 12803 -8043 12873 -7981
rect 13261 -8043 13331 -7981
rect 13717 -8043 13787 -7981
rect 14173 -8043 14243 -7981
rect 14631 -8043 14701 -7981
rect 66 -8053 400 -8043
rect 0 -8113 11 -8053
rect 71 -8113 331 -8053
rect 391 -8113 400 -8053
rect 0 -8403 14 -8113
rect 66 -8403 400 -8113
rect 0 -8463 11 -8403
rect 71 -8463 331 -8403
rect 391 -8463 400 -8403
rect 0 -8547 14 -8463
rect 66 -8473 400 -8463
rect 457 -8053 857 -8043
rect 457 -8113 467 -8053
rect 527 -8113 787 -8053
rect 847 -8113 857 -8053
rect 457 -8222 857 -8113
rect 913 -8053 1313 -8043
rect 913 -8113 923 -8053
rect 983 -8113 1243 -8053
rect 1303 -8113 1313 -8053
rect 913 -8222 1313 -8113
rect 1371 -8053 1771 -8043
rect 1371 -8113 1381 -8053
rect 1441 -8113 1701 -8053
rect 1761 -8113 1771 -8053
rect 1371 -8222 1771 -8113
rect 1827 -8053 2227 -8043
rect 1827 -8113 1837 -8053
rect 1897 -8113 2157 -8053
rect 2217 -8113 2227 -8053
rect 1827 -8222 2227 -8113
rect 2283 -8053 2683 -8043
rect 2283 -8113 2293 -8053
rect 2353 -8113 2613 -8053
rect 2673 -8113 2683 -8053
rect 2283 -8222 2683 -8113
rect 2741 -8053 3141 -8043
rect 2741 -8113 2751 -8053
rect 2811 -8113 3071 -8053
rect 3131 -8113 3141 -8053
rect 2741 -8222 3141 -8113
rect 3197 -8053 3597 -8043
rect 3197 -8113 3207 -8053
rect 3267 -8113 3527 -8053
rect 3587 -8113 3597 -8053
rect 3197 -8222 3597 -8113
rect 3653 -8053 4053 -8043
rect 3653 -8113 3663 -8053
rect 3723 -8113 3983 -8053
rect 4043 -8113 4053 -8053
rect 3653 -8222 4053 -8113
rect 457 -8292 4053 -8222
rect 457 -8293 2683 -8292
rect 457 -8403 857 -8293
rect 457 -8463 467 -8403
rect 527 -8463 787 -8403
rect 847 -8463 857 -8403
rect 457 -8473 857 -8463
rect 913 -8403 1313 -8293
rect 913 -8463 923 -8403
rect 983 -8463 1243 -8403
rect 1303 -8463 1313 -8403
rect 913 -8473 1313 -8463
rect 1371 -8403 1771 -8293
rect 1371 -8463 1381 -8403
rect 1441 -8463 1701 -8403
rect 1761 -8463 1771 -8403
rect 1371 -8473 1771 -8463
rect 1827 -8403 2227 -8293
rect 1827 -8463 1837 -8403
rect 1897 -8463 2157 -8403
rect 2217 -8463 2227 -8403
rect 1827 -8473 2227 -8463
rect 2283 -8403 2683 -8293
rect 2283 -8463 2293 -8403
rect 2353 -8463 2613 -8403
rect 2673 -8463 2683 -8403
rect 2283 -8473 2683 -8463
rect 2741 -8293 4053 -8292
rect 2741 -8403 3141 -8293
rect 2741 -8463 2751 -8403
rect 2811 -8463 3071 -8403
rect 3131 -8463 3141 -8403
rect 2741 -8473 3141 -8463
rect 3197 -8403 3597 -8293
rect 3197 -8463 3207 -8403
rect 3267 -8463 3527 -8403
rect 3587 -8463 3597 -8403
rect 3197 -8473 3597 -8463
rect 3653 -8403 4053 -8293
rect 3653 -8463 3663 -8403
rect 3723 -8463 3983 -8403
rect 4043 -8463 4053 -8403
rect 3653 -8473 4053 -8463
rect 4111 -8053 4511 -8043
rect 4111 -8113 4121 -8053
rect 4181 -8113 4441 -8053
rect 4501 -8113 4511 -8053
rect 4111 -8222 4511 -8113
rect 4567 -8053 4967 -8043
rect 4567 -8113 4577 -8053
rect 4637 -8113 4897 -8053
rect 4957 -8113 4967 -8053
rect 4567 -8222 4967 -8113
rect 5023 -8053 5423 -8043
rect 5023 -8113 5033 -8053
rect 5093 -8113 5353 -8053
rect 5413 -8113 5423 -8053
rect 5023 -8222 5423 -8113
rect 5481 -8053 5881 -8043
rect 5481 -8113 5491 -8053
rect 5551 -8113 5811 -8053
rect 5871 -8113 5881 -8053
rect 5481 -8222 5881 -8113
rect 5937 -8053 6337 -8043
rect 5937 -8113 5947 -8053
rect 6007 -8113 6267 -8053
rect 6327 -8113 6337 -8053
rect 5937 -8222 6337 -8113
rect 6393 -8053 6793 -8043
rect 6393 -8113 6403 -8053
rect 6463 -8113 6723 -8053
rect 6783 -8113 6793 -8053
rect 6393 -8222 6793 -8113
rect 6851 -8053 7251 -8043
rect 6851 -8113 6861 -8053
rect 6921 -8113 7181 -8053
rect 7241 -8113 7251 -8053
rect 6851 -8222 7251 -8113
rect 7307 -8053 7707 -8043
rect 7307 -8113 7317 -8053
rect 7377 -8113 7637 -8053
rect 7697 -8113 7707 -8053
rect 7307 -8222 7707 -8113
rect 7763 -8053 8163 -8043
rect 7763 -8113 7773 -8053
rect 7833 -8113 8093 -8053
rect 8153 -8113 8163 -8053
rect 7763 -8222 8163 -8113
rect 8237 -8053 8637 -8043
rect 8237 -8113 8247 -8053
rect 8307 -8113 8567 -8053
rect 8627 -8113 8637 -8053
rect 8237 -8222 8637 -8113
rect 8693 -8053 9093 -8043
rect 8693 -8113 8703 -8053
rect 8763 -8113 9023 -8053
rect 9083 -8113 9093 -8053
rect 8693 -8222 9093 -8113
rect 9151 -8053 9551 -8043
rect 9151 -8113 9161 -8053
rect 9221 -8113 9481 -8053
rect 9541 -8113 9551 -8053
rect 9151 -8222 9551 -8113
rect 9607 -8053 10007 -8043
rect 9607 -8113 9617 -8053
rect 9677 -8113 9937 -8053
rect 9997 -8113 10007 -8053
rect 9607 -8222 10007 -8113
rect 10063 -8053 10463 -8043
rect 10063 -8113 10073 -8053
rect 10133 -8113 10393 -8053
rect 10453 -8113 10463 -8053
rect 10063 -8222 10463 -8113
rect 10521 -8053 10921 -8043
rect 10521 -8113 10531 -8053
rect 10591 -8113 10851 -8053
rect 10911 -8113 10921 -8053
rect 10521 -8222 10921 -8113
rect 10977 -8053 11377 -8043
rect 10977 -8113 10987 -8053
rect 11047 -8113 11307 -8053
rect 11367 -8113 11377 -8053
rect 10977 -8222 11377 -8113
rect 11433 -8053 11833 -8043
rect 11433 -8113 11443 -8053
rect 11503 -8113 11763 -8053
rect 11823 -8113 11833 -8053
rect 11433 -8222 11833 -8113
rect 11891 -8053 12291 -8043
rect 11891 -8113 11901 -8053
rect 11961 -8113 12221 -8053
rect 12281 -8113 12291 -8053
rect 11891 -8222 12291 -8113
rect 12347 -8053 12747 -8043
rect 12347 -8113 12357 -8053
rect 12417 -8113 12677 -8053
rect 12737 -8113 12747 -8053
rect 12347 -8222 12747 -8113
rect 12803 -8053 13203 -8043
rect 12803 -8113 12813 -8053
rect 12873 -8113 13133 -8053
rect 13193 -8113 13203 -8053
rect 12803 -8222 13203 -8113
rect 13261 -8053 13661 -8043
rect 13261 -8113 13271 -8053
rect 13331 -8113 13591 -8053
rect 13651 -8113 13661 -8053
rect 13261 -8222 13661 -8113
rect 13717 -8053 14117 -8043
rect 13717 -8113 13727 -8053
rect 13787 -8113 14047 -8053
rect 14107 -8113 14117 -8053
rect 13717 -8222 14117 -8113
rect 14173 -8053 14573 -8043
rect 14173 -8113 14183 -8053
rect 14243 -8113 14503 -8053
rect 14563 -8113 14573 -8053
rect 14173 -8222 14573 -8113
rect 14631 -8053 15031 -8043
rect 14631 -8113 14641 -8053
rect 14701 -8113 14961 -8053
rect 15021 -8113 15031 -8053
rect 14631 -8222 15031 -8113
rect 15087 -8053 15487 -8043
rect 15087 -8113 15097 -8053
rect 15157 -8113 15417 -8053
rect 15477 -8113 15487 -8053
rect 15087 -8222 15487 -8113
rect 4111 -8292 15487 -8222
rect 4111 -8293 10463 -8292
rect 4111 -8403 4511 -8293
rect 4111 -8463 4121 -8403
rect 4181 -8463 4441 -8403
rect 4501 -8463 4511 -8403
rect 4111 -8473 4511 -8463
rect 4567 -8403 4967 -8293
rect 4567 -8463 4577 -8403
rect 4637 -8463 4897 -8403
rect 4957 -8463 4967 -8403
rect 4567 -8473 4967 -8463
rect 5023 -8403 5423 -8293
rect 5023 -8463 5033 -8403
rect 5093 -8463 5353 -8403
rect 5413 -8463 5423 -8403
rect 5023 -8473 5423 -8463
rect 5481 -8403 5881 -8293
rect 5481 -8463 5491 -8403
rect 5551 -8463 5811 -8403
rect 5871 -8463 5881 -8403
rect 5481 -8473 5881 -8463
rect 5937 -8403 6337 -8293
rect 5937 -8463 5947 -8403
rect 6007 -8463 6267 -8403
rect 6327 -8463 6337 -8403
rect 5937 -8473 6337 -8463
rect 6393 -8403 6793 -8293
rect 6393 -8463 6403 -8403
rect 6463 -8463 6723 -8403
rect 6783 -8463 6793 -8403
rect 6393 -8473 6793 -8463
rect 6851 -8403 7251 -8293
rect 6851 -8463 6861 -8403
rect 6921 -8463 7181 -8403
rect 7241 -8463 7251 -8403
rect 6851 -8473 7251 -8463
rect 7307 -8403 7707 -8293
rect 7307 -8463 7317 -8403
rect 7377 -8463 7637 -8403
rect 7697 -8463 7707 -8403
rect 7307 -8473 7707 -8463
rect 7763 -8403 8163 -8293
rect 7763 -8463 7773 -8403
rect 7833 -8463 8093 -8403
rect 8153 -8463 8163 -8403
rect 7763 -8473 8163 -8463
rect 8237 -8403 8637 -8293
rect 8237 -8463 8247 -8403
rect 8307 -8463 8567 -8403
rect 8627 -8463 8637 -8403
rect 8237 -8473 8637 -8463
rect 8693 -8403 9093 -8293
rect 8693 -8463 8703 -8403
rect 8763 -8463 9023 -8403
rect 9083 -8463 9093 -8403
rect 8693 -8473 9093 -8463
rect 9151 -8403 9551 -8293
rect 9151 -8463 9161 -8403
rect 9221 -8463 9481 -8403
rect 9541 -8463 9551 -8403
rect 9151 -8473 9551 -8463
rect 9607 -8403 10007 -8293
rect 9607 -8463 9617 -8403
rect 9677 -8463 9937 -8403
rect 9997 -8463 10007 -8403
rect 9607 -8473 10007 -8463
rect 10063 -8403 10463 -8293
rect 10063 -8463 10073 -8403
rect 10133 -8463 10393 -8403
rect 10453 -8463 10463 -8403
rect 10063 -8473 10463 -8463
rect 10521 -8293 15487 -8292
rect 10521 -8403 10921 -8293
rect 10521 -8463 10531 -8403
rect 10591 -8463 10851 -8403
rect 10911 -8463 10921 -8403
rect 10521 -8473 10921 -8463
rect 10977 -8403 11377 -8293
rect 10977 -8463 10987 -8403
rect 11047 -8463 11307 -8403
rect 11367 -8463 11377 -8403
rect 10977 -8473 11377 -8463
rect 11433 -8403 11833 -8293
rect 11433 -8463 11443 -8403
rect 11503 -8463 11763 -8403
rect 11823 -8463 11833 -8403
rect 11433 -8473 11833 -8463
rect 11891 -8403 12291 -8293
rect 11891 -8463 11901 -8403
rect 11961 -8463 12221 -8403
rect 12281 -8463 12291 -8403
rect 11891 -8473 12291 -8463
rect 12347 -8403 12747 -8293
rect 12347 -8463 12357 -8403
rect 12417 -8463 12677 -8403
rect 12737 -8463 12747 -8403
rect 12347 -8473 12747 -8463
rect 12803 -8403 13203 -8293
rect 12803 -8463 12813 -8403
rect 12873 -8463 13133 -8403
rect 13193 -8463 13203 -8403
rect 12803 -8473 13203 -8463
rect 13261 -8403 13661 -8293
rect 13261 -8463 13271 -8403
rect 13331 -8463 13591 -8403
rect 13651 -8463 13661 -8403
rect 13261 -8473 13661 -8463
rect 13717 -8403 14117 -8293
rect 13717 -8463 13727 -8403
rect 13787 -8463 14047 -8403
rect 14107 -8463 14117 -8403
rect 13717 -8473 14117 -8463
rect 14173 -8403 14573 -8293
rect 14173 -8463 14183 -8403
rect 14243 -8463 14503 -8403
rect 14563 -8463 14573 -8403
rect 14173 -8473 14573 -8463
rect 14631 -8403 15031 -8293
rect 14631 -8463 14641 -8403
rect 14701 -8463 14961 -8403
rect 15021 -8463 15031 -8403
rect 14631 -8473 15031 -8463
rect 15087 -8403 15487 -8293
rect 15087 -8463 15097 -8403
rect 15157 -8463 15417 -8403
rect 15477 -8463 15487 -8403
rect 15087 -8473 15487 -8463
rect 66 -8537 80 -8473
rect 457 -8537 527 -8473
rect 913 -8537 983 -8473
rect 1371 -8537 1441 -8473
rect 1827 -8537 1897 -8473
rect 2283 -8537 2353 -8473
rect 2741 -8537 2811 -8473
rect 3197 -8537 3267 -8473
rect 3653 -8537 3723 -8473
rect 4111 -8537 4181 -8473
rect 4567 -8537 4637 -8473
rect 5023 -8537 5093 -8473
rect 5481 -8537 5551 -8473
rect 5937 -8537 6007 -8473
rect 6393 -8537 6463 -8473
rect 6851 -8537 6921 -8473
rect 66 -8547 400 -8537
rect 0 -8607 11 -8547
rect 71 -8607 331 -8547
rect 391 -8607 400 -8547
rect 0 -8897 14 -8607
rect 66 -8897 400 -8607
rect 0 -8957 11 -8897
rect 71 -8957 331 -8897
rect 391 -8957 400 -8897
rect 0 -9049 14 -8957
rect 66 -8967 400 -8957
rect 457 -8547 857 -8537
rect 457 -8607 467 -8547
rect 527 -8607 787 -8547
rect 847 -8607 857 -8547
rect 457 -8719 857 -8607
rect 913 -8547 1313 -8537
rect 913 -8607 923 -8547
rect 983 -8607 1243 -8547
rect 1303 -8607 1313 -8547
rect 913 -8719 1313 -8607
rect 1371 -8547 1771 -8537
rect 1371 -8607 1381 -8547
rect 1441 -8607 1701 -8547
rect 1761 -8607 1771 -8547
rect 1371 -8719 1771 -8607
rect 1827 -8547 2227 -8537
rect 1827 -8607 1837 -8547
rect 1897 -8607 2157 -8547
rect 2217 -8607 2227 -8547
rect 1827 -8719 2227 -8607
rect 2283 -8547 2683 -8537
rect 2283 -8607 2293 -8547
rect 2353 -8607 2613 -8547
rect 2673 -8607 2683 -8547
rect 2283 -8719 2683 -8607
rect 2741 -8547 3141 -8537
rect 2741 -8607 2751 -8547
rect 2811 -8607 3071 -8547
rect 3131 -8607 3141 -8547
rect 2741 -8719 3141 -8607
rect 3197 -8547 3597 -8537
rect 3197 -8607 3207 -8547
rect 3267 -8607 3527 -8547
rect 3587 -8607 3597 -8547
rect 3197 -8719 3597 -8607
rect 3653 -8547 4053 -8537
rect 3653 -8607 3663 -8547
rect 3723 -8607 3983 -8547
rect 4043 -8607 4053 -8547
rect 3653 -8719 4053 -8607
rect 457 -8789 4053 -8719
rect 457 -8897 857 -8789
rect 457 -8957 467 -8897
rect 527 -8957 787 -8897
rect 847 -8957 857 -8897
rect 457 -8967 857 -8957
rect 913 -8897 1313 -8789
rect 913 -8957 923 -8897
rect 983 -8957 1243 -8897
rect 1303 -8957 1313 -8897
rect 913 -8967 1313 -8957
rect 1371 -8897 1771 -8789
rect 1371 -8957 1381 -8897
rect 1441 -8957 1701 -8897
rect 1761 -8957 1771 -8897
rect 1371 -8967 1771 -8957
rect 1827 -8897 2227 -8789
rect 1827 -8957 1837 -8897
rect 1897 -8957 2157 -8897
rect 2217 -8957 2227 -8897
rect 1827 -8967 2227 -8957
rect 2283 -8897 2683 -8789
rect 2283 -8957 2293 -8897
rect 2353 -8957 2613 -8897
rect 2673 -8957 2683 -8897
rect 2283 -8967 2683 -8957
rect 2741 -8897 3141 -8789
rect 2741 -8957 2751 -8897
rect 2811 -8957 3071 -8897
rect 3131 -8957 3141 -8897
rect 2741 -8967 3141 -8957
rect 3197 -8897 3597 -8789
rect 3197 -8957 3207 -8897
rect 3267 -8957 3527 -8897
rect 3587 -8957 3597 -8897
rect 3197 -8967 3597 -8957
rect 3653 -8897 4053 -8789
rect 3653 -8957 3663 -8897
rect 3723 -8957 3983 -8897
rect 4043 -8957 4053 -8897
rect 3653 -8967 4053 -8957
rect 4111 -8547 4511 -8537
rect 4111 -8607 4121 -8547
rect 4181 -8607 4441 -8547
rect 4501 -8607 4511 -8547
rect 4111 -8719 4511 -8607
rect 4567 -8547 4967 -8537
rect 4567 -8607 4577 -8547
rect 4637 -8607 4897 -8547
rect 4957 -8607 4967 -8547
rect 4567 -8719 4967 -8607
rect 5023 -8547 5423 -8537
rect 5023 -8607 5033 -8547
rect 5093 -8607 5353 -8547
rect 5413 -8607 5423 -8547
rect 5023 -8719 5423 -8607
rect 5481 -8547 5881 -8537
rect 5481 -8607 5491 -8547
rect 5551 -8607 5811 -8547
rect 5871 -8607 5881 -8547
rect 5481 -8719 5881 -8607
rect 5937 -8547 6337 -8537
rect 5937 -8607 5947 -8547
rect 6007 -8607 6267 -8547
rect 6327 -8607 6337 -8547
rect 5937 -8719 6337 -8607
rect 6393 -8547 6793 -8537
rect 6393 -8607 6403 -8547
rect 6463 -8607 6723 -8547
rect 6783 -8607 6793 -8547
rect 6393 -8719 6793 -8607
rect 6851 -8547 7251 -8537
rect 6851 -8607 6861 -8547
rect 6921 -8607 7181 -8547
rect 7241 -8607 7251 -8547
rect 6851 -8719 7251 -8607
rect 4111 -8789 7251 -8719
rect 4111 -8897 4511 -8789
rect 4111 -8957 4121 -8897
rect 4181 -8957 4441 -8897
rect 4501 -8957 4511 -8897
rect 4111 -8967 4511 -8957
rect 4567 -8897 4967 -8789
rect 4567 -8957 4577 -8897
rect 4637 -8957 4897 -8897
rect 4957 -8957 4967 -8897
rect 4567 -8967 4967 -8957
rect 5023 -8897 5423 -8789
rect 5023 -8957 5033 -8897
rect 5093 -8957 5353 -8897
rect 5413 -8957 5423 -8897
rect 5023 -8967 5423 -8957
rect 5481 -8897 5881 -8789
rect 5481 -8957 5491 -8897
rect 5551 -8957 5811 -8897
rect 5871 -8957 5881 -8897
rect 5481 -8967 5881 -8957
rect 5937 -8897 6337 -8789
rect 5937 -8957 5947 -8897
rect 6007 -8957 6267 -8897
rect 6327 -8957 6337 -8897
rect 5937 -8967 6337 -8957
rect 6393 -8897 6793 -8789
rect 6393 -8957 6403 -8897
rect 6463 -8957 6723 -8897
rect 6783 -8957 6793 -8897
rect 6393 -8967 6793 -8957
rect 6851 -8897 7251 -8789
rect 6851 -8957 6861 -8897
rect 6921 -8957 7181 -8897
rect 7241 -8957 7251 -8897
rect 6851 -8967 7251 -8957
rect 7307 -8547 7707 -8537
rect 7307 -8607 7317 -8547
rect 7377 -8607 7637 -8547
rect 7697 -8607 7707 -8547
rect 7307 -8719 7707 -8607
rect 7763 -8547 8163 -8537
rect 7763 -8607 7773 -8547
rect 7833 -8607 8093 -8547
rect 8153 -8607 8163 -8547
rect 7763 -8719 8163 -8607
rect 8237 -8547 8637 -8537
rect 8237 -8607 8247 -8547
rect 8307 -8607 8567 -8547
rect 8627 -8607 8637 -8547
rect 8237 -8719 8637 -8607
rect 8693 -8547 9093 -8537
rect 8693 -8607 8703 -8547
rect 8763 -8607 9023 -8547
rect 9083 -8607 9093 -8547
rect 8693 -8719 9093 -8607
rect 9151 -8547 9551 -8537
rect 9151 -8607 9161 -8547
rect 9221 -8607 9481 -8547
rect 9541 -8607 9551 -8547
rect 9151 -8719 9551 -8607
rect 9607 -8547 10007 -8537
rect 9607 -8607 9617 -8547
rect 9677 -8607 9937 -8547
rect 9997 -8607 10007 -8547
rect 9607 -8719 10007 -8607
rect 10063 -8547 10463 -8537
rect 10063 -8607 10073 -8547
rect 10133 -8607 10393 -8547
rect 10453 -8607 10463 -8547
rect 10063 -8719 10463 -8607
rect 10521 -8547 10921 -8537
rect 10521 -8607 10531 -8547
rect 10591 -8607 10851 -8547
rect 10911 -8607 10921 -8547
rect 10521 -8719 10921 -8607
rect 10977 -8547 11377 -8537
rect 10977 -8607 10987 -8547
rect 11047 -8607 11307 -8547
rect 11367 -8607 11377 -8547
rect 10977 -8719 11377 -8607
rect 11433 -8547 11833 -8537
rect 11433 -8607 11443 -8547
rect 11503 -8607 11763 -8547
rect 11823 -8607 11833 -8547
rect 11433 -8719 11833 -8607
rect 11891 -8547 12291 -8537
rect 11891 -8607 11901 -8547
rect 11961 -8607 12221 -8547
rect 12281 -8607 12291 -8547
rect 11891 -8719 12291 -8607
rect 12347 -8547 12747 -8537
rect 12347 -8607 12357 -8547
rect 12417 -8607 12677 -8547
rect 12737 -8607 12747 -8547
rect 12347 -8719 12747 -8607
rect 12803 -8547 13203 -8537
rect 12803 -8607 12813 -8547
rect 12873 -8607 13133 -8547
rect 13193 -8607 13203 -8547
rect 12803 -8719 13203 -8607
rect 13261 -8547 13661 -8537
rect 13261 -8607 13271 -8547
rect 13331 -8607 13591 -8547
rect 13651 -8607 13661 -8547
rect 13261 -8719 13661 -8607
rect 13717 -8547 14117 -8537
rect 13717 -8607 13727 -8547
rect 13787 -8607 14047 -8547
rect 14107 -8607 14117 -8547
rect 13717 -8719 14117 -8607
rect 14173 -8547 14573 -8537
rect 14173 -8607 14183 -8547
rect 14243 -8607 14503 -8547
rect 14563 -8607 14573 -8547
rect 14173 -8719 14573 -8607
rect 14631 -8547 15031 -8537
rect 14631 -8607 14641 -8547
rect 14701 -8607 14961 -8547
rect 15021 -8607 15031 -8547
rect 14631 -8719 15031 -8607
rect 15087 -8547 15487 -8537
rect 15087 -8607 15097 -8547
rect 15157 -8607 15417 -8547
rect 15477 -8607 15487 -8547
rect 15087 -8719 15487 -8607
rect 7307 -8789 15487 -8719
rect 7307 -8897 7707 -8789
rect 7307 -8957 7317 -8897
rect 7377 -8957 7637 -8897
rect 7697 -8957 7707 -8897
rect 7307 -8967 7707 -8957
rect 7763 -8897 8163 -8789
rect 7763 -8957 7773 -8897
rect 7833 -8957 8093 -8897
rect 8153 -8957 8163 -8897
rect 7763 -8967 8163 -8957
rect 8237 -8897 8637 -8789
rect 8237 -8957 8247 -8897
rect 8307 -8957 8567 -8897
rect 8627 -8957 8637 -8897
rect 8237 -8967 8637 -8957
rect 8693 -8897 9093 -8789
rect 8693 -8957 8703 -8897
rect 8763 -8957 9023 -8897
rect 9083 -8957 9093 -8897
rect 8693 -8967 9093 -8957
rect 9151 -8897 9551 -8789
rect 9151 -8957 9161 -8897
rect 9221 -8957 9481 -8897
rect 9541 -8957 9551 -8897
rect 9151 -8967 9551 -8957
rect 9607 -8897 10007 -8789
rect 9607 -8957 9617 -8897
rect 9677 -8957 9937 -8897
rect 9997 -8957 10007 -8897
rect 9607 -8967 10007 -8957
rect 10063 -8897 10463 -8789
rect 10063 -8957 10073 -8897
rect 10133 -8957 10393 -8897
rect 10453 -8957 10463 -8897
rect 10063 -8967 10463 -8957
rect 10521 -8897 10921 -8789
rect 10521 -8957 10531 -8897
rect 10591 -8957 10851 -8897
rect 10911 -8957 10921 -8897
rect 10521 -8967 10921 -8957
rect 10977 -8897 11377 -8789
rect 10977 -8957 10987 -8897
rect 11047 -8957 11307 -8897
rect 11367 -8957 11377 -8897
rect 10977 -8967 11377 -8957
rect 11433 -8897 11833 -8789
rect 11433 -8957 11443 -8897
rect 11503 -8957 11763 -8897
rect 11823 -8957 11833 -8897
rect 11433 -8967 11833 -8957
rect 11891 -8897 12291 -8789
rect 11891 -8957 11901 -8897
rect 11961 -8957 12221 -8897
rect 12281 -8957 12291 -8897
rect 11891 -8967 12291 -8957
rect 12347 -8897 12747 -8789
rect 12347 -8957 12357 -8897
rect 12417 -8957 12677 -8897
rect 12737 -8957 12747 -8897
rect 12347 -8967 12747 -8957
rect 12803 -8897 13203 -8789
rect 12803 -8957 12813 -8897
rect 12873 -8957 13133 -8897
rect 13193 -8957 13203 -8897
rect 12803 -8967 13203 -8957
rect 13261 -8897 13661 -8789
rect 13261 -8957 13271 -8897
rect 13331 -8957 13591 -8897
rect 13651 -8957 13661 -8897
rect 13261 -8967 13661 -8957
rect 13717 -8897 14117 -8789
rect 13717 -8957 13727 -8897
rect 13787 -8957 14047 -8897
rect 14107 -8957 14117 -8897
rect 13717 -8967 14117 -8957
rect 14173 -8897 14573 -8789
rect 14173 -8957 14183 -8897
rect 14243 -8957 14503 -8897
rect 14563 -8957 14573 -8897
rect 14173 -8967 14573 -8957
rect 14631 -8897 15031 -8789
rect 14631 -8957 14641 -8897
rect 14701 -8957 14961 -8897
rect 15021 -8957 15031 -8897
rect 14631 -8967 15031 -8957
rect 15087 -8897 15487 -8789
rect 15087 -8957 15097 -8897
rect 15157 -8957 15417 -8897
rect 15477 -8957 15487 -8897
rect 15087 -8967 15487 -8957
rect 66 -9039 80 -8967
rect 457 -9039 527 -8967
rect 913 -9039 984 -8967
rect 1371 -9039 1442 -8967
rect 1827 -9039 1898 -8967
rect 2283 -9039 2354 -8967
rect 2741 -9039 2812 -8967
rect 3197 -9039 3268 -8967
rect 3653 -9039 3724 -8967
rect 4111 -9039 4182 -8967
rect 4567 -9039 4638 -8967
rect 5023 -9039 5094 -8967
rect 5481 -9039 5552 -8967
rect 5937 -9039 6008 -8967
rect 6393 -9039 6464 -8967
rect 6851 -9039 6922 -8967
rect 7307 -9039 7378 -8967
rect 7763 -9039 7834 -8967
rect 8237 -9039 8308 -8967
rect 8693 -9039 8764 -8967
rect 9151 -9039 9222 -8967
rect 9607 -9039 9678 -8967
rect 10063 -9039 10134 -8967
rect 10521 -9039 10592 -8967
rect 10977 -9039 11048 -8967
rect 11433 -9039 11504 -8967
rect 11891 -9039 11962 -8967
rect 12347 -9039 12418 -8967
rect 12803 -9039 12874 -8967
rect 13261 -9039 13332 -8967
rect 13717 -9039 13788 -8967
rect 14173 -9039 14244 -8967
rect 14631 -9039 14702 -8967
rect 66 -9049 400 -9039
rect 0 -9109 11 -9049
rect 71 -9109 331 -9049
rect 391 -9109 400 -9049
rect 0 -9399 14 -9109
rect 66 -9399 400 -9109
rect 0 -9459 11 -9399
rect 71 -9459 331 -9399
rect 391 -9459 400 -9399
rect 0 -9541 14 -9459
rect 66 -9469 400 -9459
rect 457 -9049 857 -9039
rect 457 -9109 467 -9049
rect 527 -9109 787 -9049
rect 847 -9109 857 -9049
rect 457 -9219 857 -9109
rect 913 -9049 1313 -9039
rect 913 -9109 923 -9049
rect 983 -9109 1243 -9049
rect 1303 -9109 1313 -9049
rect 913 -9219 1313 -9109
rect 1371 -9049 1771 -9039
rect 1371 -9109 1381 -9049
rect 1441 -9109 1701 -9049
rect 1761 -9109 1771 -9049
rect 1371 -9219 1771 -9109
rect 1827 -9049 2227 -9039
rect 1827 -9109 1837 -9049
rect 1897 -9109 2157 -9049
rect 2217 -9109 2227 -9049
rect 1827 -9219 2227 -9109
rect 2283 -9049 2683 -9039
rect 2283 -9109 2293 -9049
rect 2353 -9109 2613 -9049
rect 2673 -9109 2683 -9049
rect 2283 -9219 2683 -9109
rect 2741 -9049 3141 -9039
rect 2741 -9109 2751 -9049
rect 2811 -9109 3071 -9049
rect 3131 -9109 3141 -9049
rect 2741 -9219 3141 -9109
rect 3197 -9049 3597 -9039
rect 3197 -9109 3207 -9049
rect 3267 -9109 3527 -9049
rect 3587 -9109 3597 -9049
rect 3197 -9219 3597 -9109
rect 3653 -9049 4053 -9039
rect 3653 -9109 3663 -9049
rect 3723 -9109 3983 -9049
rect 4043 -9109 4053 -9049
rect 3653 -9219 4053 -9109
rect 457 -9289 4053 -9219
rect 457 -9399 857 -9289
rect 457 -9459 467 -9399
rect 527 -9459 787 -9399
rect 847 -9459 857 -9399
rect 457 -9469 857 -9459
rect 913 -9399 1313 -9289
rect 913 -9459 923 -9399
rect 983 -9459 1243 -9399
rect 1303 -9459 1313 -9399
rect 913 -9469 1313 -9459
rect 1371 -9399 1771 -9289
rect 1371 -9459 1381 -9399
rect 1441 -9459 1701 -9399
rect 1761 -9459 1771 -9399
rect 1371 -9469 1771 -9459
rect 1827 -9399 2227 -9289
rect 1827 -9459 1837 -9399
rect 1897 -9459 2157 -9399
rect 2217 -9459 2227 -9399
rect 1827 -9469 2227 -9459
rect 2283 -9399 2683 -9289
rect 2283 -9459 2293 -9399
rect 2353 -9459 2613 -9399
rect 2673 -9459 2683 -9399
rect 2283 -9469 2683 -9459
rect 2741 -9399 3141 -9289
rect 2741 -9459 2751 -9399
rect 2811 -9459 3071 -9399
rect 3131 -9459 3141 -9399
rect 2741 -9469 3141 -9459
rect 3197 -9399 3597 -9289
rect 3197 -9459 3207 -9399
rect 3267 -9459 3527 -9399
rect 3587 -9459 3597 -9399
rect 3197 -9469 3597 -9459
rect 3653 -9399 4053 -9289
rect 3653 -9459 3663 -9399
rect 3723 -9459 3983 -9399
rect 4043 -9459 4053 -9399
rect 3653 -9469 4053 -9459
rect 4111 -9049 4511 -9039
rect 4111 -9109 4121 -9049
rect 4181 -9109 4441 -9049
rect 4501 -9109 4511 -9049
rect 4111 -9219 4511 -9109
rect 4567 -9049 4967 -9039
rect 4567 -9109 4577 -9049
rect 4637 -9109 4897 -9049
rect 4957 -9109 4967 -9049
rect 4567 -9219 4967 -9109
rect 5023 -9049 5423 -9039
rect 5023 -9109 5033 -9049
rect 5093 -9109 5353 -9049
rect 5413 -9109 5423 -9049
rect 5023 -9219 5423 -9109
rect 5481 -9049 5881 -9039
rect 5481 -9109 5491 -9049
rect 5551 -9109 5811 -9049
rect 5871 -9109 5881 -9049
rect 5481 -9219 5881 -9109
rect 5937 -9049 6337 -9039
rect 5937 -9109 5947 -9049
rect 6007 -9109 6267 -9049
rect 6327 -9109 6337 -9049
rect 5937 -9219 6337 -9109
rect 6393 -9049 6793 -9039
rect 6393 -9109 6403 -9049
rect 6463 -9109 6723 -9049
rect 6783 -9109 6793 -9049
rect 6393 -9219 6793 -9109
rect 6851 -9049 7251 -9039
rect 6851 -9109 6861 -9049
rect 6921 -9109 7181 -9049
rect 7241 -9109 7251 -9049
rect 6851 -9219 7251 -9109
rect 4111 -9289 7251 -9219
rect 4111 -9399 4511 -9289
rect 4111 -9459 4121 -9399
rect 4181 -9459 4441 -9399
rect 4501 -9459 4511 -9399
rect 4111 -9469 4511 -9459
rect 4567 -9399 4967 -9289
rect 4567 -9459 4577 -9399
rect 4637 -9459 4897 -9399
rect 4957 -9459 4967 -9399
rect 4567 -9469 4967 -9459
rect 5023 -9399 5423 -9289
rect 5023 -9459 5033 -9399
rect 5093 -9459 5353 -9399
rect 5413 -9459 5423 -9399
rect 5023 -9469 5423 -9459
rect 5481 -9399 5881 -9289
rect 5481 -9459 5491 -9399
rect 5551 -9459 5811 -9399
rect 5871 -9459 5881 -9399
rect 5481 -9469 5881 -9459
rect 5937 -9399 6337 -9289
rect 5937 -9459 5947 -9399
rect 6007 -9459 6267 -9399
rect 6327 -9459 6337 -9399
rect 5937 -9469 6337 -9459
rect 6393 -9399 6793 -9289
rect 6393 -9459 6403 -9399
rect 6463 -9459 6723 -9399
rect 6783 -9459 6793 -9399
rect 6393 -9469 6793 -9459
rect 6851 -9399 7251 -9289
rect 6851 -9459 6861 -9399
rect 6921 -9459 7181 -9399
rect 7241 -9459 7251 -9399
rect 6851 -9469 7251 -9459
rect 7307 -9049 7707 -9039
rect 7307 -9109 7317 -9049
rect 7377 -9109 7637 -9049
rect 7697 -9109 7707 -9049
rect 7307 -9219 7707 -9109
rect 7763 -9049 8163 -9039
rect 7763 -9109 7773 -9049
rect 7833 -9109 8093 -9049
rect 8153 -9109 8163 -9049
rect 7763 -9219 8163 -9109
rect 8237 -9049 8637 -9039
rect 8237 -9109 8247 -9049
rect 8307 -9109 8567 -9049
rect 8627 -9109 8637 -9049
rect 8237 -9219 8637 -9109
rect 8693 -9049 9093 -9039
rect 8693 -9109 8703 -9049
rect 8763 -9109 9023 -9049
rect 9083 -9109 9093 -9049
rect 8693 -9219 9093 -9109
rect 9151 -9049 9551 -9039
rect 9151 -9109 9161 -9049
rect 9221 -9109 9481 -9049
rect 9541 -9109 9551 -9049
rect 9151 -9219 9551 -9109
rect 9607 -9049 10007 -9039
rect 9607 -9109 9617 -9049
rect 9677 -9109 9937 -9049
rect 9997 -9109 10007 -9049
rect 9607 -9219 10007 -9109
rect 10063 -9049 10463 -9039
rect 10063 -9109 10073 -9049
rect 10133 -9109 10393 -9049
rect 10453 -9109 10463 -9049
rect 10063 -9219 10463 -9109
rect 10521 -9049 10921 -9039
rect 10521 -9109 10531 -9049
rect 10591 -9109 10851 -9049
rect 10911 -9109 10921 -9049
rect 10521 -9219 10921 -9109
rect 10977 -9049 11377 -9039
rect 10977 -9109 10987 -9049
rect 11047 -9109 11307 -9049
rect 11367 -9109 11377 -9049
rect 10977 -9219 11377 -9109
rect 11433 -9049 11833 -9039
rect 11433 -9109 11443 -9049
rect 11503 -9109 11763 -9049
rect 11823 -9109 11833 -9049
rect 11433 -9219 11833 -9109
rect 11891 -9049 12291 -9039
rect 11891 -9109 11901 -9049
rect 11961 -9109 12221 -9049
rect 12281 -9109 12291 -9049
rect 11891 -9219 12291 -9109
rect 12347 -9049 12747 -9039
rect 12347 -9109 12357 -9049
rect 12417 -9109 12677 -9049
rect 12737 -9109 12747 -9049
rect 12347 -9219 12747 -9109
rect 12803 -9049 13203 -9039
rect 12803 -9109 12813 -9049
rect 12873 -9109 13133 -9049
rect 13193 -9109 13203 -9049
rect 12803 -9219 13203 -9109
rect 13261 -9049 13661 -9039
rect 13261 -9109 13271 -9049
rect 13331 -9109 13591 -9049
rect 13651 -9109 13661 -9049
rect 13261 -9219 13661 -9109
rect 13717 -9049 14117 -9039
rect 13717 -9109 13727 -9049
rect 13787 -9109 14047 -9049
rect 14107 -9109 14117 -9049
rect 13717 -9219 14117 -9109
rect 14173 -9049 14573 -9039
rect 14173 -9109 14183 -9049
rect 14243 -9109 14503 -9049
rect 14563 -9109 14573 -9049
rect 14173 -9219 14573 -9109
rect 14631 -9049 15031 -9039
rect 14631 -9109 14641 -9049
rect 14701 -9109 14961 -9049
rect 15021 -9109 15031 -9049
rect 14631 -9219 15031 -9109
rect 15087 -9049 15487 -9039
rect 15087 -9109 15097 -9049
rect 15157 -9109 15417 -9049
rect 15477 -9109 15487 -9049
rect 15087 -9219 15487 -9109
rect 7307 -9289 15487 -9219
rect 7307 -9399 7707 -9289
rect 7307 -9459 7317 -9399
rect 7377 -9459 7637 -9399
rect 7697 -9459 7707 -9399
rect 7307 -9469 7707 -9459
rect 7763 -9399 8163 -9289
rect 7763 -9459 7773 -9399
rect 7833 -9459 8093 -9399
rect 8153 -9459 8163 -9399
rect 7763 -9469 8163 -9459
rect 8237 -9399 8637 -9289
rect 8237 -9459 8247 -9399
rect 8307 -9459 8567 -9399
rect 8627 -9459 8637 -9399
rect 8237 -9469 8637 -9459
rect 8693 -9399 9093 -9289
rect 8693 -9459 8703 -9399
rect 8763 -9459 9023 -9399
rect 9083 -9459 9093 -9399
rect 8693 -9469 9093 -9459
rect 9151 -9399 9551 -9289
rect 9151 -9459 9161 -9399
rect 9221 -9459 9481 -9399
rect 9541 -9459 9551 -9399
rect 9151 -9469 9551 -9459
rect 9607 -9399 10007 -9289
rect 9607 -9459 9617 -9399
rect 9677 -9459 9937 -9399
rect 9997 -9459 10007 -9399
rect 9607 -9469 10007 -9459
rect 10063 -9399 10463 -9289
rect 10063 -9459 10073 -9399
rect 10133 -9459 10393 -9399
rect 10453 -9459 10463 -9399
rect 10063 -9469 10463 -9459
rect 10521 -9399 10921 -9289
rect 10521 -9459 10531 -9399
rect 10591 -9459 10851 -9399
rect 10911 -9459 10921 -9399
rect 10521 -9469 10921 -9459
rect 10977 -9399 11377 -9289
rect 10977 -9459 10987 -9399
rect 11047 -9459 11307 -9399
rect 11367 -9459 11377 -9399
rect 10977 -9469 11377 -9459
rect 11433 -9399 11833 -9289
rect 11433 -9459 11443 -9399
rect 11503 -9459 11763 -9399
rect 11823 -9459 11833 -9399
rect 11433 -9469 11833 -9459
rect 11891 -9399 12291 -9289
rect 11891 -9459 11901 -9399
rect 11961 -9459 12221 -9399
rect 12281 -9459 12291 -9399
rect 11891 -9469 12291 -9459
rect 12347 -9399 12747 -9289
rect 12347 -9459 12357 -9399
rect 12417 -9459 12677 -9399
rect 12737 -9459 12747 -9399
rect 12347 -9469 12747 -9459
rect 12803 -9399 13203 -9289
rect 12803 -9459 12813 -9399
rect 12873 -9459 13133 -9399
rect 13193 -9459 13203 -9399
rect 12803 -9469 13203 -9459
rect 13261 -9399 13661 -9289
rect 13261 -9459 13271 -9399
rect 13331 -9459 13591 -9399
rect 13651 -9459 13661 -9399
rect 13261 -9469 13661 -9459
rect 13717 -9399 14117 -9289
rect 13717 -9459 13727 -9399
rect 13787 -9459 14047 -9399
rect 14107 -9459 14117 -9399
rect 13717 -9469 14117 -9459
rect 14173 -9399 14573 -9289
rect 14173 -9459 14183 -9399
rect 14243 -9459 14503 -9399
rect 14563 -9459 14573 -9399
rect 14173 -9469 14573 -9459
rect 14631 -9399 15031 -9289
rect 14631 -9459 14641 -9399
rect 14701 -9459 14961 -9399
rect 15021 -9459 15031 -9399
rect 14631 -9469 15031 -9459
rect 15087 -9399 15487 -9289
rect 15087 -9459 15097 -9399
rect 15157 -9459 15417 -9399
rect 15477 -9459 15487 -9399
rect 15087 -9469 15487 -9459
rect 66 -9531 80 -9469
rect 457 -9531 528 -9469
rect 913 -9531 984 -9469
rect 1371 -9531 1442 -9469
rect 1827 -9531 1898 -9469
rect 2283 -9531 2354 -9469
rect 2741 -9531 2811 -9469
rect 3197 -9531 3267 -9469
rect 3653 -9531 3723 -9469
rect 4111 -9531 4181 -9469
rect 4567 -9531 4637 -9469
rect 5023 -9531 5093 -9469
rect 5481 -9531 5551 -9469
rect 5937 -9531 6007 -9469
rect 6393 -9531 6463 -9469
rect 6851 -9531 6921 -9469
rect 7307 -9531 7377 -9469
rect 7763 -9531 7833 -9469
rect 8237 -9531 8307 -9469
rect 8693 -9531 8763 -9469
rect 9151 -9531 9221 -9469
rect 9607 -9531 9677 -9469
rect 10063 -9531 10133 -9469
rect 10521 -9531 10591 -9469
rect 10977 -9531 11047 -9469
rect 11433 -9531 11503 -9469
rect 11891 -9531 11961 -9469
rect 12347 -9531 12417 -9469
rect 12803 -9531 12873 -9469
rect 13261 -9531 13331 -9469
rect 13717 -9531 13787 -9469
rect 14173 -9531 14243 -9469
rect 14631 -9531 14701 -9469
rect 66 -9541 400 -9531
rect 0 -9601 11 -9541
rect 71 -9601 331 -9541
rect 391 -9601 400 -9541
rect 0 -9891 14 -9601
rect 66 -9891 400 -9601
rect 0 -9951 11 -9891
rect 71 -9951 331 -9891
rect 391 -9951 400 -9891
rect 0 -10057 14 -9951
rect 66 -9961 400 -9951
rect 457 -9541 857 -9531
rect 457 -9601 467 -9541
rect 527 -9601 787 -9541
rect 847 -9601 857 -9541
rect 457 -9711 857 -9601
rect 913 -9541 1313 -9531
rect 913 -9601 923 -9541
rect 983 -9601 1243 -9541
rect 1303 -9601 1313 -9541
rect 913 -9711 1313 -9601
rect 1371 -9541 1771 -9531
rect 1371 -9601 1381 -9541
rect 1441 -9601 1701 -9541
rect 1761 -9601 1771 -9541
rect 1371 -9711 1771 -9601
rect 1827 -9541 2227 -9531
rect 1827 -9601 1837 -9541
rect 1897 -9601 2157 -9541
rect 2217 -9601 2227 -9541
rect 1827 -9711 2227 -9601
rect 2283 -9541 2683 -9531
rect 2283 -9601 2293 -9541
rect 2353 -9601 2613 -9541
rect 2673 -9601 2683 -9541
rect 2283 -9711 2683 -9601
rect 2741 -9541 3141 -9531
rect 2741 -9601 2751 -9541
rect 2811 -9601 3071 -9541
rect 3131 -9601 3141 -9541
rect 2741 -9711 3141 -9601
rect 3197 -9541 3597 -9531
rect 3197 -9601 3207 -9541
rect 3267 -9601 3527 -9541
rect 3587 -9601 3597 -9541
rect 3197 -9711 3597 -9601
rect 3653 -9541 4053 -9531
rect 3653 -9601 3663 -9541
rect 3723 -9601 3983 -9541
rect 4043 -9601 4053 -9541
rect 3653 -9711 4053 -9601
rect 457 -9781 4053 -9711
rect 457 -9891 857 -9781
rect 457 -9951 467 -9891
rect 527 -9951 787 -9891
rect 847 -9951 857 -9891
rect 457 -9961 857 -9951
rect 913 -9891 1313 -9781
rect 913 -9951 923 -9891
rect 983 -9951 1243 -9891
rect 1303 -9951 1313 -9891
rect 913 -9961 1313 -9951
rect 1371 -9891 1771 -9781
rect 1371 -9951 1381 -9891
rect 1441 -9951 1701 -9891
rect 1761 -9951 1771 -9891
rect 1371 -9961 1771 -9951
rect 1827 -9891 2227 -9781
rect 1827 -9951 1837 -9891
rect 1897 -9951 2157 -9891
rect 2217 -9951 2227 -9891
rect 1827 -9961 2227 -9951
rect 2283 -9891 2683 -9781
rect 2283 -9951 2293 -9891
rect 2353 -9951 2613 -9891
rect 2673 -9951 2683 -9891
rect 2283 -9961 2683 -9951
rect 2741 -9891 3141 -9781
rect 2741 -9951 2751 -9891
rect 2811 -9951 3071 -9891
rect 3131 -9951 3141 -9891
rect 2741 -9961 3141 -9951
rect 3197 -9891 3597 -9781
rect 3197 -9951 3207 -9891
rect 3267 -9951 3527 -9891
rect 3587 -9951 3597 -9891
rect 3197 -9961 3597 -9951
rect 3653 -9891 4053 -9781
rect 3653 -9951 3663 -9891
rect 3723 -9951 3983 -9891
rect 4043 -9951 4053 -9891
rect 3653 -9961 4053 -9951
rect 4111 -9541 4511 -9531
rect 4111 -9601 4121 -9541
rect 4181 -9601 4441 -9541
rect 4501 -9601 4511 -9541
rect 4111 -9711 4511 -9601
rect 4567 -9541 4967 -9531
rect 4567 -9601 4577 -9541
rect 4637 -9601 4897 -9541
rect 4957 -9601 4967 -9541
rect 4567 -9711 4967 -9601
rect 5023 -9541 5423 -9531
rect 5023 -9601 5033 -9541
rect 5093 -9601 5353 -9541
rect 5413 -9601 5423 -9541
rect 5023 -9711 5423 -9601
rect 5481 -9541 5881 -9531
rect 5481 -9601 5491 -9541
rect 5551 -9601 5811 -9541
rect 5871 -9601 5881 -9541
rect 5481 -9711 5881 -9601
rect 5937 -9541 6337 -9531
rect 5937 -9601 5947 -9541
rect 6007 -9601 6267 -9541
rect 6327 -9601 6337 -9541
rect 5937 -9711 6337 -9601
rect 6393 -9541 6793 -9531
rect 6393 -9601 6403 -9541
rect 6463 -9601 6723 -9541
rect 6783 -9601 6793 -9541
rect 6393 -9711 6793 -9601
rect 6851 -9541 7251 -9531
rect 6851 -9601 6861 -9541
rect 6921 -9601 7181 -9541
rect 7241 -9601 7251 -9541
rect 6851 -9711 7251 -9601
rect 4111 -9781 7251 -9711
rect 4111 -9891 4511 -9781
rect 4111 -9951 4121 -9891
rect 4181 -9951 4441 -9891
rect 4501 -9951 4511 -9891
rect 4111 -9961 4511 -9951
rect 4567 -9891 4967 -9781
rect 4567 -9951 4577 -9891
rect 4637 -9951 4897 -9891
rect 4957 -9951 4967 -9891
rect 4567 -9961 4967 -9951
rect 5023 -9891 5423 -9781
rect 5023 -9951 5033 -9891
rect 5093 -9951 5353 -9891
rect 5413 -9951 5423 -9891
rect 5023 -9961 5423 -9951
rect 5481 -9891 5881 -9781
rect 5481 -9951 5491 -9891
rect 5551 -9951 5811 -9891
rect 5871 -9951 5881 -9891
rect 5481 -9961 5881 -9951
rect 5937 -9891 6337 -9781
rect 5937 -9951 5947 -9891
rect 6007 -9951 6267 -9891
rect 6327 -9951 6337 -9891
rect 5937 -9961 6337 -9951
rect 6393 -9891 6793 -9781
rect 6393 -9951 6403 -9891
rect 6463 -9951 6723 -9891
rect 6783 -9951 6793 -9891
rect 6393 -9961 6793 -9951
rect 6851 -9891 7251 -9781
rect 6851 -9951 6861 -9891
rect 6921 -9951 7181 -9891
rect 7241 -9951 7251 -9891
rect 6851 -9961 7251 -9951
rect 7307 -9541 7707 -9531
rect 7307 -9601 7317 -9541
rect 7377 -9601 7637 -9541
rect 7697 -9601 7707 -9541
rect 7307 -9711 7707 -9601
rect 7763 -9541 8163 -9531
rect 7763 -9601 7773 -9541
rect 7833 -9601 8093 -9541
rect 8153 -9601 8163 -9541
rect 7763 -9711 8163 -9601
rect 8237 -9541 8637 -9531
rect 8237 -9601 8247 -9541
rect 8307 -9601 8567 -9541
rect 8627 -9601 8637 -9541
rect 8237 -9711 8637 -9601
rect 8693 -9541 9093 -9531
rect 8693 -9601 8703 -9541
rect 8763 -9601 9023 -9541
rect 9083 -9601 9093 -9541
rect 8693 -9711 9093 -9601
rect 9151 -9541 9551 -9531
rect 9151 -9601 9161 -9541
rect 9221 -9601 9481 -9541
rect 9541 -9601 9551 -9541
rect 9151 -9711 9551 -9601
rect 9607 -9541 10007 -9531
rect 9607 -9601 9617 -9541
rect 9677 -9601 9937 -9541
rect 9997 -9601 10007 -9541
rect 9607 -9711 10007 -9601
rect 10063 -9541 10463 -9531
rect 10063 -9601 10073 -9541
rect 10133 -9601 10393 -9541
rect 10453 -9601 10463 -9541
rect 10063 -9711 10463 -9601
rect 10521 -9541 10921 -9531
rect 10521 -9601 10531 -9541
rect 10591 -9601 10851 -9541
rect 10911 -9601 10921 -9541
rect 10521 -9711 10921 -9601
rect 10977 -9541 11377 -9531
rect 10977 -9601 10987 -9541
rect 11047 -9601 11307 -9541
rect 11367 -9601 11377 -9541
rect 10977 -9711 11377 -9601
rect 11433 -9541 11833 -9531
rect 11433 -9601 11443 -9541
rect 11503 -9601 11763 -9541
rect 11823 -9601 11833 -9541
rect 11433 -9711 11833 -9601
rect 11891 -9541 12291 -9531
rect 11891 -9601 11901 -9541
rect 11961 -9601 12221 -9541
rect 12281 -9601 12291 -9541
rect 11891 -9711 12291 -9601
rect 12347 -9541 12747 -9531
rect 12347 -9601 12357 -9541
rect 12417 -9601 12677 -9541
rect 12737 -9601 12747 -9541
rect 12347 -9711 12747 -9601
rect 12803 -9541 13203 -9531
rect 12803 -9601 12813 -9541
rect 12873 -9601 13133 -9541
rect 13193 -9601 13203 -9541
rect 12803 -9711 13203 -9601
rect 13261 -9541 13661 -9531
rect 13261 -9601 13271 -9541
rect 13331 -9601 13591 -9541
rect 13651 -9601 13661 -9541
rect 13261 -9711 13661 -9601
rect 13717 -9541 14117 -9531
rect 13717 -9601 13727 -9541
rect 13787 -9601 14047 -9541
rect 14107 -9601 14117 -9541
rect 13717 -9711 14117 -9601
rect 14173 -9541 14573 -9531
rect 14173 -9601 14183 -9541
rect 14243 -9601 14503 -9541
rect 14563 -9601 14573 -9541
rect 14173 -9711 14573 -9601
rect 14631 -9541 15031 -9531
rect 14631 -9601 14641 -9541
rect 14701 -9601 14961 -9541
rect 15021 -9601 15031 -9541
rect 14631 -9711 15031 -9601
rect 15087 -9541 15487 -9531
rect 15087 -9601 15097 -9541
rect 15157 -9601 15417 -9541
rect 15477 -9601 15487 -9541
rect 15087 -9711 15487 -9601
rect 7307 -9781 15487 -9711
rect 7307 -9891 7707 -9781
rect 7307 -9951 7317 -9891
rect 7377 -9951 7637 -9891
rect 7697 -9951 7707 -9891
rect 7307 -9961 7707 -9951
rect 7763 -9891 8163 -9781
rect 7763 -9951 7773 -9891
rect 7833 -9951 8093 -9891
rect 8153 -9951 8163 -9891
rect 7763 -9961 8163 -9951
rect 8237 -9891 8637 -9781
rect 8237 -9951 8247 -9891
rect 8307 -9951 8567 -9891
rect 8627 -9951 8637 -9891
rect 8237 -9961 8637 -9951
rect 8693 -9891 9093 -9781
rect 8693 -9951 8703 -9891
rect 8763 -9951 9023 -9891
rect 9083 -9951 9093 -9891
rect 8693 -9961 9093 -9951
rect 9151 -9891 9551 -9781
rect 9151 -9951 9161 -9891
rect 9221 -9951 9481 -9891
rect 9541 -9951 9551 -9891
rect 9151 -9961 9551 -9951
rect 9607 -9891 10007 -9781
rect 9607 -9951 9617 -9891
rect 9677 -9951 9937 -9891
rect 9997 -9951 10007 -9891
rect 9607 -9961 10007 -9951
rect 10063 -9891 10463 -9781
rect 10063 -9951 10073 -9891
rect 10133 -9951 10393 -9891
rect 10453 -9951 10463 -9891
rect 10063 -9961 10463 -9951
rect 10521 -9891 10921 -9781
rect 10521 -9951 10531 -9891
rect 10591 -9951 10851 -9891
rect 10911 -9951 10921 -9891
rect 10521 -9961 10921 -9951
rect 10977 -9891 11377 -9781
rect 10977 -9951 10987 -9891
rect 11047 -9951 11307 -9891
rect 11367 -9951 11377 -9891
rect 10977 -9961 11377 -9951
rect 11433 -9891 11833 -9781
rect 11433 -9951 11443 -9891
rect 11503 -9951 11763 -9891
rect 11823 -9951 11833 -9891
rect 11433 -9961 11833 -9951
rect 11891 -9891 12291 -9781
rect 11891 -9951 11901 -9891
rect 11961 -9951 12221 -9891
rect 12281 -9951 12291 -9891
rect 11891 -9961 12291 -9951
rect 12347 -9891 12747 -9781
rect 12347 -9951 12357 -9891
rect 12417 -9951 12677 -9891
rect 12737 -9951 12747 -9891
rect 12347 -9961 12747 -9951
rect 12803 -9891 13203 -9781
rect 12803 -9951 12813 -9891
rect 12873 -9951 13133 -9891
rect 13193 -9951 13203 -9891
rect 12803 -9961 13203 -9951
rect 13261 -9891 13661 -9781
rect 13261 -9951 13271 -9891
rect 13331 -9951 13591 -9891
rect 13651 -9951 13661 -9891
rect 13261 -9961 13661 -9951
rect 13717 -9891 14117 -9781
rect 13717 -9951 13727 -9891
rect 13787 -9951 14047 -9891
rect 14107 -9951 14117 -9891
rect 13717 -9961 14117 -9951
rect 14173 -9891 14573 -9781
rect 14173 -9951 14183 -9891
rect 14243 -9951 14503 -9891
rect 14563 -9951 14573 -9891
rect 14173 -9961 14573 -9951
rect 14631 -9891 15031 -9781
rect 14631 -9951 14641 -9891
rect 14701 -9951 14961 -9891
rect 15021 -9951 15031 -9891
rect 14631 -9961 15031 -9951
rect 15087 -9891 15487 -9781
rect 15087 -9951 15097 -9891
rect 15157 -9951 15417 -9891
rect 15477 -9951 15487 -9891
rect 15087 -9961 15487 -9951
rect 66 -10047 80 -9961
rect 457 -10047 527 -9961
rect 913 -10047 983 -9961
rect 1371 -10047 1441 -9961
rect 1827 -10047 1897 -9961
rect 2283 -10047 2353 -9961
rect 2741 -10047 2811 -9961
rect 3197 -10047 3267 -9961
rect 3653 -10047 3723 -9961
rect 4111 -10047 4181 -9961
rect 4567 -10047 4637 -9961
rect 5023 -10047 5093 -9961
rect 5481 -10047 5551 -9961
rect 5937 -10047 6007 -9961
rect 6393 -10047 6463 -9961
rect 6851 -10047 6921 -9961
rect 7307 -10047 7377 -9961
rect 7763 -10047 7833 -9961
rect 8237 -10047 8307 -9961
rect 8693 -10047 8763 -9961
rect 9151 -10047 9221 -9961
rect 9607 -10047 9677 -9961
rect 10063 -10047 10133 -9961
rect 10521 -10047 10591 -9961
rect 10977 -10047 11047 -9961
rect 11433 -10047 11503 -9961
rect 11891 -10047 11961 -9961
rect 12347 -10047 12417 -9961
rect 12803 -10047 12873 -9961
rect 13261 -10047 13331 -9961
rect 13717 -10047 13787 -9961
rect 14173 -10047 14243 -9961
rect 14631 -10047 14701 -9961
rect 66 -10057 400 -10047
rect 0 -10117 11 -10057
rect 71 -10117 331 -10057
rect 391 -10117 400 -10057
rect 0 -10407 14 -10117
rect 66 -10407 400 -10117
rect 0 -10467 11 -10407
rect 71 -10467 331 -10407
rect 391 -10467 400 -10407
rect 0 -10559 14 -10467
rect 66 -10477 400 -10467
rect 457 -10057 857 -10047
rect 457 -10117 467 -10057
rect 527 -10117 787 -10057
rect 847 -10117 857 -10057
rect 457 -10227 857 -10117
rect 913 -10057 1313 -10047
rect 913 -10117 923 -10057
rect 983 -10117 1243 -10057
rect 1303 -10117 1313 -10057
rect 913 -10227 1313 -10117
rect 1371 -10057 1771 -10047
rect 1371 -10117 1381 -10057
rect 1441 -10117 1701 -10057
rect 1761 -10117 1771 -10057
rect 1371 -10227 1771 -10117
rect 1827 -10057 2227 -10047
rect 1827 -10117 1837 -10057
rect 1897 -10117 2157 -10057
rect 2217 -10117 2227 -10057
rect 1827 -10227 2227 -10117
rect 2283 -10057 2683 -10047
rect 2283 -10117 2293 -10057
rect 2353 -10117 2613 -10057
rect 2673 -10117 2683 -10057
rect 2283 -10227 2683 -10117
rect 2741 -10057 3141 -10047
rect 2741 -10117 2751 -10057
rect 2811 -10117 3071 -10057
rect 3131 -10117 3141 -10057
rect 2741 -10227 3141 -10117
rect 3197 -10057 3597 -10047
rect 3197 -10117 3207 -10057
rect 3267 -10117 3527 -10057
rect 3587 -10117 3597 -10057
rect 3197 -10227 3597 -10117
rect 3653 -10057 4053 -10047
rect 3653 -10117 3663 -10057
rect 3723 -10117 3983 -10057
rect 4043 -10117 4053 -10057
rect 3653 -10227 4053 -10117
rect 457 -10297 4053 -10227
rect 457 -10407 857 -10297
rect 457 -10467 467 -10407
rect 527 -10467 787 -10407
rect 847 -10467 857 -10407
rect 457 -10477 857 -10467
rect 913 -10407 1313 -10297
rect 913 -10467 923 -10407
rect 983 -10467 1243 -10407
rect 1303 -10467 1313 -10407
rect 913 -10477 1313 -10467
rect 1371 -10407 1771 -10297
rect 1371 -10467 1381 -10407
rect 1441 -10467 1701 -10407
rect 1761 -10467 1771 -10407
rect 1371 -10477 1771 -10467
rect 1827 -10407 2227 -10297
rect 1827 -10467 1837 -10407
rect 1897 -10467 2157 -10407
rect 2217 -10467 2227 -10407
rect 1827 -10477 2227 -10467
rect 2283 -10407 2683 -10297
rect 2283 -10467 2293 -10407
rect 2353 -10467 2613 -10407
rect 2673 -10467 2683 -10407
rect 2283 -10477 2683 -10467
rect 2741 -10407 3141 -10297
rect 2741 -10467 2751 -10407
rect 2811 -10467 3071 -10407
rect 3131 -10467 3141 -10407
rect 2741 -10477 3141 -10467
rect 3197 -10407 3597 -10297
rect 3197 -10467 3207 -10407
rect 3267 -10467 3527 -10407
rect 3587 -10467 3597 -10407
rect 3197 -10477 3597 -10467
rect 3653 -10407 4053 -10297
rect 3653 -10467 3663 -10407
rect 3723 -10467 3983 -10407
rect 4043 -10467 4053 -10407
rect 3653 -10477 4053 -10467
rect 4111 -10057 4511 -10047
rect 4111 -10117 4121 -10057
rect 4181 -10117 4441 -10057
rect 4501 -10117 4511 -10057
rect 4111 -10227 4511 -10117
rect 4567 -10057 4967 -10047
rect 4567 -10117 4577 -10057
rect 4637 -10117 4897 -10057
rect 4957 -10117 4967 -10057
rect 4567 -10227 4967 -10117
rect 5023 -10057 5423 -10047
rect 5023 -10117 5033 -10057
rect 5093 -10117 5353 -10057
rect 5413 -10117 5423 -10057
rect 5023 -10227 5423 -10117
rect 5481 -10057 5881 -10047
rect 5481 -10117 5491 -10057
rect 5551 -10117 5811 -10057
rect 5871 -10117 5881 -10057
rect 5481 -10227 5881 -10117
rect 5937 -10057 6337 -10047
rect 5937 -10117 5947 -10057
rect 6007 -10117 6267 -10057
rect 6327 -10117 6337 -10057
rect 5937 -10227 6337 -10117
rect 6393 -10057 6793 -10047
rect 6393 -10117 6403 -10057
rect 6463 -10117 6723 -10057
rect 6783 -10117 6793 -10057
rect 6393 -10227 6793 -10117
rect 6851 -10057 7251 -10047
rect 6851 -10117 6861 -10057
rect 6921 -10117 7181 -10057
rect 7241 -10117 7251 -10057
rect 6851 -10227 7251 -10117
rect 4111 -10297 7251 -10227
rect 4111 -10407 4511 -10297
rect 4111 -10467 4121 -10407
rect 4181 -10467 4441 -10407
rect 4501 -10467 4511 -10407
rect 4111 -10477 4511 -10467
rect 4567 -10407 4967 -10297
rect 4567 -10467 4577 -10407
rect 4637 -10467 4897 -10407
rect 4957 -10467 4967 -10407
rect 4567 -10477 4967 -10467
rect 5023 -10407 5423 -10297
rect 5023 -10467 5033 -10407
rect 5093 -10467 5353 -10407
rect 5413 -10467 5423 -10407
rect 5023 -10477 5423 -10467
rect 5481 -10407 5881 -10297
rect 5481 -10467 5491 -10407
rect 5551 -10467 5811 -10407
rect 5871 -10467 5881 -10407
rect 5481 -10477 5881 -10467
rect 5937 -10407 6337 -10297
rect 5937 -10467 5947 -10407
rect 6007 -10467 6267 -10407
rect 6327 -10467 6337 -10407
rect 5937 -10477 6337 -10467
rect 6393 -10407 6793 -10297
rect 6393 -10467 6403 -10407
rect 6463 -10467 6723 -10407
rect 6783 -10467 6793 -10407
rect 6393 -10477 6793 -10467
rect 6851 -10407 7251 -10297
rect 6851 -10467 6861 -10407
rect 6921 -10467 7181 -10407
rect 7241 -10467 7251 -10407
rect 6851 -10477 7251 -10467
rect 7307 -10057 7707 -10047
rect 7307 -10117 7317 -10057
rect 7377 -10117 7637 -10057
rect 7697 -10117 7707 -10057
rect 7307 -10227 7707 -10117
rect 7763 -10057 8163 -10047
rect 7763 -10117 7773 -10057
rect 7833 -10117 8093 -10057
rect 8153 -10117 8163 -10057
rect 7763 -10227 8163 -10117
rect 8237 -10057 8637 -10047
rect 8237 -10117 8247 -10057
rect 8307 -10117 8567 -10057
rect 8627 -10117 8637 -10057
rect 8237 -10227 8637 -10117
rect 8693 -10057 9093 -10047
rect 8693 -10117 8703 -10057
rect 8763 -10117 9023 -10057
rect 9083 -10117 9093 -10057
rect 8693 -10227 9093 -10117
rect 9151 -10057 9551 -10047
rect 9151 -10117 9161 -10057
rect 9221 -10117 9481 -10057
rect 9541 -10117 9551 -10057
rect 9151 -10227 9551 -10117
rect 9607 -10057 10007 -10047
rect 9607 -10117 9617 -10057
rect 9677 -10117 9937 -10057
rect 9997 -10117 10007 -10057
rect 9607 -10227 10007 -10117
rect 10063 -10057 10463 -10047
rect 10063 -10117 10073 -10057
rect 10133 -10117 10393 -10057
rect 10453 -10117 10463 -10057
rect 10063 -10227 10463 -10117
rect 10521 -10057 10921 -10047
rect 10521 -10117 10531 -10057
rect 10591 -10117 10851 -10057
rect 10911 -10117 10921 -10057
rect 10521 -10227 10921 -10117
rect 10977 -10057 11377 -10047
rect 10977 -10117 10987 -10057
rect 11047 -10117 11307 -10057
rect 11367 -10117 11377 -10057
rect 10977 -10227 11377 -10117
rect 11433 -10057 11833 -10047
rect 11433 -10117 11443 -10057
rect 11503 -10117 11763 -10057
rect 11823 -10117 11833 -10057
rect 11433 -10227 11833 -10117
rect 11891 -10057 12291 -10047
rect 11891 -10117 11901 -10057
rect 11961 -10117 12221 -10057
rect 12281 -10117 12291 -10057
rect 11891 -10227 12291 -10117
rect 12347 -10057 12747 -10047
rect 12347 -10117 12357 -10057
rect 12417 -10117 12677 -10057
rect 12737 -10117 12747 -10057
rect 12347 -10227 12747 -10117
rect 12803 -10057 13203 -10047
rect 12803 -10117 12813 -10057
rect 12873 -10117 13133 -10057
rect 13193 -10117 13203 -10057
rect 12803 -10227 13203 -10117
rect 13261 -10057 13661 -10047
rect 13261 -10117 13271 -10057
rect 13331 -10117 13591 -10057
rect 13651 -10117 13661 -10057
rect 13261 -10227 13661 -10117
rect 13717 -10057 14117 -10047
rect 13717 -10117 13727 -10057
rect 13787 -10117 14047 -10057
rect 14107 -10117 14117 -10057
rect 13717 -10227 14117 -10117
rect 14173 -10057 14573 -10047
rect 14173 -10117 14183 -10057
rect 14243 -10117 14503 -10057
rect 14563 -10117 14573 -10057
rect 14173 -10227 14573 -10117
rect 14631 -10057 15031 -10047
rect 14631 -10117 14641 -10057
rect 14701 -10117 14961 -10057
rect 15021 -10117 15031 -10057
rect 14631 -10227 15031 -10117
rect 15087 -10057 15487 -10047
rect 15087 -10117 15097 -10057
rect 15157 -10117 15417 -10057
rect 15477 -10117 15487 -10057
rect 15087 -10227 15487 -10117
rect 7307 -10297 15487 -10227
rect 7307 -10407 7707 -10297
rect 7307 -10467 7317 -10407
rect 7377 -10467 7637 -10407
rect 7697 -10467 7707 -10407
rect 7307 -10477 7707 -10467
rect 7763 -10407 8163 -10297
rect 7763 -10467 7773 -10407
rect 7833 -10467 8093 -10407
rect 8153 -10467 8163 -10407
rect 7763 -10477 8163 -10467
rect 8237 -10407 8637 -10297
rect 8237 -10467 8247 -10407
rect 8307 -10467 8567 -10407
rect 8627 -10467 8637 -10407
rect 8237 -10477 8637 -10467
rect 8693 -10407 9093 -10297
rect 8693 -10467 8703 -10407
rect 8763 -10467 9023 -10407
rect 9083 -10467 9093 -10407
rect 8693 -10477 9093 -10467
rect 9151 -10407 9551 -10297
rect 9151 -10467 9161 -10407
rect 9221 -10467 9481 -10407
rect 9541 -10467 9551 -10407
rect 9151 -10477 9551 -10467
rect 9607 -10407 10007 -10297
rect 9607 -10467 9617 -10407
rect 9677 -10467 9937 -10407
rect 9997 -10467 10007 -10407
rect 9607 -10477 10007 -10467
rect 10063 -10407 10463 -10297
rect 10063 -10467 10073 -10407
rect 10133 -10467 10393 -10407
rect 10453 -10467 10463 -10407
rect 10063 -10477 10463 -10467
rect 10521 -10407 10921 -10297
rect 10521 -10467 10531 -10407
rect 10591 -10467 10851 -10407
rect 10911 -10467 10921 -10407
rect 10521 -10477 10921 -10467
rect 10977 -10407 11377 -10297
rect 10977 -10467 10987 -10407
rect 11047 -10467 11307 -10407
rect 11367 -10467 11377 -10407
rect 10977 -10477 11377 -10467
rect 11433 -10407 11833 -10297
rect 11433 -10467 11443 -10407
rect 11503 -10467 11763 -10407
rect 11823 -10467 11833 -10407
rect 11433 -10477 11833 -10467
rect 11891 -10407 12291 -10297
rect 11891 -10467 11901 -10407
rect 11961 -10467 12221 -10407
rect 12281 -10467 12291 -10407
rect 11891 -10477 12291 -10467
rect 12347 -10407 12747 -10297
rect 12347 -10467 12357 -10407
rect 12417 -10467 12677 -10407
rect 12737 -10467 12747 -10407
rect 12347 -10477 12747 -10467
rect 12803 -10407 13203 -10297
rect 12803 -10467 12813 -10407
rect 12873 -10467 13133 -10407
rect 13193 -10467 13203 -10407
rect 12803 -10477 13203 -10467
rect 13261 -10407 13661 -10297
rect 13261 -10467 13271 -10407
rect 13331 -10467 13591 -10407
rect 13651 -10467 13661 -10407
rect 13261 -10477 13661 -10467
rect 13717 -10407 14117 -10297
rect 13717 -10467 13727 -10407
rect 13787 -10467 14047 -10407
rect 14107 -10467 14117 -10407
rect 13717 -10477 14117 -10467
rect 14173 -10407 14573 -10297
rect 14173 -10467 14183 -10407
rect 14243 -10467 14503 -10407
rect 14563 -10467 14573 -10407
rect 14173 -10477 14573 -10467
rect 14631 -10407 15031 -10297
rect 14631 -10467 14641 -10407
rect 14701 -10467 14961 -10407
rect 15021 -10467 15031 -10407
rect 14631 -10477 15031 -10467
rect 15087 -10407 15487 -10297
rect 15087 -10467 15097 -10407
rect 15157 -10467 15417 -10407
rect 15477 -10467 15487 -10407
rect 15087 -10477 15487 -10467
rect 66 -10549 80 -10477
rect 457 -10549 527 -10477
rect 913 -10549 984 -10477
rect 1371 -10549 1442 -10477
rect 1827 -10549 1898 -10477
rect 2283 -10549 2354 -10477
rect 2741 -10549 2812 -10477
rect 3197 -10549 3268 -10477
rect 3653 -10549 3724 -10477
rect 4111 -10549 4182 -10477
rect 4567 -10549 4638 -10477
rect 5023 -10549 5094 -10477
rect 5481 -10549 5552 -10477
rect 5937 -10549 6008 -10477
rect 6393 -10549 6464 -10477
rect 6851 -10549 6922 -10477
rect 7307 -10549 7378 -10477
rect 7763 -10549 7834 -10477
rect 8237 -10549 8308 -10477
rect 8693 -10549 8764 -10477
rect 9151 -10549 9222 -10477
rect 9607 -10549 9678 -10477
rect 10063 -10549 10134 -10477
rect 10521 -10549 10592 -10477
rect 10977 -10549 11048 -10477
rect 11433 -10549 11504 -10477
rect 11891 -10549 11962 -10477
rect 12347 -10549 12418 -10477
rect 12803 -10549 12874 -10477
rect 13261 -10549 13332 -10477
rect 13717 -10549 13788 -10477
rect 14173 -10549 14244 -10477
rect 14631 -10549 14702 -10477
rect 66 -10559 400 -10549
rect 0 -10619 11 -10559
rect 71 -10619 331 -10559
rect 391 -10619 400 -10559
rect 0 -10909 14 -10619
rect 66 -10909 400 -10619
rect 0 -10969 11 -10909
rect 71 -10969 331 -10909
rect 391 -10969 400 -10909
rect 0 -11051 14 -10969
rect 66 -10979 400 -10969
rect 457 -10559 857 -10549
rect 457 -10619 467 -10559
rect 527 -10619 787 -10559
rect 847 -10619 857 -10559
rect 457 -10729 857 -10619
rect 913 -10559 1313 -10549
rect 913 -10619 923 -10559
rect 983 -10619 1243 -10559
rect 1303 -10619 1313 -10559
rect 913 -10729 1313 -10619
rect 1371 -10559 1771 -10549
rect 1371 -10619 1381 -10559
rect 1441 -10619 1701 -10559
rect 1761 -10619 1771 -10559
rect 1371 -10729 1771 -10619
rect 1827 -10559 2227 -10549
rect 1827 -10619 1837 -10559
rect 1897 -10619 2157 -10559
rect 2217 -10619 2227 -10559
rect 1827 -10729 2227 -10619
rect 2283 -10559 2683 -10549
rect 2283 -10619 2293 -10559
rect 2353 -10619 2613 -10559
rect 2673 -10619 2683 -10559
rect 2283 -10729 2683 -10619
rect 457 -10730 2683 -10729
rect 2741 -10559 3141 -10549
rect 2741 -10619 2751 -10559
rect 2811 -10619 3071 -10559
rect 3131 -10619 3141 -10559
rect 2741 -10729 3141 -10619
rect 3197 -10559 3597 -10549
rect 3197 -10619 3207 -10559
rect 3267 -10619 3527 -10559
rect 3587 -10619 3597 -10559
rect 3197 -10729 3597 -10619
rect 3653 -10559 4053 -10549
rect 3653 -10619 3663 -10559
rect 3723 -10619 3983 -10559
rect 4043 -10619 4053 -10559
rect 3653 -10729 4053 -10619
rect 2741 -10730 4053 -10729
rect 457 -10800 4053 -10730
rect 457 -10909 857 -10800
rect 457 -10969 467 -10909
rect 527 -10969 787 -10909
rect 847 -10969 857 -10909
rect 457 -10979 857 -10969
rect 913 -10909 1313 -10800
rect 913 -10969 923 -10909
rect 983 -10969 1243 -10909
rect 1303 -10969 1313 -10909
rect 913 -10979 1313 -10969
rect 1371 -10909 1771 -10800
rect 1371 -10969 1381 -10909
rect 1441 -10969 1701 -10909
rect 1761 -10969 1771 -10909
rect 1371 -10979 1771 -10969
rect 1827 -10909 2227 -10800
rect 1827 -10969 1837 -10909
rect 1897 -10969 2157 -10909
rect 2217 -10969 2227 -10909
rect 1827 -10979 2227 -10969
rect 2283 -10909 2683 -10800
rect 2283 -10969 2293 -10909
rect 2353 -10969 2613 -10909
rect 2673 -10969 2683 -10909
rect 2283 -10979 2683 -10969
rect 2741 -10909 3141 -10800
rect 2741 -10969 2751 -10909
rect 2811 -10969 3071 -10909
rect 3131 -10969 3141 -10909
rect 2741 -10979 3141 -10969
rect 3197 -10909 3597 -10800
rect 3197 -10969 3207 -10909
rect 3267 -10969 3527 -10909
rect 3587 -10969 3597 -10909
rect 3197 -10979 3597 -10969
rect 3653 -10909 4053 -10800
rect 3653 -10969 3663 -10909
rect 3723 -10969 3983 -10909
rect 4043 -10969 4053 -10909
rect 3653 -10979 4053 -10969
rect 4111 -10559 4511 -10549
rect 4111 -10619 4121 -10559
rect 4181 -10619 4441 -10559
rect 4501 -10619 4511 -10559
rect 4111 -10729 4511 -10619
rect 4567 -10559 4967 -10549
rect 4567 -10619 4577 -10559
rect 4637 -10619 4897 -10559
rect 4957 -10619 4967 -10559
rect 4567 -10729 4967 -10619
rect 5023 -10559 5423 -10549
rect 5023 -10619 5033 -10559
rect 5093 -10619 5353 -10559
rect 5413 -10619 5423 -10559
rect 5023 -10729 5423 -10619
rect 5481 -10559 5881 -10549
rect 5481 -10619 5491 -10559
rect 5551 -10619 5811 -10559
rect 5871 -10619 5881 -10559
rect 5481 -10729 5881 -10619
rect 5937 -10559 6337 -10549
rect 5937 -10619 5947 -10559
rect 6007 -10619 6267 -10559
rect 6327 -10619 6337 -10559
rect 5937 -10729 6337 -10619
rect 6393 -10559 6793 -10549
rect 6393 -10619 6403 -10559
rect 6463 -10619 6723 -10559
rect 6783 -10619 6793 -10559
rect 6393 -10729 6793 -10619
rect 6851 -10559 7251 -10549
rect 6851 -10619 6861 -10559
rect 6921 -10619 7181 -10559
rect 7241 -10619 7251 -10559
rect 6851 -10729 7251 -10619
rect 4111 -10800 7251 -10729
rect 4111 -10909 4511 -10800
rect 4111 -10969 4121 -10909
rect 4181 -10969 4441 -10909
rect 4501 -10969 4511 -10909
rect 4111 -10979 4511 -10969
rect 4567 -10909 4967 -10800
rect 4567 -10969 4577 -10909
rect 4637 -10969 4897 -10909
rect 4957 -10969 4967 -10909
rect 4567 -10979 4967 -10969
rect 5023 -10909 5423 -10800
rect 5023 -10969 5033 -10909
rect 5093 -10969 5353 -10909
rect 5413 -10969 5423 -10909
rect 5023 -10979 5423 -10969
rect 5481 -10909 5881 -10800
rect 5481 -10969 5491 -10909
rect 5551 -10969 5811 -10909
rect 5871 -10969 5881 -10909
rect 5481 -10979 5881 -10969
rect 5937 -10909 6337 -10800
rect 5937 -10969 5947 -10909
rect 6007 -10969 6267 -10909
rect 6327 -10969 6337 -10909
rect 5937 -10979 6337 -10969
rect 6393 -10909 6793 -10800
rect 6393 -10969 6403 -10909
rect 6463 -10969 6723 -10909
rect 6783 -10969 6793 -10909
rect 6393 -10979 6793 -10969
rect 6851 -10909 7251 -10800
rect 6851 -10969 6861 -10909
rect 6921 -10969 7181 -10909
rect 7241 -10969 7251 -10909
rect 6851 -10979 7251 -10969
rect 7307 -10559 7707 -10549
rect 7307 -10619 7317 -10559
rect 7377 -10619 7637 -10559
rect 7697 -10619 7707 -10559
rect 7307 -10729 7707 -10619
rect 7763 -10559 8163 -10549
rect 7763 -10619 7773 -10559
rect 7833 -10619 8093 -10559
rect 8153 -10619 8163 -10559
rect 7763 -10729 8163 -10619
rect 8237 -10559 8637 -10549
rect 8237 -10619 8247 -10559
rect 8307 -10619 8567 -10559
rect 8627 -10619 8637 -10559
rect 8237 -10729 8637 -10619
rect 8693 -10559 9093 -10549
rect 8693 -10619 8703 -10559
rect 8763 -10619 9023 -10559
rect 9083 -10619 9093 -10559
rect 8693 -10729 9093 -10619
rect 9151 -10559 9551 -10549
rect 9151 -10619 9161 -10559
rect 9221 -10619 9481 -10559
rect 9541 -10619 9551 -10559
rect 9151 -10729 9551 -10619
rect 9607 -10559 10007 -10549
rect 9607 -10619 9617 -10559
rect 9677 -10619 9937 -10559
rect 9997 -10619 10007 -10559
rect 9607 -10729 10007 -10619
rect 10063 -10559 10463 -10549
rect 10063 -10619 10073 -10559
rect 10133 -10619 10393 -10559
rect 10453 -10619 10463 -10559
rect 10063 -10729 10463 -10619
rect 7307 -10730 10463 -10729
rect 10521 -10559 10921 -10549
rect 10521 -10619 10531 -10559
rect 10591 -10619 10851 -10559
rect 10911 -10619 10921 -10559
rect 10521 -10729 10921 -10619
rect 10977 -10559 11377 -10549
rect 10977 -10619 10987 -10559
rect 11047 -10619 11307 -10559
rect 11367 -10619 11377 -10559
rect 10977 -10729 11377 -10619
rect 11433 -10559 11833 -10549
rect 11433 -10619 11443 -10559
rect 11503 -10619 11763 -10559
rect 11823 -10619 11833 -10559
rect 11433 -10729 11833 -10619
rect 11891 -10559 12291 -10549
rect 11891 -10619 11901 -10559
rect 11961 -10619 12221 -10559
rect 12281 -10619 12291 -10559
rect 11891 -10729 12291 -10619
rect 12347 -10559 12747 -10549
rect 12347 -10619 12357 -10559
rect 12417 -10619 12677 -10559
rect 12737 -10619 12747 -10559
rect 12347 -10729 12747 -10619
rect 12803 -10559 13203 -10549
rect 12803 -10619 12813 -10559
rect 12873 -10619 13133 -10559
rect 13193 -10619 13203 -10559
rect 12803 -10729 13203 -10619
rect 13261 -10559 13661 -10549
rect 13261 -10619 13271 -10559
rect 13331 -10619 13591 -10559
rect 13651 -10619 13661 -10559
rect 13261 -10729 13661 -10619
rect 13717 -10559 14117 -10549
rect 13717 -10619 13727 -10559
rect 13787 -10619 14047 -10559
rect 14107 -10619 14117 -10559
rect 13717 -10729 14117 -10619
rect 14173 -10559 14573 -10549
rect 14173 -10619 14183 -10559
rect 14243 -10619 14503 -10559
rect 14563 -10619 14573 -10559
rect 14173 -10729 14573 -10619
rect 14631 -10559 15031 -10549
rect 14631 -10619 14641 -10559
rect 14701 -10619 14961 -10559
rect 15021 -10619 15031 -10559
rect 14631 -10729 15031 -10619
rect 15087 -10559 15487 -10549
rect 15087 -10619 15097 -10559
rect 15157 -10619 15417 -10559
rect 15477 -10619 15487 -10559
rect 15087 -10729 15487 -10619
rect 10521 -10730 15487 -10729
rect 7307 -10800 15487 -10730
rect 7307 -10909 7707 -10800
rect 7307 -10969 7317 -10909
rect 7377 -10969 7637 -10909
rect 7697 -10969 7707 -10909
rect 7307 -10979 7707 -10969
rect 7763 -10909 8163 -10800
rect 7763 -10969 7773 -10909
rect 7833 -10969 8093 -10909
rect 8153 -10969 8163 -10909
rect 7763 -10979 8163 -10969
rect 8237 -10909 8637 -10800
rect 8237 -10969 8247 -10909
rect 8307 -10969 8567 -10909
rect 8627 -10969 8637 -10909
rect 8237 -10979 8637 -10969
rect 8693 -10909 9093 -10800
rect 8693 -10969 8703 -10909
rect 8763 -10969 9023 -10909
rect 9083 -10969 9093 -10909
rect 8693 -10979 9093 -10969
rect 9151 -10909 9551 -10800
rect 9151 -10969 9161 -10909
rect 9221 -10969 9481 -10909
rect 9541 -10969 9551 -10909
rect 9151 -10979 9551 -10969
rect 9607 -10909 10007 -10800
rect 9607 -10969 9617 -10909
rect 9677 -10969 9937 -10909
rect 9997 -10969 10007 -10909
rect 9607 -10979 10007 -10969
rect 10063 -10909 10463 -10800
rect 10063 -10969 10073 -10909
rect 10133 -10969 10393 -10909
rect 10453 -10969 10463 -10909
rect 10063 -10979 10463 -10969
rect 10521 -10909 10921 -10800
rect 10521 -10969 10531 -10909
rect 10591 -10969 10851 -10909
rect 10911 -10969 10921 -10909
rect 10521 -10979 10921 -10969
rect 10977 -10909 11377 -10800
rect 10977 -10969 10987 -10909
rect 11047 -10969 11307 -10909
rect 11367 -10969 11377 -10909
rect 10977 -10979 11377 -10969
rect 11433 -10909 11833 -10800
rect 11433 -10969 11443 -10909
rect 11503 -10969 11763 -10909
rect 11823 -10969 11833 -10909
rect 11433 -10979 11833 -10969
rect 11891 -10909 12291 -10800
rect 11891 -10969 11901 -10909
rect 11961 -10969 12221 -10909
rect 12281 -10969 12291 -10909
rect 11891 -10979 12291 -10969
rect 12347 -10909 12747 -10800
rect 12347 -10969 12357 -10909
rect 12417 -10969 12677 -10909
rect 12737 -10969 12747 -10909
rect 12347 -10979 12747 -10969
rect 12803 -10909 13203 -10800
rect 12803 -10969 12813 -10909
rect 12873 -10969 13133 -10909
rect 13193 -10969 13203 -10909
rect 12803 -10979 13203 -10969
rect 13261 -10909 13661 -10800
rect 13261 -10969 13271 -10909
rect 13331 -10969 13591 -10909
rect 13651 -10969 13661 -10909
rect 13261 -10979 13661 -10969
rect 13717 -10909 14117 -10800
rect 13717 -10969 13727 -10909
rect 13787 -10969 14047 -10909
rect 14107 -10969 14117 -10909
rect 13717 -10979 14117 -10969
rect 14173 -10909 14573 -10800
rect 14173 -10969 14183 -10909
rect 14243 -10969 14503 -10909
rect 14563 -10969 14573 -10909
rect 14173 -10979 14573 -10969
rect 14631 -10909 15031 -10800
rect 14631 -10969 14641 -10909
rect 14701 -10969 14961 -10909
rect 15021 -10969 15031 -10909
rect 14631 -10979 15031 -10969
rect 15087 -10909 15487 -10800
rect 15087 -10969 15097 -10909
rect 15157 -10969 15417 -10909
rect 15477 -10969 15487 -10909
rect 15087 -10979 15487 -10969
rect 66 -11041 80 -10979
rect 457 -11041 528 -10979
rect 913 -11041 984 -10979
rect 1371 -11041 1442 -10979
rect 1827 -11041 1898 -10979
rect 2283 -11041 2354 -10979
rect 2741 -11041 2811 -10979
rect 3197 -11041 3267 -10979
rect 3653 -11041 3723 -10979
rect 4111 -11041 4181 -10979
rect 4567 -11041 4637 -10979
rect 5023 -11041 5093 -10979
rect 5481 -11041 5551 -10979
rect 5937 -11041 6007 -10979
rect 6393 -11041 6463 -10979
rect 6851 -11041 6921 -10979
rect 7307 -11041 7377 -10979
rect 7763 -11041 7833 -10979
rect 8237 -11041 8307 -10979
rect 8693 -11041 8763 -10979
rect 9151 -11041 9221 -10979
rect 66 -11051 400 -11041
rect 0 -11111 11 -11051
rect 71 -11111 331 -11051
rect 391 -11111 400 -11051
rect 0 -11401 14 -11111
rect 66 -11401 400 -11111
rect 0 -11461 11 -11401
rect 71 -11461 331 -11401
rect 391 -11461 400 -11401
rect 0 -11544 14 -11461
rect 66 -11471 400 -11461
rect 457 -11051 857 -11041
rect 457 -11111 467 -11051
rect 527 -11111 787 -11051
rect 847 -11111 857 -11051
rect 457 -11221 857 -11111
rect 913 -11051 1313 -11041
rect 913 -11111 923 -11051
rect 983 -11111 1243 -11051
rect 1303 -11111 1313 -11051
rect 913 -11221 1313 -11111
rect 1371 -11051 1771 -11041
rect 1371 -11111 1381 -11051
rect 1441 -11111 1701 -11051
rect 1761 -11111 1771 -11051
rect 1371 -11221 1771 -11111
rect 1827 -11051 2227 -11041
rect 1827 -11111 1837 -11051
rect 1897 -11111 2157 -11051
rect 2217 -11111 2227 -11051
rect 1827 -11221 2227 -11111
rect 2283 -11051 2683 -11041
rect 2283 -11111 2293 -11051
rect 2353 -11111 2613 -11051
rect 2673 -11111 2683 -11051
rect 2283 -11221 2683 -11111
rect 2741 -11051 3141 -11041
rect 2741 -11111 2751 -11051
rect 2811 -11111 3071 -11051
rect 3131 -11111 3141 -11051
rect 2741 -11221 3141 -11111
rect 3197 -11051 3597 -11041
rect 3197 -11111 3207 -11051
rect 3267 -11111 3527 -11051
rect 3587 -11111 3597 -11051
rect 3197 -11221 3597 -11111
rect 3653 -11051 4053 -11041
rect 3653 -11111 3663 -11051
rect 3723 -11111 3983 -11051
rect 4043 -11111 4053 -11051
rect 3653 -11221 4053 -11111
rect 457 -11291 4053 -11221
rect 457 -11401 857 -11291
rect 457 -11461 467 -11401
rect 527 -11461 787 -11401
rect 847 -11461 857 -11401
rect 457 -11471 857 -11461
rect 913 -11401 1313 -11291
rect 913 -11461 923 -11401
rect 983 -11461 1243 -11401
rect 1303 -11461 1313 -11401
rect 913 -11471 1313 -11461
rect 1371 -11401 1771 -11291
rect 1371 -11461 1381 -11401
rect 1441 -11461 1701 -11401
rect 1761 -11461 1771 -11401
rect 1371 -11471 1771 -11461
rect 1827 -11401 2227 -11291
rect 1827 -11461 1837 -11401
rect 1897 -11461 2157 -11401
rect 2217 -11461 2227 -11401
rect 1827 -11471 2227 -11461
rect 2283 -11401 2683 -11291
rect 2283 -11461 2293 -11401
rect 2353 -11461 2613 -11401
rect 2673 -11461 2683 -11401
rect 2283 -11471 2683 -11461
rect 2741 -11401 3141 -11291
rect 2741 -11461 2751 -11401
rect 2811 -11461 3071 -11401
rect 3131 -11461 3141 -11401
rect 2741 -11471 3141 -11461
rect 3197 -11401 3597 -11291
rect 3197 -11461 3207 -11401
rect 3267 -11461 3527 -11401
rect 3587 -11461 3597 -11401
rect 3197 -11471 3597 -11461
rect 3653 -11401 4053 -11291
rect 3653 -11461 3663 -11401
rect 3723 -11461 3983 -11401
rect 4043 -11461 4053 -11401
rect 3653 -11471 4053 -11461
rect 4111 -11051 4511 -11041
rect 4111 -11111 4121 -11051
rect 4181 -11111 4441 -11051
rect 4501 -11111 4511 -11051
rect 4111 -11221 4511 -11111
rect 4567 -11051 4967 -11041
rect 4567 -11111 4577 -11051
rect 4637 -11111 4897 -11051
rect 4957 -11111 4967 -11051
rect 4567 -11221 4967 -11111
rect 5023 -11051 5423 -11041
rect 5023 -11111 5033 -11051
rect 5093 -11111 5353 -11051
rect 5413 -11111 5423 -11051
rect 5023 -11221 5423 -11111
rect 5481 -11051 5881 -11041
rect 5481 -11111 5491 -11051
rect 5551 -11111 5811 -11051
rect 5871 -11111 5881 -11051
rect 5481 -11221 5881 -11111
rect 5937 -11051 6337 -11041
rect 5937 -11111 5947 -11051
rect 6007 -11111 6267 -11051
rect 6327 -11111 6337 -11051
rect 5937 -11221 6337 -11111
rect 6393 -11051 6793 -11041
rect 6393 -11111 6403 -11051
rect 6463 -11111 6723 -11051
rect 6783 -11111 6793 -11051
rect 6393 -11221 6793 -11111
rect 6851 -11051 7251 -11041
rect 6851 -11111 6861 -11051
rect 6921 -11111 7181 -11051
rect 7241 -11111 7251 -11051
rect 6851 -11221 7251 -11111
rect 4111 -11291 7251 -11221
rect 4111 -11401 4511 -11291
rect 4111 -11461 4121 -11401
rect 4181 -11461 4441 -11401
rect 4501 -11461 4511 -11401
rect 4111 -11471 4511 -11461
rect 4567 -11401 4967 -11291
rect 4567 -11461 4577 -11401
rect 4637 -11461 4897 -11401
rect 4957 -11461 4967 -11401
rect 4567 -11471 4967 -11461
rect 5023 -11401 5423 -11291
rect 5023 -11461 5033 -11401
rect 5093 -11461 5353 -11401
rect 5413 -11461 5423 -11401
rect 5023 -11471 5423 -11461
rect 5481 -11401 5881 -11291
rect 5481 -11461 5491 -11401
rect 5551 -11461 5811 -11401
rect 5871 -11461 5881 -11401
rect 5481 -11471 5881 -11461
rect 5937 -11401 6337 -11291
rect 5937 -11461 5947 -11401
rect 6007 -11461 6267 -11401
rect 6327 -11461 6337 -11401
rect 5937 -11471 6337 -11461
rect 6393 -11401 6793 -11291
rect 6393 -11461 6403 -11401
rect 6463 -11461 6723 -11401
rect 6783 -11461 6793 -11401
rect 6393 -11471 6793 -11461
rect 6851 -11401 7251 -11291
rect 6851 -11461 6861 -11401
rect 6921 -11461 7181 -11401
rect 7241 -11461 7251 -11401
rect 6851 -11471 7251 -11461
rect 7307 -11051 7707 -11041
rect 7307 -11111 7317 -11051
rect 7377 -11111 7637 -11051
rect 7697 -11111 7707 -11051
rect 7307 -11221 7707 -11111
rect 7763 -11051 8163 -11041
rect 7763 -11111 7773 -11051
rect 7833 -11111 8093 -11051
rect 8153 -11111 8163 -11051
rect 7763 -11221 8163 -11111
rect 8237 -11051 8637 -11041
rect 8237 -11111 8247 -11051
rect 8307 -11111 8567 -11051
rect 8627 -11111 8637 -11051
rect 8237 -11221 8637 -11111
rect 8693 -11051 9093 -11041
rect 8693 -11111 8703 -11051
rect 8763 -11111 9023 -11051
rect 9083 -11111 9093 -11051
rect 8693 -11221 9093 -11111
rect 9151 -11051 9551 -11041
rect 9151 -11111 9161 -11051
rect 9221 -11111 9481 -11051
rect 9541 -11111 9551 -11051
rect 9151 -11170 9551 -11111
rect 9607 -11051 10007 -11041
rect 9607 -11111 9617 -11051
rect 9677 -11111 9937 -11051
rect 9997 -11111 10007 -11051
rect 9151 -11221 9550 -11170
rect 7307 -11291 9550 -11221
rect 7307 -11401 7707 -11291
rect 7307 -11461 7317 -11401
rect 7377 -11461 7637 -11401
rect 7697 -11461 7707 -11401
rect 7307 -11471 7707 -11461
rect 7763 -11401 8163 -11291
rect 7763 -11461 7773 -11401
rect 7833 -11461 8093 -11401
rect 8153 -11461 8163 -11401
rect 7763 -11471 8163 -11461
rect 8237 -11401 8637 -11291
rect 8237 -11461 8247 -11401
rect 8307 -11461 8567 -11401
rect 8627 -11461 8637 -11401
rect 8237 -11471 8637 -11461
rect 8693 -11401 9093 -11291
rect 8693 -11461 8703 -11401
rect 8763 -11461 9023 -11401
rect 9083 -11461 9093 -11401
rect 8693 -11471 9093 -11461
rect 9151 -11401 9550 -11291
rect 9151 -11461 9161 -11401
rect 9221 -11461 9481 -11401
rect 9541 -11461 9550 -11401
rect 9151 -11471 9550 -11461
rect 9607 -11221 10007 -11111
rect 10063 -11051 10463 -11041
rect 10063 -11111 10073 -11051
rect 10133 -11111 10393 -11051
rect 10453 -11111 10463 -11051
rect 10063 -11221 10463 -11111
rect 10521 -11051 10921 -11041
rect 10521 -11111 10531 -11051
rect 10591 -11111 10851 -11051
rect 10911 -11111 10921 -11051
rect 10521 -11221 10921 -11111
rect 10977 -11051 11377 -11041
rect 10977 -11111 10987 -11051
rect 11047 -11111 11307 -11051
rect 11367 -11111 11377 -11051
rect 10977 -11221 11377 -11111
rect 11433 -11051 11833 -11041
rect 11433 -11111 11443 -11051
rect 11503 -11111 11763 -11051
rect 11823 -11111 11833 -11051
rect 11433 -11221 11833 -11111
rect 11891 -11051 12291 -11041
rect 11891 -11111 11901 -11051
rect 11961 -11111 12221 -11051
rect 12281 -11111 12291 -11051
rect 11891 -11221 12291 -11111
rect 12347 -11051 12747 -11041
rect 12347 -11111 12357 -11051
rect 12417 -11111 12677 -11051
rect 12737 -11111 12747 -11051
rect 12347 -11221 12747 -11111
rect 12803 -11051 13203 -11041
rect 12803 -11111 12813 -11051
rect 12873 -11111 13133 -11051
rect 13193 -11111 13203 -11051
rect 12803 -11221 13203 -11111
rect 13261 -11051 13661 -11041
rect 13261 -11111 13271 -11051
rect 13331 -11111 13591 -11051
rect 13651 -11111 13661 -11051
rect 13261 -11221 13661 -11111
rect 13717 -11051 14117 -11041
rect 13717 -11111 13727 -11051
rect 13787 -11111 14047 -11051
rect 14107 -11111 14117 -11051
rect 13717 -11221 14117 -11111
rect 14173 -11051 14573 -11041
rect 14173 -11111 14183 -11051
rect 14243 -11111 14503 -11051
rect 14563 -11111 14573 -11051
rect 14173 -11221 14573 -11111
rect 14631 -11051 15031 -11041
rect 14631 -11111 14641 -11051
rect 14701 -11111 14961 -11051
rect 15021 -11111 15031 -11051
rect 14631 -11221 15031 -11111
rect 15087 -11051 15487 -11041
rect 15087 -11111 15097 -11051
rect 15157 -11111 15417 -11051
rect 15477 -11111 15487 -11051
rect 15087 -11221 15487 -11111
rect 9607 -11291 15487 -11221
rect 9607 -11401 10007 -11291
rect 9607 -11461 9617 -11401
rect 9677 -11461 9937 -11401
rect 9997 -11461 10007 -11401
rect 9607 -11471 10007 -11461
rect 10063 -11401 10463 -11291
rect 10063 -11461 10073 -11401
rect 10133 -11461 10393 -11401
rect 10453 -11461 10463 -11401
rect 10063 -11471 10463 -11461
rect 10521 -11401 10921 -11291
rect 10521 -11461 10531 -11401
rect 10591 -11461 10851 -11401
rect 10911 -11461 10921 -11401
rect 10521 -11471 10921 -11461
rect 10977 -11401 11377 -11291
rect 10977 -11461 10987 -11401
rect 11047 -11461 11307 -11401
rect 11367 -11461 11377 -11401
rect 10977 -11471 11377 -11461
rect 11433 -11401 11833 -11291
rect 11433 -11461 11443 -11401
rect 11503 -11461 11763 -11401
rect 11823 -11461 11833 -11401
rect 11433 -11471 11833 -11461
rect 11891 -11401 12291 -11291
rect 11891 -11461 11901 -11401
rect 11961 -11461 12221 -11401
rect 12281 -11461 12291 -11401
rect 11891 -11471 12291 -11461
rect 12347 -11401 12747 -11291
rect 12347 -11461 12357 -11401
rect 12417 -11461 12677 -11401
rect 12737 -11461 12747 -11401
rect 12347 -11471 12747 -11461
rect 12803 -11401 13203 -11291
rect 12803 -11461 12813 -11401
rect 12873 -11461 13133 -11401
rect 13193 -11461 13203 -11401
rect 12803 -11471 13203 -11461
rect 13261 -11401 13661 -11291
rect 13261 -11461 13271 -11401
rect 13331 -11461 13591 -11401
rect 13651 -11461 13661 -11401
rect 13261 -11471 13661 -11461
rect 13717 -11401 14117 -11291
rect 13717 -11461 13727 -11401
rect 13787 -11461 14047 -11401
rect 14107 -11461 14117 -11401
rect 13717 -11471 14117 -11461
rect 14173 -11401 14573 -11291
rect 14173 -11461 14183 -11401
rect 14243 -11461 14503 -11401
rect 14563 -11461 14573 -11401
rect 14173 -11471 14573 -11461
rect 14631 -11401 15031 -11291
rect 14631 -11461 14641 -11401
rect 14701 -11461 14961 -11401
rect 15021 -11461 15031 -11401
rect 14631 -11471 15031 -11461
rect 15087 -11401 15487 -11291
rect 15087 -11461 15097 -11401
rect 15157 -11461 15417 -11401
rect 15477 -11461 15487 -11401
rect 15087 -11471 15487 -11461
rect 66 -11534 80 -11471
rect 457 -11489 527 -11471
rect 913 -11489 983 -11471
rect 1371 -11489 1441 -11471
rect 1827 -11489 1897 -11471
rect 2283 -11489 2353 -11471
rect 2741 -11489 2811 -11471
rect 3197 -11489 3267 -11471
rect 3653 -11489 3723 -11471
rect 4111 -11489 4181 -11471
rect 4567 -11489 4637 -11471
rect 5023 -11489 5093 -11471
rect 5481 -11489 5551 -11471
rect 5937 -11489 6007 -11471
rect 6393 -11489 6463 -11471
rect 6851 -11489 6921 -11471
rect 7307 -11489 7377 -11471
rect 7763 -11489 7833 -11471
rect 8237 -11489 8307 -11471
rect 8693 -11489 8763 -11471
rect 9151 -11489 9221 -11471
rect 456 -11534 527 -11489
rect 912 -11534 983 -11489
rect 1370 -11534 1441 -11489
rect 1826 -11534 1897 -11489
rect 2282 -11534 2353 -11489
rect 2740 -11534 2811 -11489
rect 3196 -11534 3267 -11489
rect 3652 -11534 3723 -11489
rect 4110 -11534 4181 -11489
rect 4566 -11534 4637 -11489
rect 5022 -11534 5093 -11489
rect 5480 -11534 5551 -11489
rect 5936 -11534 6007 -11489
rect 6392 -11534 6463 -11489
rect 6850 -11534 6921 -11489
rect 7306 -11534 7377 -11489
rect 7762 -11534 7833 -11489
rect 8236 -11534 8307 -11489
rect 8692 -11534 8763 -11489
rect 9150 -11534 9221 -11489
rect 9607 -11534 9677 -11471
rect 10063 -11489 10133 -11471
rect 10521 -11489 10591 -11471
rect 10977 -11489 11047 -11471
rect 11433 -11489 11503 -11471
rect 11891 -11489 11961 -11471
rect 12347 -11489 12417 -11471
rect 12803 -11489 12873 -11471
rect 13261 -11489 13331 -11471
rect 13717 -11489 13787 -11471
rect 14173 -11489 14243 -11471
rect 14631 -11489 14701 -11471
rect 10062 -11534 10133 -11489
rect 10520 -11534 10591 -11489
rect 10976 -11534 11047 -11489
rect 11432 -11534 11503 -11489
rect 11890 -11534 11961 -11489
rect 12346 -11534 12417 -11489
rect 12802 -11534 12873 -11489
rect 13260 -11534 13331 -11489
rect 13716 -11534 13787 -11489
rect 14172 -11534 14243 -11489
rect 14630 -11534 14701 -11489
rect 66 -11544 400 -11534
rect 0 -11604 10 -11544
rect 70 -11604 330 -11544
rect 390 -11604 400 -11544
rect 0 -11894 14 -11604
rect 66 -11894 400 -11604
rect 0 -11954 10 -11894
rect 70 -11954 330 -11894
rect 390 -11954 400 -11894
rect 0 -12036 14 -11954
rect 66 -11964 400 -11954
rect 456 -11544 856 -11534
rect 456 -11604 466 -11544
rect 526 -11604 786 -11544
rect 846 -11604 856 -11544
rect 456 -11714 856 -11604
rect 912 -11544 1312 -11534
rect 912 -11604 922 -11544
rect 982 -11604 1242 -11544
rect 1302 -11604 1312 -11544
rect 912 -11714 1312 -11604
rect 1370 -11544 1770 -11534
rect 1370 -11604 1380 -11544
rect 1440 -11604 1700 -11544
rect 1760 -11604 1770 -11544
rect 1370 -11714 1770 -11604
rect 1826 -11544 2226 -11534
rect 1826 -11604 1836 -11544
rect 1896 -11604 2156 -11544
rect 2216 -11604 2226 -11544
rect 1826 -11714 2226 -11604
rect 2282 -11544 2682 -11534
rect 2282 -11604 2292 -11544
rect 2352 -11604 2612 -11544
rect 2672 -11604 2682 -11544
rect 2282 -11714 2682 -11604
rect 2740 -11544 3140 -11534
rect 2740 -11604 2750 -11544
rect 2810 -11604 3070 -11544
rect 3130 -11604 3140 -11544
rect 2740 -11714 3140 -11604
rect 3196 -11544 3596 -11534
rect 3196 -11604 3206 -11544
rect 3266 -11604 3526 -11544
rect 3586 -11604 3596 -11544
rect 3196 -11714 3596 -11604
rect 3652 -11544 4052 -11534
rect 3652 -11604 3662 -11544
rect 3722 -11604 3982 -11544
rect 4042 -11604 4052 -11544
rect 3652 -11714 4052 -11604
rect 456 -11784 4052 -11714
rect 456 -11894 856 -11784
rect 456 -11954 466 -11894
rect 526 -11954 786 -11894
rect 846 -11954 856 -11894
rect 456 -11964 856 -11954
rect 912 -11894 1312 -11784
rect 912 -11954 922 -11894
rect 982 -11954 1242 -11894
rect 1302 -11954 1312 -11894
rect 912 -11964 1312 -11954
rect 1370 -11894 1770 -11784
rect 1370 -11954 1380 -11894
rect 1440 -11954 1700 -11894
rect 1760 -11954 1770 -11894
rect 1370 -11964 1770 -11954
rect 1826 -11894 2226 -11784
rect 1826 -11954 1836 -11894
rect 1896 -11954 2156 -11894
rect 2216 -11954 2226 -11894
rect 1826 -11964 2226 -11954
rect 2282 -11894 2682 -11784
rect 2282 -11954 2292 -11894
rect 2352 -11954 2612 -11894
rect 2672 -11954 2682 -11894
rect 2282 -11964 2682 -11954
rect 2740 -11894 3140 -11784
rect 2740 -11954 2750 -11894
rect 2810 -11954 3070 -11894
rect 3130 -11954 3140 -11894
rect 2740 -11964 3140 -11954
rect 3196 -11894 3596 -11784
rect 3196 -11954 3206 -11894
rect 3266 -11954 3526 -11894
rect 3586 -11954 3596 -11894
rect 3196 -11964 3596 -11954
rect 3652 -11894 4052 -11784
rect 3652 -11954 3662 -11894
rect 3722 -11954 3982 -11894
rect 4042 -11954 4052 -11894
rect 3652 -11964 4052 -11954
rect 4110 -11544 4510 -11534
rect 4110 -11604 4120 -11544
rect 4180 -11604 4440 -11544
rect 4500 -11604 4510 -11544
rect 4110 -11714 4510 -11604
rect 4566 -11544 4966 -11534
rect 4566 -11604 4576 -11544
rect 4636 -11604 4896 -11544
rect 4956 -11604 4966 -11544
rect 4566 -11714 4966 -11604
rect 5022 -11544 5422 -11534
rect 5022 -11604 5032 -11544
rect 5092 -11604 5352 -11544
rect 5412 -11604 5422 -11544
rect 5022 -11714 5422 -11604
rect 5480 -11544 5880 -11534
rect 5480 -11604 5490 -11544
rect 5550 -11604 5810 -11544
rect 5870 -11604 5880 -11544
rect 5480 -11714 5880 -11604
rect 5936 -11544 6336 -11534
rect 5936 -11604 5946 -11544
rect 6006 -11604 6266 -11544
rect 6326 -11604 6336 -11544
rect 5936 -11714 6336 -11604
rect 6392 -11544 6792 -11534
rect 6392 -11604 6402 -11544
rect 6462 -11604 6722 -11544
rect 6782 -11604 6792 -11544
rect 6392 -11714 6792 -11604
rect 6850 -11544 7250 -11534
rect 6850 -11604 6860 -11544
rect 6920 -11604 7180 -11544
rect 7240 -11604 7250 -11544
rect 6850 -11714 7250 -11604
rect 4110 -11784 7250 -11714
rect 4110 -11894 4510 -11784
rect 4110 -11954 4120 -11894
rect 4180 -11954 4440 -11894
rect 4500 -11954 4510 -11894
rect 4110 -11964 4510 -11954
rect 4566 -11894 4966 -11784
rect 4566 -11954 4576 -11894
rect 4636 -11954 4896 -11894
rect 4956 -11954 4966 -11894
rect 4566 -11964 4966 -11954
rect 5022 -11894 5422 -11784
rect 5022 -11954 5032 -11894
rect 5092 -11954 5352 -11894
rect 5412 -11954 5422 -11894
rect 5022 -11964 5422 -11954
rect 5480 -11894 5880 -11784
rect 5480 -11954 5490 -11894
rect 5550 -11954 5810 -11894
rect 5870 -11954 5880 -11894
rect 5480 -11964 5880 -11954
rect 5936 -11894 6336 -11784
rect 5936 -11954 5946 -11894
rect 6006 -11954 6266 -11894
rect 6326 -11954 6336 -11894
rect 5936 -11964 6336 -11954
rect 6392 -11894 6792 -11784
rect 6392 -11954 6402 -11894
rect 6462 -11954 6722 -11894
rect 6782 -11954 6792 -11894
rect 6392 -11964 6792 -11954
rect 6850 -11894 7250 -11784
rect 6850 -11954 6860 -11894
rect 6920 -11954 7180 -11894
rect 7240 -11954 7250 -11894
rect 6850 -11964 7250 -11954
rect 7306 -11544 7706 -11534
rect 7306 -11604 7316 -11544
rect 7376 -11604 7636 -11544
rect 7696 -11604 7706 -11544
rect 7306 -11714 7706 -11604
rect 7762 -11544 8162 -11534
rect 7762 -11604 7772 -11544
rect 7832 -11604 8092 -11544
rect 8152 -11604 8162 -11544
rect 7762 -11714 8162 -11604
rect 8236 -11544 8636 -11534
rect 8236 -11604 8246 -11544
rect 8306 -11604 8566 -11544
rect 8626 -11604 8636 -11544
rect 8236 -11714 8636 -11604
rect 8692 -11544 9092 -11534
rect 8692 -11604 8702 -11544
rect 8762 -11604 9022 -11544
rect 9082 -11604 9092 -11544
rect 8692 -11714 9092 -11604
rect 9150 -11544 9550 -11534
rect 9150 -11604 9160 -11544
rect 9220 -11604 9480 -11544
rect 9540 -11604 9550 -11544
rect 9150 -11714 9550 -11604
rect 7306 -11784 9550 -11714
rect 7306 -11894 7706 -11784
rect 7306 -11954 7316 -11894
rect 7376 -11954 7636 -11894
rect 7696 -11954 7706 -11894
rect 7306 -11964 7706 -11954
rect 7762 -11894 8162 -11784
rect 7762 -11954 7772 -11894
rect 7832 -11954 8092 -11894
rect 8152 -11954 8162 -11894
rect 7762 -11964 8162 -11954
rect 8236 -11894 8636 -11784
rect 8236 -11954 8246 -11894
rect 8306 -11954 8566 -11894
rect 8626 -11954 8636 -11894
rect 8236 -11964 8636 -11954
rect 8692 -11894 9092 -11784
rect 8692 -11954 8702 -11894
rect 8762 -11954 9022 -11894
rect 9082 -11954 9092 -11894
rect 8692 -11964 9092 -11954
rect 9150 -11894 9550 -11784
rect 9607 -11544 10006 -11534
rect 9607 -11604 9616 -11544
rect 9676 -11604 9936 -11544
rect 9996 -11604 10006 -11544
rect 9607 -11714 10006 -11604
rect 10062 -11544 10462 -11534
rect 10062 -11604 10072 -11544
rect 10132 -11604 10392 -11544
rect 10452 -11604 10462 -11544
rect 10062 -11714 10462 -11604
rect 10520 -11544 10920 -11534
rect 10520 -11604 10530 -11544
rect 10590 -11604 10850 -11544
rect 10910 -11604 10920 -11544
rect 10520 -11714 10920 -11604
rect 10976 -11544 11376 -11534
rect 10976 -11604 10986 -11544
rect 11046 -11604 11306 -11544
rect 11366 -11604 11376 -11544
rect 10976 -11714 11376 -11604
rect 11432 -11544 11832 -11534
rect 11432 -11604 11442 -11544
rect 11502 -11604 11762 -11544
rect 11822 -11604 11832 -11544
rect 11432 -11714 11832 -11604
rect 11890 -11544 12290 -11534
rect 11890 -11604 11900 -11544
rect 11960 -11604 12220 -11544
rect 12280 -11604 12290 -11544
rect 11890 -11714 12290 -11604
rect 12346 -11544 12746 -11534
rect 12346 -11604 12356 -11544
rect 12416 -11604 12676 -11544
rect 12736 -11604 12746 -11544
rect 12346 -11714 12746 -11604
rect 12802 -11544 13202 -11534
rect 12802 -11604 12812 -11544
rect 12872 -11604 13132 -11544
rect 13192 -11604 13202 -11544
rect 12802 -11714 13202 -11604
rect 13260 -11544 13660 -11534
rect 13260 -11604 13270 -11544
rect 13330 -11604 13590 -11544
rect 13650 -11604 13660 -11544
rect 13260 -11714 13660 -11604
rect 13716 -11544 14116 -11534
rect 13716 -11604 13726 -11544
rect 13786 -11604 14046 -11544
rect 14106 -11604 14116 -11544
rect 13716 -11714 14116 -11604
rect 14172 -11544 14572 -11534
rect 14172 -11604 14182 -11544
rect 14242 -11604 14502 -11544
rect 14562 -11604 14572 -11544
rect 14172 -11714 14572 -11604
rect 14630 -11544 15030 -11534
rect 14630 -11604 14640 -11544
rect 14700 -11604 14960 -11544
rect 15020 -11604 15030 -11544
rect 14630 -11714 15030 -11604
rect 15086 -11544 15486 -11534
rect 15086 -11604 15096 -11544
rect 15156 -11604 15416 -11544
rect 15476 -11604 15486 -11544
rect 15086 -11714 15486 -11604
rect 9607 -11784 15486 -11714
rect 9607 -11787 10006 -11784
rect 9150 -11954 9160 -11894
rect 9220 -11954 9480 -11894
rect 9540 -11954 9550 -11894
rect 9150 -11964 9550 -11954
rect 9606 -11894 10006 -11787
rect 9606 -11954 9616 -11894
rect 9676 -11954 9936 -11894
rect 9996 -11954 10006 -11894
rect 9606 -11964 10006 -11954
rect 10062 -11894 10462 -11784
rect 10062 -11954 10072 -11894
rect 10132 -11954 10392 -11894
rect 10452 -11954 10462 -11894
rect 10062 -11964 10462 -11954
rect 10520 -11894 10920 -11784
rect 10520 -11954 10530 -11894
rect 10590 -11954 10850 -11894
rect 10910 -11954 10920 -11894
rect 10520 -11964 10920 -11954
rect 10976 -11894 11376 -11784
rect 10976 -11954 10986 -11894
rect 11046 -11954 11306 -11894
rect 11366 -11954 11376 -11894
rect 10976 -11964 11376 -11954
rect 11432 -11894 11832 -11784
rect 11432 -11954 11442 -11894
rect 11502 -11954 11762 -11894
rect 11822 -11954 11832 -11894
rect 11432 -11964 11832 -11954
rect 11890 -11894 12290 -11784
rect 11890 -11954 11900 -11894
rect 11960 -11954 12220 -11894
rect 12280 -11954 12290 -11894
rect 11890 -11964 12290 -11954
rect 12346 -11894 12746 -11784
rect 12346 -11954 12356 -11894
rect 12416 -11954 12676 -11894
rect 12736 -11954 12746 -11894
rect 12346 -11964 12746 -11954
rect 12802 -11894 13202 -11784
rect 12802 -11954 12812 -11894
rect 12872 -11954 13132 -11894
rect 13192 -11954 13202 -11894
rect 12802 -11964 13202 -11954
rect 13260 -11894 13660 -11784
rect 13260 -11954 13270 -11894
rect 13330 -11954 13590 -11894
rect 13650 -11954 13660 -11894
rect 13260 -11964 13660 -11954
rect 13716 -11894 14116 -11784
rect 13716 -11954 13726 -11894
rect 13786 -11954 14046 -11894
rect 14106 -11954 14116 -11894
rect 13716 -11964 14116 -11954
rect 14172 -11894 14572 -11784
rect 14172 -11954 14182 -11894
rect 14242 -11954 14502 -11894
rect 14562 -11954 14572 -11894
rect 14172 -11964 14572 -11954
rect 14630 -11894 15030 -11784
rect 14630 -11954 14640 -11894
rect 14700 -11954 14960 -11894
rect 15020 -11954 15030 -11894
rect 14630 -11964 15030 -11954
rect 15086 -11894 15486 -11784
rect 15086 -11954 15096 -11894
rect 15156 -11954 15416 -11894
rect 15476 -11954 15486 -11894
rect 15086 -11964 15486 -11954
rect 66 -12026 80 -11964
rect 456 -12026 527 -11964
rect 912 -12026 983 -11964
rect 1370 -12026 1441 -11964
rect 1826 -12026 1897 -11964
rect 2282 -12026 2353 -11964
rect 2740 -12026 2810 -11964
rect 3196 -12026 3266 -11964
rect 4110 -12026 4180 -11964
rect 4566 -12026 4636 -11964
rect 5022 -12026 5092 -11964
rect 5480 -12026 5550 -11964
rect 5936 -12026 6006 -11964
rect 6392 -12026 6462 -11964
rect 6850 -12026 6920 -11964
rect 7306 -12026 7376 -11964
rect 7762 -12026 7832 -11964
rect 8236 -12026 8306 -11964
rect 8692 -12026 8762 -11964
rect 9606 -12026 9676 -11964
rect 10062 -12026 10132 -11964
rect 10520 -12026 10590 -11964
rect 10976 -12026 11046 -11964
rect 11432 -12026 11502 -11964
rect 11890 -12026 11960 -11964
rect 12346 -12026 12416 -11964
rect 12802 -12026 12872 -11964
rect 13260 -12026 13330 -11964
rect 13716 -12026 13786 -11964
rect 14172 -12026 14242 -11964
rect 14630 -12026 14700 -11964
rect 66 -12036 400 -12026
rect 0 -12096 10 -12036
rect 70 -12096 330 -12036
rect 390 -12096 400 -12036
rect 0 -12386 14 -12096
rect 66 -12386 400 -12096
rect 0 -12446 10 -12386
rect 70 -12446 330 -12386
rect 390 -12446 400 -12386
rect 0 -12552 14 -12446
rect 66 -12456 400 -12446
rect 456 -12036 856 -12026
rect 456 -12096 466 -12036
rect 526 -12096 786 -12036
rect 846 -12096 856 -12036
rect 456 -12206 856 -12096
rect 912 -12036 1312 -12026
rect 912 -12096 922 -12036
rect 982 -12096 1242 -12036
rect 1302 -12096 1312 -12036
rect 912 -12206 1312 -12096
rect 1370 -12036 1770 -12026
rect 1370 -12096 1380 -12036
rect 1440 -12096 1700 -12036
rect 1760 -12096 1770 -12036
rect 1370 -12206 1770 -12096
rect 1826 -12036 2226 -12026
rect 1826 -12096 1836 -12036
rect 1896 -12096 2156 -12036
rect 2216 -12096 2226 -12036
rect 1826 -12206 2226 -12096
rect 2282 -12036 2682 -12026
rect 2282 -12096 2292 -12036
rect 2352 -12096 2612 -12036
rect 2672 -12096 2682 -12036
rect 2282 -12206 2682 -12096
rect 456 -12207 2682 -12206
rect 2740 -12036 3140 -12026
rect 2740 -12096 2750 -12036
rect 2810 -12096 3070 -12036
rect 3130 -12096 3140 -12036
rect 2740 -12206 3140 -12096
rect 3196 -12036 3596 -12026
rect 3196 -12096 3206 -12036
rect 3266 -12096 3526 -12036
rect 3586 -12096 3596 -12036
rect 3196 -12206 3596 -12096
rect 2740 -12207 3596 -12206
rect 456 -12277 3596 -12207
rect 456 -12386 856 -12277
rect 456 -12446 466 -12386
rect 526 -12446 786 -12386
rect 846 -12446 856 -12386
rect 456 -12456 856 -12446
rect 912 -12386 1312 -12277
rect 912 -12446 922 -12386
rect 982 -12446 1242 -12386
rect 1302 -12446 1312 -12386
rect 912 -12456 1312 -12446
rect 1370 -12386 1770 -12277
rect 1370 -12446 1380 -12386
rect 1440 -12446 1700 -12386
rect 1760 -12446 1770 -12386
rect 1370 -12456 1770 -12446
rect 1826 -12386 2226 -12277
rect 1826 -12446 1836 -12386
rect 1896 -12446 2156 -12386
rect 2216 -12446 2226 -12386
rect 1826 -12456 2226 -12446
rect 2282 -12386 2682 -12277
rect 2282 -12446 2292 -12386
rect 2352 -12446 2612 -12386
rect 2672 -12446 2682 -12386
rect 2282 -12456 2682 -12446
rect 2740 -12386 3140 -12277
rect 2740 -12446 2750 -12386
rect 2810 -12446 3070 -12386
rect 3130 -12446 3140 -12386
rect 2740 -12456 3140 -12446
rect 3196 -12386 3596 -12277
rect 3196 -12446 3206 -12386
rect 3266 -12446 3526 -12386
rect 3586 -12446 3596 -12386
rect 3196 -12456 3596 -12446
rect 3652 -12036 4052 -12026
rect 3652 -12096 3662 -12036
rect 3722 -12096 3982 -12036
rect 4042 -12096 4052 -12036
rect 3652 -12206 4052 -12096
rect 4110 -12036 4510 -12026
rect 4110 -12096 4120 -12036
rect 4180 -12096 4440 -12036
rect 4500 -12096 4510 -12036
rect 4110 -12206 4510 -12096
rect 4566 -12036 4966 -12026
rect 4566 -12096 4576 -12036
rect 4636 -12096 4896 -12036
rect 4956 -12096 4966 -12036
rect 4566 -12206 4966 -12096
rect 5022 -12036 5422 -12026
rect 5022 -12096 5032 -12036
rect 5092 -12096 5352 -12036
rect 5412 -12096 5422 -12036
rect 5022 -12206 5422 -12096
rect 5480 -12036 5880 -12026
rect 5480 -12096 5490 -12036
rect 5550 -12096 5810 -12036
rect 5870 -12096 5880 -12036
rect 5480 -12206 5880 -12096
rect 5936 -12036 6336 -12026
rect 5936 -12096 5946 -12036
rect 6006 -12096 6266 -12036
rect 6326 -12096 6336 -12036
rect 5936 -12206 6336 -12096
rect 6392 -12036 6792 -12026
rect 6392 -12096 6402 -12036
rect 6462 -12096 6722 -12036
rect 6782 -12096 6792 -12036
rect 6392 -12206 6792 -12096
rect 6850 -12036 7250 -12026
rect 6850 -12096 6860 -12036
rect 6920 -12096 7180 -12036
rect 7240 -12096 7250 -12036
rect 6850 -12206 7250 -12096
rect 3652 -12277 7250 -12206
rect 3652 -12386 4052 -12277
rect 3652 -12446 3662 -12386
rect 3722 -12446 3982 -12386
rect 4042 -12446 4052 -12386
rect 3652 -12456 4052 -12446
rect 4110 -12386 4510 -12277
rect 4110 -12446 4120 -12386
rect 4180 -12446 4440 -12386
rect 4500 -12446 4510 -12386
rect 4110 -12456 4510 -12446
rect 4566 -12386 4966 -12277
rect 4566 -12446 4576 -12386
rect 4636 -12446 4896 -12386
rect 4956 -12446 4966 -12386
rect 4566 -12456 4966 -12446
rect 5022 -12386 5422 -12277
rect 5022 -12446 5032 -12386
rect 5092 -12446 5352 -12386
rect 5412 -12446 5422 -12386
rect 5022 -12456 5422 -12446
rect 5480 -12386 5880 -12277
rect 5480 -12446 5490 -12386
rect 5550 -12446 5810 -12386
rect 5870 -12446 5880 -12386
rect 5480 -12456 5880 -12446
rect 5936 -12386 6336 -12277
rect 5936 -12446 5946 -12386
rect 6006 -12446 6266 -12386
rect 6326 -12446 6336 -12386
rect 5936 -12456 6336 -12446
rect 6392 -12386 6792 -12277
rect 6392 -12446 6402 -12386
rect 6462 -12446 6722 -12386
rect 6782 -12446 6792 -12386
rect 6392 -12456 6792 -12446
rect 6850 -12386 7250 -12277
rect 6850 -12446 6860 -12386
rect 6920 -12446 7180 -12386
rect 7240 -12446 7250 -12386
rect 6850 -12456 7250 -12446
rect 7306 -12036 7706 -12026
rect 7306 -12096 7316 -12036
rect 7376 -12096 7636 -12036
rect 7696 -12096 7706 -12036
rect 7306 -12206 7706 -12096
rect 7762 -12036 8162 -12026
rect 7762 -12096 7772 -12036
rect 7832 -12096 8092 -12036
rect 8152 -12096 8162 -12036
rect 7762 -12206 8162 -12096
rect 8236 -12036 8636 -12026
rect 8236 -12096 8246 -12036
rect 8306 -12096 8566 -12036
rect 8626 -12096 8636 -12036
rect 8236 -12206 8636 -12096
rect 8692 -12036 9092 -12026
rect 8692 -12096 8702 -12036
rect 8762 -12096 9022 -12036
rect 9082 -12096 9092 -12036
rect 8692 -12206 9092 -12096
rect 9150 -12036 9550 -12026
rect 9150 -12096 9160 -12036
rect 9220 -12096 9480 -12036
rect 9540 -12096 9550 -12036
rect 9150 -12206 9550 -12096
rect 9606 -12036 10006 -12026
rect 9606 -12096 9616 -12036
rect 9676 -12096 9936 -12036
rect 9996 -12096 10006 -12036
rect 9606 -12206 10006 -12096
rect 10062 -12036 10462 -12026
rect 10062 -12096 10072 -12036
rect 10132 -12096 10392 -12036
rect 10452 -12096 10462 -12036
rect 10062 -12206 10462 -12096
rect 7306 -12277 9093 -12206
rect 9150 -12207 10462 -12206
rect 10520 -12036 10920 -12026
rect 10520 -12096 10530 -12036
rect 10590 -12096 10850 -12036
rect 10910 -12096 10920 -12036
rect 10520 -12206 10920 -12096
rect 10976 -12036 11376 -12026
rect 10976 -12096 10986 -12036
rect 11046 -12096 11306 -12036
rect 11366 -12096 11376 -12036
rect 10976 -12206 11376 -12096
rect 11432 -12036 11832 -12026
rect 11432 -12096 11442 -12036
rect 11502 -12096 11762 -12036
rect 11822 -12096 11832 -12036
rect 11432 -12206 11832 -12096
rect 11890 -12036 12290 -12026
rect 11890 -12096 11900 -12036
rect 11960 -12096 12220 -12036
rect 12280 -12096 12290 -12036
rect 11890 -12206 12290 -12096
rect 12346 -12036 12746 -12026
rect 12346 -12096 12356 -12036
rect 12416 -12096 12676 -12036
rect 12736 -12096 12746 -12036
rect 12346 -12206 12746 -12096
rect 12802 -12036 13202 -12026
rect 12802 -12096 12812 -12036
rect 12872 -12096 13132 -12036
rect 13192 -12096 13202 -12036
rect 12802 -12206 13202 -12096
rect 13260 -12036 13660 -12026
rect 13260 -12096 13270 -12036
rect 13330 -12096 13590 -12036
rect 13650 -12096 13660 -12036
rect 13260 -12206 13660 -12096
rect 13716 -12036 14116 -12026
rect 13716 -12096 13726 -12036
rect 13786 -12096 14046 -12036
rect 14106 -12096 14116 -12036
rect 13716 -12206 14116 -12096
rect 14172 -12036 14572 -12026
rect 14172 -12096 14182 -12036
rect 14242 -12096 14502 -12036
rect 14562 -12096 14572 -12036
rect 14172 -12206 14572 -12096
rect 14630 -12036 15030 -12026
rect 14630 -12096 14640 -12036
rect 14700 -12096 14960 -12036
rect 15020 -12096 15030 -12036
rect 14630 -12206 15030 -12096
rect 15086 -12036 15486 -12026
rect 15086 -12096 15096 -12036
rect 15156 -12096 15416 -12036
rect 15476 -12096 15486 -12036
rect 15086 -12206 15486 -12096
rect 10520 -12207 15486 -12206
rect 9150 -12277 15486 -12207
rect 7306 -12386 7706 -12277
rect 7306 -12446 7316 -12386
rect 7376 -12446 7636 -12386
rect 7696 -12446 7706 -12386
rect 7306 -12456 7706 -12446
rect 7762 -12386 8162 -12277
rect 7762 -12446 7772 -12386
rect 7832 -12446 8092 -12386
rect 8152 -12446 8162 -12386
rect 7762 -12456 8162 -12446
rect 8236 -12386 8636 -12277
rect 8236 -12446 8246 -12386
rect 8306 -12446 8566 -12386
rect 8626 -12446 8636 -12386
rect 8236 -12456 8636 -12446
rect 8692 -12386 9092 -12277
rect 8692 -12446 8702 -12386
rect 8762 -12446 9022 -12386
rect 9082 -12446 9092 -12386
rect 8692 -12456 9092 -12446
rect 9150 -12386 9550 -12277
rect 9150 -12446 9160 -12386
rect 9220 -12446 9480 -12386
rect 9540 -12446 9550 -12386
rect 9150 -12456 9550 -12446
rect 9606 -12386 10006 -12277
rect 9606 -12446 9616 -12386
rect 9676 -12446 9936 -12386
rect 9996 -12446 10006 -12386
rect 9606 -12456 10006 -12446
rect 10062 -12386 10462 -12277
rect 10062 -12446 10072 -12386
rect 10132 -12446 10392 -12386
rect 10452 -12446 10462 -12386
rect 10062 -12456 10462 -12446
rect 10520 -12386 10920 -12277
rect 10520 -12446 10530 -12386
rect 10590 -12446 10850 -12386
rect 10910 -12446 10920 -12386
rect 10520 -12456 10920 -12446
rect 10976 -12386 11376 -12277
rect 10976 -12446 10986 -12386
rect 11046 -12446 11306 -12386
rect 11366 -12446 11376 -12386
rect 10976 -12456 11376 -12446
rect 11432 -12386 11832 -12277
rect 11432 -12446 11442 -12386
rect 11502 -12446 11762 -12386
rect 11822 -12446 11832 -12386
rect 11432 -12456 11832 -12446
rect 11890 -12386 12290 -12277
rect 11890 -12446 11900 -12386
rect 11960 -12446 12220 -12386
rect 12280 -12446 12290 -12386
rect 11890 -12456 12290 -12446
rect 12346 -12386 12746 -12277
rect 12346 -12446 12356 -12386
rect 12416 -12446 12676 -12386
rect 12736 -12446 12746 -12386
rect 12346 -12456 12746 -12446
rect 12802 -12386 13202 -12277
rect 12802 -12446 12812 -12386
rect 12872 -12446 13132 -12386
rect 13192 -12446 13202 -12386
rect 12802 -12456 13202 -12446
rect 13260 -12386 13660 -12277
rect 13260 -12446 13270 -12386
rect 13330 -12446 13590 -12386
rect 13650 -12446 13660 -12386
rect 13260 -12456 13660 -12446
rect 13716 -12386 14116 -12277
rect 13716 -12446 13726 -12386
rect 13786 -12446 14046 -12386
rect 14106 -12446 14116 -12386
rect 13716 -12456 14116 -12446
rect 14172 -12386 14572 -12277
rect 14172 -12446 14182 -12386
rect 14242 -12446 14502 -12386
rect 14562 -12446 14572 -12386
rect 14172 -12456 14572 -12446
rect 14630 -12386 15030 -12277
rect 14630 -12446 14640 -12386
rect 14700 -12446 14960 -12386
rect 15020 -12446 15030 -12386
rect 14630 -12456 15030 -12446
rect 15086 -12386 15486 -12277
rect 15086 -12446 15096 -12386
rect 15156 -12446 15416 -12386
rect 15476 -12446 15486 -12386
rect 15086 -12456 15486 -12446
rect 66 -12542 80 -12456
rect 456 -12542 526 -12456
rect 912 -12542 982 -12456
rect 1370 -12542 1440 -12456
rect 1826 -12542 1896 -12456
rect 2282 -12542 2352 -12456
rect 2740 -12542 2810 -12456
rect 3196 -12542 3266 -12456
rect 3652 -12542 3722 -12456
rect 4110 -12542 4180 -12456
rect 4566 -12542 4636 -12456
rect 5022 -12542 5092 -12456
rect 5480 -12542 5550 -12456
rect 5936 -12542 6006 -12456
rect 6392 -12542 6462 -12456
rect 6850 -12542 6920 -12456
rect 7306 -12542 7376 -12456
rect 7762 -12542 7832 -12456
rect 8236 -12542 8306 -12456
rect 8692 -12542 8762 -12456
rect 9150 -12542 9220 -12456
rect 9606 -12542 9676 -12456
rect 10062 -12542 10132 -12456
rect 10520 -12542 10590 -12456
rect 66 -12552 400 -12542
rect 0 -12612 10 -12552
rect 70 -12612 330 -12552
rect 390 -12612 400 -12552
rect 0 -12902 14 -12612
rect 66 -12902 400 -12612
rect 0 -12962 10 -12902
rect 70 -12962 330 -12902
rect 390 -12962 400 -12902
rect 0 -13054 14 -12962
rect 66 -12972 400 -12962
rect 456 -12552 856 -12542
rect 456 -12612 466 -12552
rect 526 -12612 786 -12552
rect 846 -12612 856 -12552
rect 456 -12722 856 -12612
rect 912 -12552 1312 -12542
rect 912 -12612 922 -12552
rect 982 -12612 1242 -12552
rect 1302 -12612 1312 -12552
rect 912 -12722 1312 -12612
rect 1370 -12552 1770 -12542
rect 1370 -12612 1380 -12552
rect 1440 -12612 1700 -12552
rect 1760 -12612 1770 -12552
rect 1370 -12722 1770 -12612
rect 1826 -12552 2226 -12542
rect 1826 -12612 1836 -12552
rect 1896 -12612 2156 -12552
rect 2216 -12612 2226 -12552
rect 1826 -12722 2226 -12612
rect 2282 -12552 2682 -12542
rect 2282 -12612 2292 -12552
rect 2352 -12612 2612 -12552
rect 2672 -12612 2682 -12552
rect 2282 -12722 2682 -12612
rect 2740 -12552 3140 -12542
rect 2740 -12612 2750 -12552
rect 2810 -12612 3070 -12552
rect 3130 -12612 3140 -12552
rect 2740 -12722 3140 -12612
rect 3196 -12552 3596 -12542
rect 3196 -12612 3206 -12552
rect 3266 -12612 3526 -12552
rect 3586 -12612 3596 -12552
rect 3196 -12722 3596 -12612
rect 456 -12792 3596 -12722
rect 456 -12902 856 -12792
rect 456 -12962 466 -12902
rect 526 -12962 786 -12902
rect 846 -12962 856 -12902
rect 456 -12972 856 -12962
rect 912 -12902 1312 -12792
rect 912 -12962 922 -12902
rect 982 -12962 1242 -12902
rect 1302 -12962 1312 -12902
rect 912 -12972 1312 -12962
rect 1370 -12902 1770 -12792
rect 1370 -12962 1380 -12902
rect 1440 -12962 1700 -12902
rect 1760 -12962 1770 -12902
rect 1370 -12972 1770 -12962
rect 1826 -12902 2226 -12792
rect 1826 -12962 1836 -12902
rect 1896 -12962 2156 -12902
rect 2216 -12962 2226 -12902
rect 1826 -12972 2226 -12962
rect 2282 -12902 2682 -12792
rect 2282 -12962 2292 -12902
rect 2352 -12962 2612 -12902
rect 2672 -12962 2682 -12902
rect 2282 -12972 2682 -12962
rect 2740 -12902 3140 -12792
rect 2740 -12962 2750 -12902
rect 2810 -12962 3070 -12902
rect 3130 -12962 3140 -12902
rect 2740 -12972 3140 -12962
rect 3196 -12902 3596 -12792
rect 3196 -12962 3206 -12902
rect 3266 -12962 3526 -12902
rect 3586 -12962 3596 -12902
rect 3196 -12972 3596 -12962
rect 3652 -12552 4052 -12542
rect 3652 -12612 3662 -12552
rect 3722 -12612 3982 -12552
rect 4042 -12612 4052 -12552
rect 3652 -12722 4052 -12612
rect 4110 -12552 4510 -12542
rect 4110 -12612 4120 -12552
rect 4180 -12612 4440 -12552
rect 4500 -12612 4510 -12552
rect 4110 -12722 4510 -12612
rect 4566 -12552 4966 -12542
rect 4566 -12612 4576 -12552
rect 4636 -12612 4896 -12552
rect 4956 -12612 4966 -12552
rect 4566 -12722 4966 -12612
rect 5022 -12552 5422 -12542
rect 5022 -12612 5032 -12552
rect 5092 -12612 5352 -12552
rect 5412 -12612 5422 -12552
rect 5022 -12722 5422 -12612
rect 5480 -12552 5880 -12542
rect 5480 -12612 5490 -12552
rect 5550 -12612 5810 -12552
rect 5870 -12612 5880 -12552
rect 5480 -12722 5880 -12612
rect 5936 -12552 6336 -12542
rect 5936 -12612 5946 -12552
rect 6006 -12612 6266 -12552
rect 6326 -12612 6336 -12552
rect 5936 -12722 6336 -12612
rect 6392 -12552 6792 -12542
rect 6392 -12612 6402 -12552
rect 6462 -12612 6722 -12552
rect 6782 -12612 6792 -12552
rect 6392 -12722 6792 -12612
rect 6850 -12552 7250 -12542
rect 6850 -12612 6860 -12552
rect 6920 -12612 7180 -12552
rect 7240 -12612 7250 -12552
rect 6850 -12722 7250 -12612
rect 3652 -12792 7250 -12722
rect 3652 -12902 4052 -12792
rect 3652 -12962 3662 -12902
rect 3722 -12962 3982 -12902
rect 4042 -12962 4052 -12902
rect 3652 -12972 4052 -12962
rect 4110 -12902 4510 -12792
rect 4110 -12962 4120 -12902
rect 4180 -12962 4440 -12902
rect 4500 -12962 4510 -12902
rect 4110 -12972 4510 -12962
rect 4566 -12902 4966 -12792
rect 4566 -12962 4576 -12902
rect 4636 -12962 4896 -12902
rect 4956 -12962 4966 -12902
rect 4566 -12972 4966 -12962
rect 5022 -12902 5422 -12792
rect 5022 -12962 5032 -12902
rect 5092 -12962 5352 -12902
rect 5412 -12962 5422 -12902
rect 5022 -12972 5422 -12962
rect 5480 -12902 5880 -12792
rect 5480 -12962 5490 -12902
rect 5550 -12962 5810 -12902
rect 5870 -12962 5880 -12902
rect 5480 -12972 5880 -12962
rect 5936 -12902 6336 -12792
rect 5936 -12962 5946 -12902
rect 6006 -12962 6266 -12902
rect 6326 -12962 6336 -12902
rect 5936 -12972 6336 -12962
rect 6392 -12902 6792 -12792
rect 6392 -12962 6402 -12902
rect 6462 -12962 6722 -12902
rect 6782 -12962 6792 -12902
rect 6392 -12972 6792 -12962
rect 6850 -12902 7250 -12792
rect 6850 -12962 6860 -12902
rect 6920 -12962 7180 -12902
rect 7240 -12962 7250 -12902
rect 6850 -12972 7250 -12962
rect 7306 -12552 7706 -12542
rect 7306 -12612 7316 -12552
rect 7376 -12612 7636 -12552
rect 7696 -12612 7706 -12552
rect 7306 -12722 7706 -12612
rect 7762 -12552 8162 -12542
rect 7762 -12612 7772 -12552
rect 7832 -12612 8092 -12552
rect 8152 -12612 8162 -12552
rect 7762 -12722 8162 -12612
rect 8236 -12552 8636 -12542
rect 8236 -12612 8246 -12552
rect 8306 -12612 8566 -12552
rect 8626 -12612 8636 -12552
rect 8236 -12722 8636 -12612
rect 8692 -12552 9092 -12542
rect 8692 -12612 8702 -12552
rect 8762 -12612 9022 -12552
rect 9082 -12612 9092 -12552
rect 8692 -12722 9092 -12612
rect 9150 -12552 9550 -12542
rect 9150 -12612 9160 -12552
rect 9220 -12612 9480 -12552
rect 9540 -12612 9550 -12552
rect 9150 -12722 9550 -12612
rect 9606 -12552 10006 -12542
rect 9606 -12612 9616 -12552
rect 9676 -12612 9936 -12552
rect 9996 -12612 10006 -12552
rect 9606 -12722 10006 -12612
rect 10062 -12552 10462 -12542
rect 10062 -12612 10072 -12552
rect 10132 -12612 10392 -12552
rect 10452 -12612 10462 -12552
rect 10062 -12722 10462 -12612
rect 10520 -12552 10920 -12542
rect 10520 -12612 10530 -12552
rect 10590 -12612 10850 -12552
rect 10910 -12612 10920 -12552
rect 10520 -12722 10920 -12612
rect 7306 -12792 9093 -12722
rect 9150 -12792 10920 -12722
rect 7306 -12902 7706 -12792
rect 7306 -12962 7316 -12902
rect 7376 -12962 7636 -12902
rect 7696 -12962 7706 -12902
rect 7306 -12972 7706 -12962
rect 7762 -12902 8162 -12792
rect 7762 -12962 7772 -12902
rect 7832 -12962 8092 -12902
rect 8152 -12962 8162 -12902
rect 7762 -12972 8162 -12962
rect 8236 -12902 8636 -12792
rect 8236 -12962 8246 -12902
rect 8306 -12962 8566 -12902
rect 8626 -12962 8636 -12902
rect 8236 -12972 8636 -12962
rect 8692 -12902 9092 -12792
rect 8692 -12962 8702 -12902
rect 8762 -12962 9022 -12902
rect 9082 -12962 9092 -12902
rect 8692 -12972 9092 -12962
rect 9150 -12902 9550 -12792
rect 9150 -12962 9160 -12902
rect 9220 -12962 9480 -12902
rect 9540 -12962 9550 -12902
rect 9150 -12972 9550 -12962
rect 9606 -12902 10006 -12792
rect 9606 -12962 9616 -12902
rect 9676 -12962 9936 -12902
rect 9996 -12962 10006 -12902
rect 9606 -12972 10006 -12962
rect 10062 -12902 10462 -12792
rect 10062 -12962 10072 -12902
rect 10132 -12962 10392 -12902
rect 10452 -12962 10462 -12902
rect 10062 -12972 10462 -12962
rect 10520 -12902 10920 -12792
rect 10520 -12962 10530 -12902
rect 10590 -12962 10850 -12902
rect 10910 -12962 10920 -12902
rect 10520 -12972 10920 -12962
rect 10976 -12552 11376 -12542
rect 10976 -12612 10986 -12552
rect 11046 -12612 11306 -12552
rect 11366 -12612 11376 -12552
rect 10976 -12722 11376 -12612
rect 11432 -12552 11832 -12542
rect 11432 -12612 11442 -12552
rect 11502 -12612 11762 -12552
rect 11822 -12612 11832 -12552
rect 11432 -12722 11832 -12612
rect 11890 -12552 12290 -12542
rect 11890 -12612 11900 -12552
rect 11960 -12612 12220 -12552
rect 12280 -12612 12290 -12552
rect 11890 -12722 12290 -12612
rect 12346 -12552 12746 -12542
rect 12346 -12612 12356 -12552
rect 12416 -12612 12676 -12552
rect 12736 -12612 12746 -12552
rect 12346 -12722 12746 -12612
rect 12802 -12552 13202 -12542
rect 12802 -12612 12812 -12552
rect 12872 -12612 13132 -12552
rect 13192 -12612 13202 -12552
rect 12802 -12722 13202 -12612
rect 13260 -12552 13660 -12542
rect 13260 -12612 13270 -12552
rect 13330 -12612 13590 -12552
rect 13650 -12612 13660 -12552
rect 13260 -12722 13660 -12612
rect 13716 -12552 14116 -12542
rect 13716 -12612 13726 -12552
rect 13786 -12612 14046 -12552
rect 14106 -12612 14116 -12552
rect 13716 -12722 14116 -12612
rect 14172 -12552 14572 -12542
rect 14172 -12612 14182 -12552
rect 14242 -12612 14502 -12552
rect 14562 -12612 14572 -12552
rect 14172 -12722 14572 -12612
rect 14630 -12552 15030 -12542
rect 14630 -12612 14640 -12552
rect 14700 -12612 14960 -12552
rect 15020 -12612 15030 -12552
rect 14630 -12722 15030 -12612
rect 15086 -12552 15486 -12542
rect 15086 -12612 15096 -12552
rect 15156 -12612 15416 -12552
rect 15476 -12612 15486 -12552
rect 15086 -12722 15486 -12612
rect 10976 -12792 15486 -12722
rect 10976 -12902 11376 -12792
rect 10976 -12962 10986 -12902
rect 11046 -12962 11306 -12902
rect 11366 -12962 11376 -12902
rect 10976 -12972 11376 -12962
rect 11432 -12902 11832 -12792
rect 11432 -12962 11442 -12902
rect 11502 -12962 11762 -12902
rect 11822 -12962 11832 -12902
rect 11432 -12972 11832 -12962
rect 11890 -12902 12290 -12792
rect 11890 -12962 11900 -12902
rect 11960 -12962 12220 -12902
rect 12280 -12962 12290 -12902
rect 11890 -12972 12290 -12962
rect 12346 -12902 12746 -12792
rect 12346 -12962 12356 -12902
rect 12416 -12962 12676 -12902
rect 12736 -12962 12746 -12902
rect 12346 -12972 12746 -12962
rect 12802 -12902 13202 -12792
rect 12802 -12962 12812 -12902
rect 12872 -12962 13132 -12902
rect 13192 -12962 13202 -12902
rect 12802 -12972 13202 -12962
rect 13260 -12902 13660 -12792
rect 13260 -12962 13270 -12902
rect 13330 -12962 13590 -12902
rect 13650 -12962 13660 -12902
rect 13260 -12972 13660 -12962
rect 13716 -12902 14116 -12792
rect 13716 -12962 13726 -12902
rect 13786 -12962 14046 -12902
rect 14106 -12962 14116 -12902
rect 13716 -12972 14116 -12962
rect 14172 -12902 14572 -12792
rect 14172 -12962 14182 -12902
rect 14242 -12962 14502 -12902
rect 14562 -12962 14572 -12902
rect 14172 -12972 14572 -12962
rect 14630 -12902 15030 -12792
rect 14630 -12962 14640 -12902
rect 14700 -12962 14960 -12902
rect 15020 -12962 15030 -12902
rect 14630 -12972 15030 -12962
rect 15086 -12902 15486 -12792
rect 15086 -12962 15096 -12902
rect 15156 -12962 15416 -12902
rect 15476 -12962 15486 -12902
rect 15086 -12972 15486 -12962
rect 66 -13044 80 -12972
rect 456 -13044 526 -12972
rect 912 -13044 983 -12972
rect 1370 -13044 1441 -12972
rect 1826 -13044 1897 -12972
rect 2282 -13044 2353 -12972
rect 2740 -13044 2811 -12972
rect 3196 -13044 3267 -12972
rect 3652 -13044 3723 -12972
rect 4110 -13044 4181 -12972
rect 4566 -13044 4637 -12972
rect 5022 -13044 5093 -12972
rect 5480 -13044 5551 -12972
rect 5936 -13044 6007 -12972
rect 6392 -13044 6463 -12972
rect 6850 -13044 6921 -12972
rect 7306 -13044 7377 -12972
rect 7762 -13044 7833 -12972
rect 8236 -13044 8307 -12972
rect 8692 -13044 8763 -12972
rect 9150 -13044 9221 -12972
rect 9606 -13044 9677 -12972
rect 10062 -13044 10133 -12972
rect 10520 -13044 10591 -12972
rect 10976 -13044 11047 -12972
rect 11432 -13044 11503 -12972
rect 11890 -13044 11961 -12972
rect 12346 -13044 12417 -12972
rect 12802 -13044 12873 -12972
rect 13260 -13044 13331 -12972
rect 13716 -13044 13787 -12972
rect 14172 -13044 14243 -12972
rect 14630 -13044 14701 -12972
rect 66 -13054 400 -13044
rect 0 -13114 10 -13054
rect 70 -13114 330 -13054
rect 390 -13114 400 -13054
rect 0 -13404 14 -13114
rect 66 -13404 400 -13114
rect 0 -13464 10 -13404
rect 70 -13464 330 -13404
rect 390 -13464 400 -13404
rect 0 -13546 14 -13464
rect 66 -13474 400 -13464
rect 456 -13054 856 -13044
rect 456 -13114 466 -13054
rect 526 -13114 786 -13054
rect 846 -13114 856 -13054
rect 456 -13224 856 -13114
rect 912 -13054 1312 -13044
rect 912 -13114 922 -13054
rect 982 -13114 1242 -13054
rect 1302 -13114 1312 -13054
rect 912 -13224 1312 -13114
rect 1370 -13054 1770 -13044
rect 1370 -13114 1380 -13054
rect 1440 -13114 1700 -13054
rect 1760 -13114 1770 -13054
rect 1370 -13224 1770 -13114
rect 1826 -13054 2226 -13044
rect 1826 -13114 1836 -13054
rect 1896 -13114 2156 -13054
rect 2216 -13114 2226 -13054
rect 1826 -13224 2226 -13114
rect 2282 -13054 2682 -13044
rect 2282 -13114 2292 -13054
rect 2352 -13114 2612 -13054
rect 2672 -13114 2682 -13054
rect 2282 -13224 2682 -13114
rect 2740 -13054 3140 -13044
rect 2740 -13114 2750 -13054
rect 2810 -13114 3070 -13054
rect 3130 -13114 3140 -13054
rect 2740 -13224 3140 -13114
rect 3196 -13054 3596 -13044
rect 3196 -13114 3206 -13054
rect 3266 -13114 3526 -13054
rect 3586 -13114 3596 -13054
rect 3196 -13224 3596 -13114
rect 456 -13294 3596 -13224
rect 456 -13404 856 -13294
rect 456 -13464 466 -13404
rect 526 -13464 786 -13404
rect 846 -13464 856 -13404
rect 456 -13474 856 -13464
rect 912 -13404 1312 -13294
rect 912 -13464 922 -13404
rect 982 -13464 1242 -13404
rect 1302 -13464 1312 -13404
rect 912 -13474 1312 -13464
rect 1370 -13404 1770 -13294
rect 1370 -13464 1380 -13404
rect 1440 -13464 1700 -13404
rect 1760 -13464 1770 -13404
rect 1370 -13474 1770 -13464
rect 1826 -13404 2226 -13294
rect 1826 -13464 1836 -13404
rect 1896 -13464 2156 -13404
rect 2216 -13464 2226 -13404
rect 1826 -13474 2226 -13464
rect 2282 -13404 2682 -13294
rect 2282 -13464 2292 -13404
rect 2352 -13464 2612 -13404
rect 2672 -13464 2682 -13404
rect 2282 -13474 2682 -13464
rect 2740 -13404 3140 -13294
rect 2740 -13464 2750 -13404
rect 2810 -13464 3070 -13404
rect 3130 -13464 3140 -13404
rect 2740 -13474 3140 -13464
rect 3196 -13404 3596 -13294
rect 3196 -13464 3206 -13404
rect 3266 -13464 3526 -13404
rect 3586 -13464 3596 -13404
rect 3196 -13474 3596 -13464
rect 3652 -13054 4052 -13044
rect 3652 -13114 3662 -13054
rect 3722 -13114 3982 -13054
rect 4042 -13114 4052 -13054
rect 3652 -13224 4052 -13114
rect 4110 -13054 4510 -13044
rect 4110 -13114 4120 -13054
rect 4180 -13114 4440 -13054
rect 4500 -13114 4510 -13054
rect 4110 -13224 4510 -13114
rect 4566 -13054 4966 -13044
rect 4566 -13114 4576 -13054
rect 4636 -13114 4896 -13054
rect 4956 -13114 4966 -13054
rect 4566 -13224 4966 -13114
rect 5022 -13054 5422 -13044
rect 5022 -13114 5032 -13054
rect 5092 -13114 5352 -13054
rect 5412 -13114 5422 -13054
rect 5022 -13224 5422 -13114
rect 5480 -13054 5880 -13044
rect 5480 -13114 5490 -13054
rect 5550 -13114 5810 -13054
rect 5870 -13114 5880 -13054
rect 5480 -13224 5880 -13114
rect 5936 -13054 6336 -13044
rect 5936 -13114 5946 -13054
rect 6006 -13114 6266 -13054
rect 6326 -13114 6336 -13054
rect 5936 -13224 6336 -13114
rect 6392 -13054 6792 -13044
rect 6392 -13114 6402 -13054
rect 6462 -13114 6722 -13054
rect 6782 -13114 6792 -13054
rect 6392 -13224 6792 -13114
rect 6850 -13054 7250 -13044
rect 6850 -13114 6860 -13054
rect 6920 -13114 7180 -13054
rect 7240 -13114 7250 -13054
rect 6850 -13224 7250 -13114
rect 3652 -13294 7250 -13224
rect 3652 -13404 4052 -13294
rect 3652 -13464 3662 -13404
rect 3722 -13464 3982 -13404
rect 4042 -13464 4052 -13404
rect 3652 -13474 4052 -13464
rect 4110 -13404 4510 -13294
rect 4110 -13464 4120 -13404
rect 4180 -13464 4440 -13404
rect 4500 -13464 4510 -13404
rect 4110 -13474 4510 -13464
rect 4566 -13404 4966 -13294
rect 4566 -13464 4576 -13404
rect 4636 -13464 4896 -13404
rect 4956 -13464 4966 -13404
rect 4566 -13474 4966 -13464
rect 5022 -13404 5422 -13294
rect 5022 -13464 5032 -13404
rect 5092 -13464 5352 -13404
rect 5412 -13464 5422 -13404
rect 5022 -13474 5422 -13464
rect 5480 -13404 5880 -13294
rect 5480 -13464 5490 -13404
rect 5550 -13464 5810 -13404
rect 5870 -13464 5880 -13404
rect 5480 -13474 5880 -13464
rect 5936 -13404 6336 -13294
rect 5936 -13464 5946 -13404
rect 6006 -13464 6266 -13404
rect 6326 -13464 6336 -13404
rect 5936 -13474 6336 -13464
rect 6392 -13404 6792 -13294
rect 6392 -13464 6402 -13404
rect 6462 -13464 6722 -13404
rect 6782 -13464 6792 -13404
rect 6392 -13474 6792 -13464
rect 6850 -13404 7250 -13294
rect 6850 -13464 6860 -13404
rect 6920 -13464 7180 -13404
rect 7240 -13464 7250 -13404
rect 6850 -13474 7250 -13464
rect 7306 -13054 7706 -13044
rect 7306 -13114 7316 -13054
rect 7376 -13114 7636 -13054
rect 7696 -13114 7706 -13054
rect 7306 -13224 7706 -13114
rect 7762 -13054 8162 -13044
rect 7762 -13114 7772 -13054
rect 7832 -13114 8092 -13054
rect 8152 -13114 8162 -13054
rect 7762 -13224 8162 -13114
rect 8236 -13054 8636 -13044
rect 8236 -13114 8246 -13054
rect 8306 -13114 8566 -13054
rect 8626 -13114 8636 -13054
rect 8236 -13224 8636 -13114
rect 8692 -13054 9092 -13044
rect 8692 -13114 8702 -13054
rect 8762 -13114 9022 -13054
rect 9082 -13114 9092 -13054
rect 8692 -13224 9092 -13114
rect 9150 -13054 9550 -13044
rect 9150 -13114 9160 -13054
rect 9220 -13114 9480 -13054
rect 9540 -13114 9550 -13054
rect 9150 -13224 9550 -13114
rect 9606 -13054 10006 -13044
rect 9606 -13114 9616 -13054
rect 9676 -13114 9936 -13054
rect 9996 -13114 10006 -13054
rect 9606 -13224 10006 -13114
rect 10062 -13054 10462 -13044
rect 10062 -13114 10072 -13054
rect 10132 -13114 10392 -13054
rect 10452 -13114 10462 -13054
rect 10062 -13224 10462 -13114
rect 10520 -13054 10920 -13044
rect 10520 -13114 10530 -13054
rect 10590 -13114 10850 -13054
rect 10910 -13114 10920 -13054
rect 10520 -13224 10920 -13114
rect 7306 -13294 9093 -13224
rect 9150 -13294 10920 -13224
rect 7306 -13404 7706 -13294
rect 7306 -13464 7316 -13404
rect 7376 -13464 7636 -13404
rect 7696 -13464 7706 -13404
rect 7306 -13474 7706 -13464
rect 7762 -13404 8162 -13294
rect 7762 -13464 7772 -13404
rect 7832 -13464 8092 -13404
rect 8152 -13464 8162 -13404
rect 7762 -13474 8162 -13464
rect 8236 -13404 8636 -13294
rect 8236 -13464 8246 -13404
rect 8306 -13464 8566 -13404
rect 8626 -13464 8636 -13404
rect 8236 -13474 8636 -13464
rect 8692 -13404 9092 -13294
rect 8692 -13464 8702 -13404
rect 8762 -13464 9022 -13404
rect 9082 -13464 9092 -13404
rect 8692 -13474 9092 -13464
rect 9150 -13404 9550 -13294
rect 9150 -13464 9160 -13404
rect 9220 -13464 9480 -13404
rect 9540 -13464 9550 -13404
rect 9150 -13474 9550 -13464
rect 9606 -13404 10006 -13294
rect 9606 -13464 9616 -13404
rect 9676 -13464 9936 -13404
rect 9996 -13464 10006 -13404
rect 9606 -13474 10006 -13464
rect 10062 -13404 10462 -13294
rect 10062 -13464 10072 -13404
rect 10132 -13464 10392 -13404
rect 10452 -13464 10462 -13404
rect 10062 -13474 10462 -13464
rect 10520 -13404 10920 -13294
rect 10520 -13464 10530 -13404
rect 10590 -13464 10850 -13404
rect 10910 -13464 10920 -13404
rect 10520 -13474 10920 -13464
rect 10976 -13054 11376 -13044
rect 10976 -13114 10986 -13054
rect 11046 -13114 11306 -13054
rect 11366 -13114 11376 -13054
rect 10976 -13224 11376 -13114
rect 11432 -13054 11832 -13044
rect 11432 -13114 11442 -13054
rect 11502 -13114 11762 -13054
rect 11822 -13114 11832 -13054
rect 11432 -13224 11832 -13114
rect 11890 -13054 12290 -13044
rect 11890 -13114 11900 -13054
rect 11960 -13114 12220 -13054
rect 12280 -13114 12290 -13054
rect 11890 -13224 12290 -13114
rect 12346 -13054 12746 -13044
rect 12346 -13114 12356 -13054
rect 12416 -13114 12676 -13054
rect 12736 -13114 12746 -13054
rect 12346 -13224 12746 -13114
rect 12802 -13054 13202 -13044
rect 12802 -13114 12812 -13054
rect 12872 -13114 13132 -13054
rect 13192 -13114 13202 -13054
rect 12802 -13224 13202 -13114
rect 13260 -13054 13660 -13044
rect 13260 -13114 13270 -13054
rect 13330 -13114 13590 -13054
rect 13650 -13114 13660 -13054
rect 13260 -13224 13660 -13114
rect 13716 -13054 14116 -13044
rect 13716 -13114 13726 -13054
rect 13786 -13114 14046 -13054
rect 14106 -13114 14116 -13054
rect 13716 -13224 14116 -13114
rect 14172 -13054 14572 -13044
rect 14172 -13114 14182 -13054
rect 14242 -13114 14502 -13054
rect 14562 -13114 14572 -13054
rect 14172 -13224 14572 -13114
rect 14630 -13054 15030 -13044
rect 14630 -13114 14640 -13054
rect 14700 -13114 14960 -13054
rect 15020 -13114 15030 -13054
rect 14630 -13224 15030 -13114
rect 15086 -13054 15486 -13044
rect 15086 -13114 15096 -13054
rect 15156 -13114 15416 -13054
rect 15476 -13114 15486 -13054
rect 15086 -13224 15486 -13114
rect 10976 -13294 15486 -13224
rect 10976 -13404 11376 -13294
rect 10976 -13464 10986 -13404
rect 11046 -13464 11306 -13404
rect 11366 -13464 11376 -13404
rect 10976 -13474 11376 -13464
rect 11432 -13404 11832 -13294
rect 11432 -13464 11442 -13404
rect 11502 -13464 11762 -13404
rect 11822 -13464 11832 -13404
rect 11432 -13474 11832 -13464
rect 11890 -13404 12290 -13294
rect 11890 -13464 11900 -13404
rect 11960 -13464 12220 -13404
rect 12280 -13464 12290 -13404
rect 11890 -13474 12290 -13464
rect 12346 -13404 12746 -13294
rect 12346 -13464 12356 -13404
rect 12416 -13464 12676 -13404
rect 12736 -13464 12746 -13404
rect 12346 -13474 12746 -13464
rect 12802 -13404 13202 -13294
rect 12802 -13464 12812 -13404
rect 12872 -13464 13132 -13404
rect 13192 -13464 13202 -13404
rect 12802 -13474 13202 -13464
rect 13260 -13404 13660 -13294
rect 13260 -13464 13270 -13404
rect 13330 -13464 13590 -13404
rect 13650 -13464 13660 -13404
rect 13260 -13474 13660 -13464
rect 13716 -13404 14116 -13294
rect 13716 -13464 13726 -13404
rect 13786 -13464 14046 -13404
rect 14106 -13464 14116 -13404
rect 13716 -13474 14116 -13464
rect 14172 -13404 14572 -13294
rect 14172 -13464 14182 -13404
rect 14242 -13464 14502 -13404
rect 14562 -13464 14572 -13404
rect 14172 -13474 14572 -13464
rect 14630 -13404 15030 -13294
rect 14630 -13464 14640 -13404
rect 14700 -13464 14960 -13404
rect 15020 -13464 15030 -13404
rect 14630 -13474 15030 -13464
rect 15086 -13404 15486 -13294
rect 15086 -13464 15096 -13404
rect 15156 -13464 15416 -13404
rect 15476 -13464 15486 -13404
rect 15086 -13474 15486 -13464
rect 66 -13536 80 -13474
rect 456 -13536 527 -13474
rect 912 -13536 983 -13474
rect 1370 -13536 1441 -13474
rect 1826 -13536 1897 -13474
rect 2282 -13536 2353 -13474
rect 2740 -13536 2810 -13474
rect 3196 -13536 3266 -13474
rect 3652 -13536 3722 -13474
rect 4110 -13536 4180 -13474
rect 4566 -13536 4636 -13474
rect 5022 -13536 5092 -13474
rect 5480 -13536 5550 -13474
rect 5936 -13536 6006 -13474
rect 6392 -13536 6462 -13474
rect 6850 -13536 6920 -13474
rect 7306 -13536 7376 -13474
rect 7762 -13536 7832 -13474
rect 8236 -13536 8306 -13474
rect 8692 -13536 8762 -13474
rect 9150 -13536 9220 -13474
rect 9606 -13536 9676 -13474
rect 10062 -13536 10132 -13474
rect 10520 -13536 10590 -13474
rect 10976 -13536 11046 -13474
rect 11432 -13536 11502 -13474
rect 11890 -13536 11960 -13474
rect 66 -13546 400 -13536
rect 0 -13606 10 -13546
rect 70 -13606 330 -13546
rect 390 -13606 400 -13546
rect 0 -13896 14 -13606
rect 66 -13896 400 -13606
rect 0 -13956 10 -13896
rect 70 -13956 330 -13896
rect 390 -13956 400 -13896
rect 0 -14040 14 -13956
rect 66 -13966 400 -13956
rect 456 -13546 856 -13536
rect 456 -13606 466 -13546
rect 526 -13606 786 -13546
rect 846 -13606 856 -13546
rect 456 -13716 856 -13606
rect 912 -13546 1312 -13536
rect 912 -13606 922 -13546
rect 982 -13606 1242 -13546
rect 1302 -13606 1312 -13546
rect 912 -13716 1312 -13606
rect 1370 -13546 1770 -13536
rect 1370 -13606 1380 -13546
rect 1440 -13606 1700 -13546
rect 1760 -13606 1770 -13546
rect 1370 -13716 1770 -13606
rect 1826 -13546 2226 -13536
rect 1826 -13606 1836 -13546
rect 1896 -13606 2156 -13546
rect 2216 -13606 2226 -13546
rect 1826 -13716 2226 -13606
rect 2282 -13546 2682 -13536
rect 2282 -13606 2292 -13546
rect 2352 -13606 2612 -13546
rect 2672 -13606 2682 -13546
rect 2282 -13716 2682 -13606
rect 2740 -13546 3140 -13536
rect 2740 -13606 2750 -13546
rect 2810 -13606 3070 -13546
rect 3130 -13606 3140 -13546
rect 2740 -13716 3140 -13606
rect 3196 -13546 3596 -13536
rect 3196 -13606 3206 -13546
rect 3266 -13606 3526 -13546
rect 3586 -13606 3596 -13546
rect 3196 -13716 3596 -13606
rect 456 -13786 3596 -13716
rect 456 -13896 856 -13786
rect 456 -13956 466 -13896
rect 526 -13956 786 -13896
rect 846 -13956 856 -13896
rect 456 -13966 856 -13956
rect 912 -13896 1312 -13786
rect 912 -13956 922 -13896
rect 982 -13956 1242 -13896
rect 1302 -13956 1312 -13896
rect 912 -13966 1312 -13956
rect 1370 -13896 1770 -13786
rect 1370 -13956 1380 -13896
rect 1440 -13956 1700 -13896
rect 1760 -13956 1770 -13896
rect 1370 -13966 1770 -13956
rect 1826 -13896 2226 -13786
rect 1826 -13956 1836 -13896
rect 1896 -13956 2156 -13896
rect 2216 -13956 2226 -13896
rect 1826 -13966 2226 -13956
rect 2282 -13896 2682 -13786
rect 2282 -13956 2292 -13896
rect 2352 -13956 2612 -13896
rect 2672 -13956 2682 -13896
rect 2282 -13966 2682 -13956
rect 2740 -13896 3140 -13786
rect 2740 -13956 2750 -13896
rect 2810 -13956 3070 -13896
rect 3130 -13956 3140 -13896
rect 2740 -13966 3140 -13956
rect 3196 -13896 3596 -13786
rect 3196 -13956 3206 -13896
rect 3266 -13956 3526 -13896
rect 3586 -13956 3596 -13896
rect 3196 -13966 3596 -13956
rect 3652 -13546 4052 -13536
rect 3652 -13606 3662 -13546
rect 3722 -13606 3982 -13546
rect 4042 -13606 4052 -13546
rect 3652 -13716 4052 -13606
rect 4110 -13546 4510 -13536
rect 4110 -13606 4120 -13546
rect 4180 -13606 4440 -13546
rect 4500 -13606 4510 -13546
rect 4110 -13716 4510 -13606
rect 4566 -13546 4966 -13536
rect 4566 -13606 4576 -13546
rect 4636 -13606 4896 -13546
rect 4956 -13606 4966 -13546
rect 4566 -13716 4966 -13606
rect 5022 -13546 5422 -13536
rect 5022 -13606 5032 -13546
rect 5092 -13606 5352 -13546
rect 5412 -13606 5422 -13546
rect 5022 -13716 5422 -13606
rect 5480 -13546 5880 -13536
rect 5480 -13606 5490 -13546
rect 5550 -13606 5810 -13546
rect 5870 -13606 5880 -13546
rect 5480 -13716 5880 -13606
rect 5936 -13546 6336 -13536
rect 5936 -13606 5946 -13546
rect 6006 -13606 6266 -13546
rect 6326 -13606 6336 -13546
rect 5936 -13716 6336 -13606
rect 6392 -13546 6792 -13536
rect 6392 -13606 6402 -13546
rect 6462 -13606 6722 -13546
rect 6782 -13606 6792 -13546
rect 6392 -13716 6792 -13606
rect 6850 -13546 7250 -13536
rect 6850 -13606 6860 -13546
rect 6920 -13606 7180 -13546
rect 7240 -13606 7250 -13546
rect 6850 -13716 7250 -13606
rect 3652 -13786 7250 -13716
rect 3652 -13896 4052 -13786
rect 3652 -13956 3662 -13896
rect 3722 -13956 3982 -13896
rect 4042 -13956 4052 -13896
rect 3652 -13966 4052 -13956
rect 4110 -13896 4510 -13786
rect 4110 -13956 4120 -13896
rect 4180 -13956 4440 -13896
rect 4500 -13956 4510 -13896
rect 4110 -13966 4510 -13956
rect 4566 -13896 4966 -13786
rect 4566 -13956 4576 -13896
rect 4636 -13956 4896 -13896
rect 4956 -13956 4966 -13896
rect 4566 -13966 4966 -13956
rect 5022 -13896 5422 -13786
rect 5022 -13956 5032 -13896
rect 5092 -13956 5352 -13896
rect 5412 -13956 5422 -13896
rect 5022 -13966 5422 -13956
rect 5480 -13896 5880 -13786
rect 5480 -13956 5490 -13896
rect 5550 -13956 5810 -13896
rect 5870 -13956 5880 -13896
rect 5480 -13966 5880 -13956
rect 5936 -13896 6336 -13786
rect 5936 -13956 5946 -13896
rect 6006 -13956 6266 -13896
rect 6326 -13956 6336 -13896
rect 5936 -13966 6336 -13956
rect 6392 -13896 6792 -13786
rect 6392 -13956 6402 -13896
rect 6462 -13956 6722 -13896
rect 6782 -13956 6792 -13896
rect 6392 -13966 6792 -13956
rect 6850 -13896 7250 -13786
rect 6850 -13956 6860 -13896
rect 6920 -13956 7180 -13896
rect 7240 -13956 7250 -13896
rect 6850 -13966 7250 -13956
rect 7306 -13546 7706 -13536
rect 7306 -13606 7316 -13546
rect 7376 -13606 7636 -13546
rect 7696 -13606 7706 -13546
rect 7306 -13716 7706 -13606
rect 7762 -13546 8162 -13536
rect 7762 -13606 7772 -13546
rect 7832 -13606 8092 -13546
rect 8152 -13606 8162 -13546
rect 7762 -13716 8162 -13606
rect 8236 -13546 8636 -13536
rect 8236 -13606 8246 -13546
rect 8306 -13606 8566 -13546
rect 8626 -13606 8636 -13546
rect 8236 -13716 8636 -13606
rect 8692 -13546 9092 -13536
rect 8692 -13606 8702 -13546
rect 8762 -13606 9022 -13546
rect 9082 -13606 9092 -13546
rect 8692 -13716 9092 -13606
rect 9150 -13546 9550 -13536
rect 9150 -13606 9160 -13546
rect 9220 -13606 9480 -13546
rect 9540 -13606 9550 -13546
rect 9150 -13716 9550 -13606
rect 9606 -13546 10006 -13536
rect 9606 -13606 9616 -13546
rect 9676 -13606 9936 -13546
rect 9996 -13606 10006 -13546
rect 9606 -13716 10006 -13606
rect 10062 -13546 10462 -13536
rect 10062 -13606 10072 -13546
rect 10132 -13606 10392 -13546
rect 10452 -13606 10462 -13546
rect 10062 -13716 10462 -13606
rect 10520 -13546 10920 -13536
rect 10520 -13606 10530 -13546
rect 10590 -13606 10850 -13546
rect 10910 -13606 10920 -13546
rect 10520 -13716 10920 -13606
rect 7306 -13786 9093 -13716
rect 9150 -13786 10920 -13716
rect 7306 -13896 7706 -13786
rect 7306 -13956 7316 -13896
rect 7376 -13956 7636 -13896
rect 7696 -13956 7706 -13896
rect 7306 -13966 7706 -13956
rect 7762 -13896 8162 -13786
rect 7762 -13956 7772 -13896
rect 7832 -13956 8092 -13896
rect 8152 -13956 8162 -13896
rect 7762 -13966 8162 -13956
rect 8236 -13896 8636 -13786
rect 8236 -13956 8246 -13896
rect 8306 -13956 8566 -13896
rect 8626 -13956 8636 -13896
rect 8236 -13966 8636 -13956
rect 8692 -13896 9092 -13786
rect 8692 -13956 8702 -13896
rect 8762 -13956 9022 -13896
rect 9082 -13956 9092 -13896
rect 8692 -13966 9092 -13956
rect 9150 -13896 9550 -13786
rect 9150 -13956 9160 -13896
rect 9220 -13956 9480 -13896
rect 9540 -13956 9550 -13896
rect 9150 -13966 9550 -13956
rect 9606 -13896 10006 -13786
rect 9606 -13956 9616 -13896
rect 9676 -13956 9936 -13896
rect 9996 -13956 10006 -13896
rect 9606 -13966 10006 -13956
rect 10062 -13896 10462 -13786
rect 10062 -13956 10072 -13896
rect 10132 -13956 10392 -13896
rect 10452 -13956 10462 -13896
rect 10062 -13966 10462 -13956
rect 10520 -13896 10920 -13786
rect 10520 -13956 10530 -13896
rect 10590 -13956 10850 -13896
rect 10910 -13956 10920 -13896
rect 10520 -13966 10920 -13956
rect 10976 -13546 11376 -13536
rect 10976 -13606 10986 -13546
rect 11046 -13606 11306 -13546
rect 11366 -13606 11376 -13546
rect 10976 -13716 11376 -13606
rect 11432 -13546 11832 -13536
rect 11432 -13606 11442 -13546
rect 11502 -13606 11762 -13546
rect 11822 -13606 11832 -13546
rect 11432 -13716 11832 -13606
rect 11890 -13546 12290 -13536
rect 11890 -13606 11900 -13546
rect 11960 -13606 12220 -13546
rect 12280 -13606 12290 -13546
rect 11890 -13716 12290 -13606
rect 10976 -13786 12290 -13716
rect 10976 -13896 11376 -13786
rect 10976 -13956 10986 -13896
rect 11046 -13956 11306 -13896
rect 11366 -13956 11376 -13896
rect 10976 -13966 11376 -13956
rect 11432 -13896 11832 -13786
rect 11432 -13956 11442 -13896
rect 11502 -13956 11762 -13896
rect 11822 -13956 11832 -13896
rect 11432 -13966 11832 -13956
rect 11890 -13896 12290 -13786
rect 11890 -13956 11900 -13896
rect 11960 -13956 12220 -13896
rect 12280 -13956 12290 -13896
rect 11890 -13966 12290 -13956
rect 12346 -13546 12746 -13536
rect 12346 -13606 12356 -13546
rect 12416 -13606 12676 -13546
rect 12736 -13606 12746 -13546
rect 12346 -13716 12746 -13606
rect 12802 -13546 13202 -13536
rect 12802 -13606 12812 -13546
rect 12872 -13606 13132 -13546
rect 13192 -13606 13202 -13546
rect 12802 -13716 13202 -13606
rect 13260 -13546 13660 -13536
rect 13260 -13606 13270 -13546
rect 13330 -13606 13590 -13546
rect 13650 -13606 13660 -13546
rect 13260 -13716 13660 -13606
rect 13716 -13546 14116 -13536
rect 13716 -13606 13726 -13546
rect 13786 -13606 14046 -13546
rect 14106 -13606 14116 -13546
rect 13716 -13716 14116 -13606
rect 14172 -13546 14572 -13536
rect 14172 -13606 14182 -13546
rect 14242 -13606 14502 -13546
rect 14562 -13606 14572 -13546
rect 14172 -13716 14572 -13606
rect 14630 -13546 15030 -13536
rect 14630 -13606 14640 -13546
rect 14700 -13606 14960 -13546
rect 15020 -13606 15030 -13546
rect 14630 -13716 15030 -13606
rect 15086 -13546 15486 -13536
rect 15086 -13606 15096 -13546
rect 15156 -13606 15416 -13546
rect 15476 -13606 15486 -13546
rect 15086 -13716 15486 -13606
rect 12346 -13786 15486 -13716
rect 12346 -13896 12746 -13786
rect 12346 -13956 12356 -13896
rect 12416 -13956 12676 -13896
rect 12736 -13956 12746 -13896
rect 12346 -13966 12746 -13956
rect 12802 -13896 13202 -13786
rect 12802 -13956 12812 -13896
rect 12872 -13956 13132 -13896
rect 13192 -13956 13202 -13896
rect 12802 -13966 13202 -13956
rect 13260 -13896 13660 -13786
rect 13260 -13956 13270 -13896
rect 13330 -13956 13590 -13896
rect 13650 -13956 13660 -13896
rect 13260 -13966 13660 -13956
rect 13716 -13896 14116 -13786
rect 13716 -13956 13726 -13896
rect 13786 -13956 14046 -13896
rect 14106 -13956 14116 -13896
rect 13716 -13966 14116 -13956
rect 14172 -13896 14572 -13786
rect 14172 -13956 14182 -13896
rect 14242 -13956 14502 -13896
rect 14562 -13956 14572 -13896
rect 14172 -13966 14572 -13956
rect 14630 -13896 15030 -13786
rect 14630 -13956 14640 -13896
rect 14700 -13956 14960 -13896
rect 15020 -13956 15030 -13896
rect 14630 -13966 15030 -13956
rect 15086 -13896 15486 -13786
rect 15086 -13956 15096 -13896
rect 15156 -13956 15416 -13896
rect 15476 -13956 15486 -13896
rect 15086 -13966 15486 -13956
rect 66 -14030 80 -13966
rect 456 -14030 526 -13966
rect 912 -14030 982 -13966
rect 1370 -14030 1440 -13966
rect 1826 -14030 1896 -13966
rect 2282 -14030 2352 -13966
rect 2740 -14030 2810 -13966
rect 3196 -14030 3266 -13966
rect 3652 -14030 3722 -13966
rect 4110 -14030 4180 -13966
rect 4566 -14030 4636 -13966
rect 5022 -14030 5092 -13966
rect 5480 -14030 5550 -13966
rect 5936 -14030 6006 -13966
rect 6392 -14030 6462 -13966
rect 6850 -14030 6920 -13966
rect 7306 -14030 7376 -13966
rect 7762 -14030 7832 -13966
rect 8236 -14030 8306 -13966
rect 8692 -14030 8762 -13966
rect 9150 -14030 9220 -13966
rect 9606 -14030 9676 -13966
rect 10062 -14030 10132 -13966
rect 10520 -14030 10590 -13966
rect 10976 -14030 11047 -13966
rect 11432 -14030 11503 -13966
rect 11890 -14030 11961 -13966
rect 12346 -14030 12417 -13966
rect 12802 -14030 12873 -13966
rect 66 -14040 400 -14030
rect 0 -14100 10 -14040
rect 70 -14100 330 -14040
rect 390 -14100 400 -14040
rect 0 -14390 14 -14100
rect 66 -14390 400 -14100
rect 0 -14450 10 -14390
rect 70 -14450 330 -14390
rect 390 -14450 400 -14390
rect 0 -14542 14 -14450
rect 66 -14460 400 -14450
rect 456 -14040 856 -14030
rect 456 -14100 466 -14040
rect 526 -14100 786 -14040
rect 846 -14100 856 -14040
rect 456 -14209 856 -14100
rect 912 -14040 1312 -14030
rect 912 -14100 922 -14040
rect 982 -14100 1242 -14040
rect 1302 -14100 1312 -14040
rect 912 -14209 1312 -14100
rect 1370 -14040 1770 -14030
rect 1370 -14100 1380 -14040
rect 1440 -14100 1700 -14040
rect 1760 -14100 1770 -14040
rect 1370 -14209 1770 -14100
rect 1826 -14040 2226 -14030
rect 1826 -14100 1836 -14040
rect 1896 -14100 2156 -14040
rect 2216 -14100 2226 -14040
rect 1826 -14209 2226 -14100
rect 2282 -14040 2682 -14030
rect 2282 -14100 2292 -14040
rect 2352 -14100 2612 -14040
rect 2672 -14100 2682 -14040
rect 2282 -14209 2682 -14100
rect 2740 -14040 3140 -14030
rect 2740 -14100 2750 -14040
rect 2810 -14100 3070 -14040
rect 3130 -14100 3140 -14040
rect 2740 -14209 3140 -14100
rect 3196 -14040 3596 -14030
rect 3196 -14100 3206 -14040
rect 3266 -14100 3526 -14040
rect 3586 -14100 3596 -14040
rect 3196 -14209 3596 -14100
rect 456 -14279 3596 -14209
rect 456 -14390 856 -14279
rect 456 -14450 466 -14390
rect 526 -14450 786 -14390
rect 846 -14450 856 -14390
rect 456 -14460 856 -14450
rect 912 -14390 1312 -14279
rect 912 -14450 922 -14390
rect 982 -14450 1242 -14390
rect 1302 -14450 1312 -14390
rect 912 -14460 1312 -14450
rect 1370 -14390 1770 -14279
rect 1370 -14450 1380 -14390
rect 1440 -14450 1700 -14390
rect 1760 -14450 1770 -14390
rect 1370 -14460 1770 -14450
rect 1826 -14390 2226 -14279
rect 1826 -14450 1836 -14390
rect 1896 -14450 2156 -14390
rect 2216 -14450 2226 -14390
rect 1826 -14460 2226 -14450
rect 2282 -14390 2682 -14279
rect 2282 -14450 2292 -14390
rect 2352 -14450 2612 -14390
rect 2672 -14450 2682 -14390
rect 2282 -14460 2682 -14450
rect 2740 -14390 3140 -14279
rect 2740 -14450 2750 -14390
rect 2810 -14450 3070 -14390
rect 3130 -14450 3140 -14390
rect 2740 -14460 3140 -14450
rect 3196 -14390 3596 -14279
rect 3196 -14450 3206 -14390
rect 3266 -14450 3526 -14390
rect 3586 -14450 3596 -14390
rect 3196 -14460 3596 -14450
rect 3652 -14040 4052 -14030
rect 3652 -14100 3662 -14040
rect 3722 -14100 3982 -14040
rect 4042 -14100 4052 -14040
rect 3652 -14209 4052 -14100
rect 4110 -14040 4510 -14030
rect 4110 -14100 4120 -14040
rect 4180 -14100 4440 -14040
rect 4500 -14100 4510 -14040
rect 4110 -14209 4510 -14100
rect 4566 -14040 4966 -14030
rect 4566 -14100 4576 -14040
rect 4636 -14100 4896 -14040
rect 4956 -14100 4966 -14040
rect 4566 -14209 4966 -14100
rect 5022 -14040 5422 -14030
rect 5022 -14100 5032 -14040
rect 5092 -14100 5352 -14040
rect 5412 -14100 5422 -14040
rect 5022 -14209 5422 -14100
rect 5480 -14040 5880 -14030
rect 5480 -14100 5490 -14040
rect 5550 -14100 5810 -14040
rect 5870 -14100 5880 -14040
rect 5480 -14209 5880 -14100
rect 5936 -14040 6336 -14030
rect 5936 -14100 5946 -14040
rect 6006 -14100 6266 -14040
rect 6326 -14100 6336 -14040
rect 5936 -14209 6336 -14100
rect 6392 -14040 6792 -14030
rect 6392 -14100 6402 -14040
rect 6462 -14100 6722 -14040
rect 6782 -14100 6792 -14040
rect 6392 -14209 6792 -14100
rect 6850 -14040 7250 -14030
rect 6850 -14100 6860 -14040
rect 6920 -14100 7180 -14040
rect 7240 -14100 7250 -14040
rect 6850 -14209 7250 -14100
rect 3652 -14279 7250 -14209
rect 3652 -14390 4052 -14279
rect 3652 -14450 3662 -14390
rect 3722 -14450 3982 -14390
rect 4042 -14450 4052 -14390
rect 3652 -14460 4052 -14450
rect 4110 -14390 4510 -14279
rect 4110 -14450 4120 -14390
rect 4180 -14450 4440 -14390
rect 4500 -14450 4510 -14390
rect 4110 -14460 4510 -14450
rect 4566 -14390 4966 -14279
rect 4566 -14450 4576 -14390
rect 4636 -14450 4896 -14390
rect 4956 -14450 4966 -14390
rect 4566 -14460 4966 -14450
rect 5022 -14390 5422 -14279
rect 5022 -14450 5032 -14390
rect 5092 -14450 5352 -14390
rect 5412 -14450 5422 -14390
rect 5022 -14460 5422 -14450
rect 5480 -14390 5880 -14279
rect 5480 -14450 5490 -14390
rect 5550 -14450 5810 -14390
rect 5870 -14450 5880 -14390
rect 5480 -14460 5880 -14450
rect 5936 -14390 6336 -14279
rect 5936 -14450 5946 -14390
rect 6006 -14450 6266 -14390
rect 6326 -14450 6336 -14390
rect 5936 -14460 6336 -14450
rect 6392 -14390 6792 -14279
rect 6392 -14450 6402 -14390
rect 6462 -14450 6722 -14390
rect 6782 -14450 6792 -14390
rect 6392 -14460 6792 -14450
rect 6850 -14390 7250 -14279
rect 6850 -14450 6860 -14390
rect 6920 -14450 7180 -14390
rect 7240 -14450 7250 -14390
rect 6850 -14460 7250 -14450
rect 7306 -14040 7706 -14030
rect 7306 -14100 7316 -14040
rect 7376 -14100 7636 -14040
rect 7696 -14100 7706 -14040
rect 7306 -14209 7706 -14100
rect 7762 -14040 8162 -14030
rect 7762 -14100 7772 -14040
rect 7832 -14100 8092 -14040
rect 8152 -14100 8162 -14040
rect 7762 -14209 8162 -14100
rect 8236 -14040 8636 -14030
rect 8236 -14100 8246 -14040
rect 8306 -14100 8566 -14040
rect 8626 -14100 8636 -14040
rect 8236 -14209 8636 -14100
rect 8692 -14040 9092 -14030
rect 8692 -14100 8702 -14040
rect 8762 -14100 9022 -14040
rect 9082 -14100 9092 -14040
rect 8692 -14209 9092 -14100
rect 9150 -14040 9550 -14030
rect 9150 -14100 9160 -14040
rect 9220 -14100 9480 -14040
rect 9540 -14100 9550 -14040
rect 9150 -14209 9550 -14100
rect 9606 -14040 10006 -14030
rect 9606 -14100 9616 -14040
rect 9676 -14100 9936 -14040
rect 9996 -14100 10006 -14040
rect 9606 -14209 10006 -14100
rect 10062 -14040 10462 -14030
rect 10062 -14100 10072 -14040
rect 10132 -14100 10392 -14040
rect 10452 -14100 10462 -14040
rect 10062 -14209 10462 -14100
rect 10520 -14040 10920 -14030
rect 10520 -14100 10530 -14040
rect 10590 -14100 10850 -14040
rect 10910 -14100 10920 -14040
rect 10520 -14209 10920 -14100
rect 7306 -14279 9093 -14209
rect 9150 -14279 10920 -14209
rect 7306 -14390 7706 -14279
rect 7306 -14450 7316 -14390
rect 7376 -14450 7636 -14390
rect 7696 -14450 7706 -14390
rect 7306 -14460 7706 -14450
rect 7762 -14390 8162 -14279
rect 7762 -14450 7772 -14390
rect 7832 -14450 8092 -14390
rect 8152 -14450 8162 -14390
rect 7762 -14460 8162 -14450
rect 8236 -14390 8636 -14279
rect 8236 -14450 8246 -14390
rect 8306 -14450 8566 -14390
rect 8626 -14450 8636 -14390
rect 8236 -14460 8636 -14450
rect 8692 -14390 9092 -14279
rect 8692 -14450 8702 -14390
rect 8762 -14450 9022 -14390
rect 9082 -14450 9092 -14390
rect 8692 -14460 9092 -14450
rect 9150 -14390 9550 -14279
rect 9150 -14450 9160 -14390
rect 9220 -14450 9480 -14390
rect 9540 -14450 9550 -14390
rect 9150 -14460 9550 -14450
rect 9606 -14390 10006 -14279
rect 9606 -14450 9616 -14390
rect 9676 -14450 9936 -14390
rect 9996 -14450 10006 -14390
rect 9606 -14460 10006 -14450
rect 10062 -14390 10462 -14279
rect 10062 -14450 10072 -14390
rect 10132 -14450 10392 -14390
rect 10452 -14450 10462 -14390
rect 10062 -14460 10462 -14450
rect 10520 -14390 10920 -14279
rect 10520 -14450 10530 -14390
rect 10590 -14450 10850 -14390
rect 10910 -14450 10920 -14390
rect 10520 -14460 10920 -14450
rect 10976 -14040 11376 -14030
rect 10976 -14100 10986 -14040
rect 11046 -14100 11306 -14040
rect 11366 -14100 11376 -14040
rect 10976 -14209 11376 -14100
rect 11432 -14040 11832 -14030
rect 11432 -14100 11442 -14040
rect 11502 -14100 11762 -14040
rect 11822 -14100 11832 -14040
rect 11432 -14209 11832 -14100
rect 11890 -14040 12290 -14030
rect 11890 -14100 11900 -14040
rect 11960 -14100 12220 -14040
rect 12280 -14100 12290 -14040
rect 11890 -14209 12290 -14100
rect 10976 -14279 12290 -14209
rect 10976 -14390 11376 -14279
rect 10976 -14450 10986 -14390
rect 11046 -14450 11306 -14390
rect 11366 -14450 11376 -14390
rect 10976 -14460 11376 -14450
rect 11432 -14390 11832 -14279
rect 11432 -14450 11442 -14390
rect 11502 -14450 11762 -14390
rect 11822 -14450 11832 -14390
rect 11432 -14460 11832 -14450
rect 11890 -14390 12290 -14279
rect 11890 -14450 11900 -14390
rect 11960 -14450 12220 -14390
rect 12280 -14450 12290 -14390
rect 11890 -14460 12290 -14450
rect 12346 -14040 12746 -14030
rect 12346 -14100 12356 -14040
rect 12416 -14100 12676 -14040
rect 12736 -14100 12746 -14040
rect 12346 -14209 12746 -14100
rect 12802 -14040 13202 -14030
rect 12802 -14100 12812 -14040
rect 12872 -14100 13132 -14040
rect 13192 -14100 13202 -14040
rect 12802 -14209 13202 -14100
rect 12346 -14279 13202 -14209
rect 12346 -14390 12746 -14279
rect 12346 -14450 12356 -14390
rect 12416 -14450 12676 -14390
rect 12736 -14450 12746 -14390
rect 12346 -14460 12746 -14450
rect 12802 -14390 13202 -14279
rect 12802 -14450 12812 -14390
rect 12872 -14450 13132 -14390
rect 13192 -14450 13202 -14390
rect 12802 -14460 13202 -14450
rect 13260 -14040 13660 -14030
rect 13260 -14100 13270 -14040
rect 13330 -14100 13590 -14040
rect 13650 -14100 13660 -14040
rect 13260 -14209 13660 -14100
rect 13716 -14040 14116 -14030
rect 13716 -14100 13726 -14040
rect 13786 -14100 14046 -14040
rect 14106 -14100 14116 -14040
rect 13716 -14209 14116 -14100
rect 14172 -14040 14572 -14030
rect 14172 -14100 14182 -14040
rect 14242 -14100 14502 -14040
rect 14562 -14100 14572 -14040
rect 14172 -14209 14572 -14100
rect 14630 -14040 15030 -14030
rect 14630 -14100 14640 -14040
rect 14700 -14100 14960 -14040
rect 15020 -14100 15030 -14040
rect 14630 -14209 15030 -14100
rect 15086 -14040 15486 -14030
rect 15086 -14100 15096 -14040
rect 15156 -14100 15416 -14040
rect 15476 -14100 15486 -14040
rect 15086 -14209 15486 -14100
rect 13260 -14279 15486 -14209
rect 13260 -14390 13660 -14279
rect 13260 -14450 13270 -14390
rect 13330 -14450 13590 -14390
rect 13650 -14450 13660 -14390
rect 13260 -14460 13660 -14450
rect 13716 -14390 14116 -14279
rect 13716 -14450 13726 -14390
rect 13786 -14450 14046 -14390
rect 14106 -14450 14116 -14390
rect 13716 -14460 14116 -14450
rect 14172 -14390 14572 -14279
rect 14172 -14450 14182 -14390
rect 14242 -14450 14502 -14390
rect 14562 -14450 14572 -14390
rect 14172 -14460 14572 -14450
rect 14630 -14390 15030 -14279
rect 14630 -14450 14640 -14390
rect 14700 -14450 14960 -14390
rect 15020 -14450 15030 -14390
rect 14630 -14460 15030 -14450
rect 15086 -14390 15486 -14279
rect 15086 -14450 15096 -14390
rect 15156 -14450 15416 -14390
rect 15476 -14450 15486 -14390
rect 15086 -14460 15486 -14450
rect 66 -14532 80 -14460
rect 456 -14532 526 -14460
rect 912 -14532 983 -14460
rect 1370 -14532 1441 -14460
rect 1826 -14532 1897 -14460
rect 2282 -14532 2353 -14460
rect 2740 -14532 2811 -14460
rect 3196 -14532 3267 -14460
rect 3652 -14532 3723 -14460
rect 4110 -14532 4181 -14460
rect 4566 -14532 4637 -14460
rect 5022 -14532 5093 -14460
rect 5480 -14532 5551 -14460
rect 5936 -14532 6007 -14460
rect 6392 -14532 6463 -14460
rect 6850 -14532 6921 -14460
rect 7306 -14532 7377 -14460
rect 7762 -14532 7833 -14460
rect 8236 -14532 8307 -14460
rect 8692 -14532 8763 -14460
rect 9150 -14532 9221 -14460
rect 9606 -14532 9677 -14460
rect 10062 -14532 10133 -14460
rect 10520 -14532 10591 -14460
rect 10976 -14532 11047 -14460
rect 11432 -14532 11503 -14460
rect 11890 -14532 11961 -14460
rect 12346 -14532 12417 -14460
rect 12802 -14532 12873 -14460
rect 13260 -14532 13331 -14460
rect 66 -14542 400 -14532
rect 0 -14602 10 -14542
rect 70 -14602 330 -14542
rect 390 -14602 400 -14542
rect 0 -14892 14 -14602
rect 66 -14892 400 -14602
rect 0 -14952 10 -14892
rect 70 -14952 330 -14892
rect 390 -14952 400 -14892
rect 0 -15034 14 -14952
rect 66 -14962 400 -14952
rect 456 -14542 856 -14532
rect 456 -14602 466 -14542
rect 526 -14602 786 -14542
rect 846 -14602 856 -14542
rect 456 -14711 856 -14602
rect 912 -14542 1312 -14532
rect 912 -14602 922 -14542
rect 982 -14602 1242 -14542
rect 1302 -14602 1312 -14542
rect 912 -14711 1312 -14602
rect 1370 -14542 1770 -14532
rect 1370 -14602 1380 -14542
rect 1440 -14602 1700 -14542
rect 1760 -14602 1770 -14542
rect 1370 -14711 1770 -14602
rect 1826 -14542 2226 -14532
rect 1826 -14602 1836 -14542
rect 1896 -14602 2156 -14542
rect 2216 -14602 2226 -14542
rect 1826 -14711 2226 -14602
rect 2282 -14542 2682 -14532
rect 2282 -14602 2292 -14542
rect 2352 -14602 2612 -14542
rect 2672 -14602 2682 -14542
rect 2282 -14711 2682 -14602
rect 2740 -14542 3140 -14532
rect 2740 -14602 2750 -14542
rect 2810 -14602 3070 -14542
rect 3130 -14602 3140 -14542
rect 2740 -14711 3140 -14602
rect 3196 -14542 3596 -14532
rect 3196 -14602 3206 -14542
rect 3266 -14602 3526 -14542
rect 3586 -14602 3596 -14542
rect 3196 -14711 3596 -14602
rect 456 -14781 3596 -14711
rect 456 -14782 2682 -14781
rect 456 -14892 856 -14782
rect 456 -14952 466 -14892
rect 526 -14952 786 -14892
rect 846 -14952 856 -14892
rect 456 -14962 856 -14952
rect 912 -14892 1312 -14782
rect 912 -14952 922 -14892
rect 982 -14952 1242 -14892
rect 1302 -14952 1312 -14892
rect 912 -14962 1312 -14952
rect 1370 -14892 1770 -14782
rect 1370 -14952 1380 -14892
rect 1440 -14952 1700 -14892
rect 1760 -14952 1770 -14892
rect 1370 -14962 1770 -14952
rect 1826 -14892 2226 -14782
rect 1826 -14952 1836 -14892
rect 1896 -14952 2156 -14892
rect 2216 -14952 2226 -14892
rect 1826 -14962 2226 -14952
rect 2282 -14892 2682 -14782
rect 2282 -14952 2292 -14892
rect 2352 -14952 2612 -14892
rect 2672 -14952 2682 -14892
rect 2282 -14962 2682 -14952
rect 2740 -14782 3596 -14781
rect 2740 -14892 3140 -14782
rect 2740 -14952 2750 -14892
rect 2810 -14952 3070 -14892
rect 3130 -14952 3140 -14892
rect 2740 -14962 3140 -14952
rect 3196 -14892 3596 -14782
rect 3196 -14952 3206 -14892
rect 3266 -14952 3526 -14892
rect 3586 -14952 3596 -14892
rect 3196 -14962 3596 -14952
rect 3652 -14542 4052 -14532
rect 3652 -14602 3662 -14542
rect 3722 -14602 3982 -14542
rect 4042 -14602 4052 -14542
rect 3652 -14711 4052 -14602
rect 4110 -14542 4510 -14532
rect 4110 -14602 4120 -14542
rect 4180 -14602 4440 -14542
rect 4500 -14602 4510 -14542
rect 4110 -14711 4510 -14602
rect 4566 -14542 4966 -14532
rect 4566 -14602 4576 -14542
rect 4636 -14602 4896 -14542
rect 4956 -14602 4966 -14542
rect 4566 -14711 4966 -14602
rect 5022 -14542 5422 -14532
rect 5022 -14602 5032 -14542
rect 5092 -14602 5352 -14542
rect 5412 -14602 5422 -14542
rect 5022 -14711 5422 -14602
rect 5480 -14542 5880 -14532
rect 5480 -14602 5490 -14542
rect 5550 -14602 5810 -14542
rect 5870 -14602 5880 -14542
rect 5480 -14711 5880 -14602
rect 5936 -14542 6336 -14532
rect 5936 -14602 5946 -14542
rect 6006 -14602 6266 -14542
rect 6326 -14602 6336 -14542
rect 5936 -14711 6336 -14602
rect 6392 -14542 6792 -14532
rect 6392 -14602 6402 -14542
rect 6462 -14602 6722 -14542
rect 6782 -14602 6792 -14542
rect 6392 -14711 6792 -14602
rect 6850 -14542 7250 -14532
rect 6850 -14602 6860 -14542
rect 6920 -14602 7180 -14542
rect 7240 -14602 7250 -14542
rect 6850 -14711 7250 -14602
rect 3652 -14782 7250 -14711
rect 3652 -14892 4052 -14782
rect 3652 -14952 3662 -14892
rect 3722 -14952 3982 -14892
rect 4042 -14952 4052 -14892
rect 3652 -14962 4052 -14952
rect 4110 -14892 4510 -14782
rect 4110 -14952 4120 -14892
rect 4180 -14952 4440 -14892
rect 4500 -14952 4510 -14892
rect 4110 -14962 4510 -14952
rect 4566 -14892 4966 -14782
rect 4566 -14952 4576 -14892
rect 4636 -14952 4896 -14892
rect 4956 -14952 4966 -14892
rect 4566 -14962 4966 -14952
rect 5022 -14892 5422 -14782
rect 5022 -14952 5032 -14892
rect 5092 -14952 5352 -14892
rect 5412 -14952 5422 -14892
rect 5022 -14962 5422 -14952
rect 5480 -14892 5880 -14782
rect 5480 -14952 5490 -14892
rect 5550 -14952 5810 -14892
rect 5870 -14952 5880 -14892
rect 5480 -14962 5880 -14952
rect 5936 -14892 6336 -14782
rect 5936 -14952 5946 -14892
rect 6006 -14952 6266 -14892
rect 6326 -14952 6336 -14892
rect 5936 -14962 6336 -14952
rect 6392 -14892 6792 -14782
rect 6392 -14952 6402 -14892
rect 6462 -14952 6722 -14892
rect 6782 -14952 6792 -14892
rect 6392 -14962 6792 -14952
rect 6850 -14892 7250 -14782
rect 6850 -14952 6860 -14892
rect 6920 -14952 7180 -14892
rect 7240 -14952 7250 -14892
rect 6850 -14962 7250 -14952
rect 7306 -14542 7706 -14532
rect 7306 -14602 7316 -14542
rect 7376 -14602 7636 -14542
rect 7696 -14602 7706 -14542
rect 7306 -14711 7706 -14602
rect 7762 -14542 8162 -14532
rect 7762 -14602 7772 -14542
rect 7832 -14602 8092 -14542
rect 8152 -14602 8162 -14542
rect 7762 -14711 8162 -14602
rect 8236 -14542 8636 -14532
rect 8236 -14602 8246 -14542
rect 8306 -14602 8566 -14542
rect 8626 -14602 8636 -14542
rect 8236 -14711 8636 -14602
rect 8692 -14542 9092 -14532
rect 8692 -14602 8702 -14542
rect 8762 -14602 9022 -14542
rect 9082 -14602 9092 -14542
rect 8692 -14711 9092 -14602
rect 9150 -14542 9550 -14532
rect 9150 -14602 9160 -14542
rect 9220 -14602 9480 -14542
rect 9540 -14602 9550 -14542
rect 9150 -14711 9550 -14602
rect 9606 -14542 10006 -14532
rect 9606 -14602 9616 -14542
rect 9676 -14602 9936 -14542
rect 9996 -14602 10006 -14542
rect 9606 -14711 10006 -14602
rect 10062 -14542 10462 -14532
rect 10062 -14602 10072 -14542
rect 10132 -14602 10392 -14542
rect 10452 -14602 10462 -14542
rect 10062 -14711 10462 -14602
rect 10520 -14542 10920 -14532
rect 10520 -14602 10530 -14542
rect 10590 -14602 10850 -14542
rect 10910 -14602 10920 -14542
rect 10520 -14711 10920 -14602
rect 7306 -14782 9093 -14711
rect 9150 -14781 10920 -14711
rect 9150 -14782 10462 -14781
rect 7306 -14892 7706 -14782
rect 7306 -14952 7316 -14892
rect 7376 -14952 7636 -14892
rect 7696 -14952 7706 -14892
rect 7306 -14962 7706 -14952
rect 7762 -14892 8162 -14782
rect 7762 -14952 7772 -14892
rect 7832 -14952 8092 -14892
rect 8152 -14952 8162 -14892
rect 7762 -14962 8162 -14952
rect 8236 -14892 8636 -14782
rect 8236 -14952 8246 -14892
rect 8306 -14952 8566 -14892
rect 8626 -14952 8636 -14892
rect 8236 -14962 8636 -14952
rect 8692 -14892 9092 -14782
rect 8692 -14952 8702 -14892
rect 8762 -14952 9022 -14892
rect 9082 -14952 9092 -14892
rect 8692 -14962 9092 -14952
rect 9150 -14892 9550 -14782
rect 9150 -14952 9160 -14892
rect 9220 -14952 9480 -14892
rect 9540 -14952 9550 -14892
rect 9150 -14962 9550 -14952
rect 9606 -14892 10006 -14782
rect 9606 -14952 9616 -14892
rect 9676 -14952 9936 -14892
rect 9996 -14952 10006 -14892
rect 9606 -14962 10006 -14952
rect 10062 -14892 10462 -14782
rect 10062 -14952 10072 -14892
rect 10132 -14952 10392 -14892
rect 10452 -14952 10462 -14892
rect 10062 -14962 10462 -14952
rect 10520 -14892 10920 -14781
rect 10520 -14952 10530 -14892
rect 10590 -14952 10850 -14892
rect 10910 -14952 10920 -14892
rect 10520 -14962 10920 -14952
rect 10976 -14542 11376 -14532
rect 10976 -14602 10986 -14542
rect 11046 -14602 11306 -14542
rect 11366 -14602 11376 -14542
rect 10976 -14711 11376 -14602
rect 11432 -14542 11832 -14532
rect 11432 -14602 11442 -14542
rect 11502 -14602 11762 -14542
rect 11822 -14602 11832 -14542
rect 11432 -14711 11832 -14602
rect 11890 -14542 12290 -14532
rect 11890 -14602 11900 -14542
rect 11960 -14602 12220 -14542
rect 12280 -14602 12290 -14542
rect 11890 -14711 12290 -14602
rect 10976 -14782 12290 -14711
rect 10976 -14892 11376 -14782
rect 10976 -14952 10986 -14892
rect 11046 -14952 11306 -14892
rect 11366 -14952 11376 -14892
rect 10976 -14962 11376 -14952
rect 11432 -14892 11832 -14782
rect 11432 -14952 11442 -14892
rect 11502 -14952 11762 -14892
rect 11822 -14952 11832 -14892
rect 11432 -14962 11832 -14952
rect 11890 -14892 12290 -14782
rect 11890 -14952 11900 -14892
rect 11960 -14952 12220 -14892
rect 12280 -14952 12290 -14892
rect 11890 -14962 12290 -14952
rect 12346 -14542 12746 -14532
rect 12346 -14602 12356 -14542
rect 12416 -14602 12676 -14542
rect 12736 -14602 12746 -14542
rect 12346 -14711 12746 -14602
rect 12802 -14542 13202 -14532
rect 12802 -14602 12812 -14542
rect 12872 -14602 13132 -14542
rect 13192 -14602 13202 -14542
rect 12802 -14711 13202 -14602
rect 12346 -14782 13202 -14711
rect 12346 -14892 12746 -14782
rect 12346 -14952 12356 -14892
rect 12416 -14952 12676 -14892
rect 12736 -14952 12746 -14892
rect 12346 -14962 12746 -14952
rect 12802 -14892 13202 -14782
rect 12802 -14952 12812 -14892
rect 12872 -14952 13132 -14892
rect 13192 -14952 13202 -14892
rect 12802 -14962 13202 -14952
rect 13260 -14542 13660 -14532
rect 13260 -14602 13270 -14542
rect 13330 -14602 13590 -14542
rect 13650 -14602 13660 -14542
rect 13260 -14892 13660 -14602
rect 13260 -14952 13270 -14892
rect 13330 -14952 13590 -14892
rect 13650 -14952 13660 -14892
rect 13260 -14962 13660 -14952
rect 13716 -14542 14116 -14532
rect 13716 -14602 13726 -14542
rect 13786 -14602 14046 -14542
rect 14106 -14602 14116 -14542
rect 13716 -14711 14116 -14602
rect 14172 -14542 14572 -14532
rect 14172 -14602 14182 -14542
rect 14242 -14602 14502 -14542
rect 14562 -14602 14572 -14542
rect 14172 -14711 14572 -14602
rect 14630 -14542 15030 -14532
rect 14630 -14602 14640 -14542
rect 14700 -14602 14960 -14542
rect 15020 -14602 15030 -14542
rect 14630 -14711 15030 -14602
rect 15086 -14542 15486 -14532
rect 15086 -14602 15096 -14542
rect 15156 -14602 15416 -14542
rect 15476 -14602 15486 -14542
rect 15086 -14710 15486 -14602
rect 15086 -14711 15721 -14710
rect 13716 -14781 15721 -14711
rect 13716 -14782 15486 -14781
rect 13716 -14892 14116 -14782
rect 13716 -14952 13726 -14892
rect 13786 -14952 14046 -14892
rect 14106 -14952 14116 -14892
rect 13716 -14962 14116 -14952
rect 14172 -14892 14572 -14782
rect 14172 -14952 14182 -14892
rect 14242 -14952 14502 -14892
rect 14562 -14952 14572 -14892
rect 14172 -14962 14572 -14952
rect 14630 -14892 15030 -14782
rect 14630 -14952 14640 -14892
rect 14700 -14952 14960 -14892
rect 15020 -14952 15030 -14892
rect 14630 -14962 15030 -14952
rect 15086 -14892 15486 -14782
rect 15086 -14952 15096 -14892
rect 15156 -14952 15416 -14892
rect 15476 -14952 15486 -14892
rect 15086 -14962 15486 -14952
rect 66 -15024 80 -14962
rect 456 -15024 527 -14962
rect 912 -15024 983 -14962
rect 1370 -15024 1441 -14962
rect 1826 -15024 1897 -14962
rect 2282 -15024 2353 -14962
rect 2740 -15024 2810 -14962
rect 3196 -15024 3266 -14962
rect 3652 -15024 3722 -14962
rect 4110 -15024 4180 -14962
rect 4566 -15024 4636 -14962
rect 5022 -15024 5092 -14962
rect 5480 -15024 5550 -14962
rect 5936 -15024 6006 -14962
rect 6392 -15024 6462 -14962
rect 6850 -15024 6920 -14962
rect 7306 -15024 7376 -14962
rect 7762 -15024 7832 -14962
rect 8236 -15024 8306 -14962
rect 8692 -15024 8762 -14962
rect 9150 -15024 9220 -14962
rect 9606 -15024 9676 -14962
rect 10062 -15024 10132 -14962
rect 10520 -15024 10590 -14962
rect 10976 -15024 11046 -14962
rect 11432 -15024 11502 -14962
rect 12346 -15024 12416 -14962
rect 12802 -15024 12872 -14962
rect 13260 -15024 13330 -14962
rect 13716 -15024 13786 -14962
rect 66 -15034 400 -15024
rect 0 -15094 10 -15034
rect 70 -15094 330 -15034
rect 390 -15094 400 -15034
rect 0 -15384 14 -15094
rect 66 -15384 400 -15094
rect 0 -15444 10 -15384
rect 70 -15444 330 -15384
rect 390 -15444 400 -15384
rect 0 -15550 14 -15444
rect 66 -15454 400 -15444
rect 456 -15034 856 -15024
rect 456 -15094 466 -15034
rect 526 -15094 786 -15034
rect 846 -15094 856 -15034
rect 456 -15204 856 -15094
rect 912 -15034 1312 -15024
rect 912 -15094 922 -15034
rect 982 -15094 1242 -15034
rect 1302 -15094 1312 -15034
rect 912 -15204 1312 -15094
rect 1370 -15034 1770 -15024
rect 1370 -15094 1380 -15034
rect 1440 -15094 1700 -15034
rect 1760 -15094 1770 -15034
rect 1370 -15204 1770 -15094
rect 1826 -15034 2226 -15024
rect 1826 -15094 1836 -15034
rect 1896 -15094 2156 -15034
rect 2216 -15094 2226 -15034
rect 1826 -15204 2226 -15094
rect 2282 -15034 2682 -15024
rect 2282 -15094 2292 -15034
rect 2352 -15094 2612 -15034
rect 2672 -15094 2682 -15034
rect 2282 -15204 2682 -15094
rect 2740 -15034 3140 -15024
rect 2740 -15094 2750 -15034
rect 2810 -15094 3070 -15034
rect 3130 -15094 3140 -15034
rect 2740 -15204 3140 -15094
rect 3196 -15034 3596 -15024
rect 3196 -15094 3206 -15034
rect 3266 -15094 3526 -15034
rect 3586 -15094 3596 -15034
rect 3196 -15204 3596 -15094
rect 456 -15274 3596 -15204
rect 456 -15384 856 -15274
rect 456 -15444 466 -15384
rect 526 -15444 786 -15384
rect 846 -15444 856 -15384
rect 456 -15454 856 -15444
rect 912 -15384 1312 -15274
rect 912 -15444 922 -15384
rect 982 -15444 1242 -15384
rect 1302 -15444 1312 -15384
rect 912 -15454 1312 -15444
rect 1370 -15384 1770 -15274
rect 1370 -15444 1380 -15384
rect 1440 -15444 1700 -15384
rect 1760 -15444 1770 -15384
rect 1370 -15454 1770 -15444
rect 1826 -15384 2226 -15274
rect 1826 -15444 1836 -15384
rect 1896 -15444 2156 -15384
rect 2216 -15444 2226 -15384
rect 1826 -15454 2226 -15444
rect 2282 -15384 2682 -15274
rect 2282 -15444 2292 -15384
rect 2352 -15444 2612 -15384
rect 2672 -15444 2682 -15384
rect 2282 -15454 2682 -15444
rect 2740 -15384 3140 -15274
rect 2740 -15444 2750 -15384
rect 2810 -15444 3070 -15384
rect 3130 -15444 3140 -15384
rect 2740 -15454 3140 -15444
rect 3196 -15384 3596 -15274
rect 3196 -15444 3206 -15384
rect 3266 -15444 3526 -15384
rect 3586 -15444 3596 -15384
rect 3196 -15454 3596 -15444
rect 3652 -15034 4052 -15024
rect 3652 -15094 3662 -15034
rect 3722 -15094 3982 -15034
rect 4042 -15094 4052 -15034
rect 3652 -15204 4052 -15094
rect 4110 -15034 4510 -15024
rect 4110 -15094 4120 -15034
rect 4180 -15094 4440 -15034
rect 4500 -15094 4510 -15034
rect 4110 -15204 4510 -15094
rect 4566 -15034 4966 -15024
rect 4566 -15094 4576 -15034
rect 4636 -15094 4896 -15034
rect 4956 -15094 4966 -15034
rect 4566 -15204 4966 -15094
rect 5022 -15034 5422 -15024
rect 5022 -15094 5032 -15034
rect 5092 -15094 5352 -15034
rect 5412 -15094 5422 -15034
rect 5022 -15204 5422 -15094
rect 5480 -15034 5880 -15024
rect 5480 -15094 5490 -15034
rect 5550 -15094 5810 -15034
rect 5870 -15094 5880 -15034
rect 5480 -15204 5880 -15094
rect 5936 -15034 6336 -15024
rect 5936 -15094 5946 -15034
rect 6006 -15094 6266 -15034
rect 6326 -15094 6336 -15034
rect 5936 -15204 6336 -15094
rect 6392 -15034 6792 -15024
rect 6392 -15094 6402 -15034
rect 6462 -15094 6722 -15034
rect 6782 -15094 6792 -15034
rect 6392 -15204 6792 -15094
rect 6850 -15034 7250 -15024
rect 6850 -15094 6860 -15034
rect 6920 -15094 7180 -15034
rect 7240 -15094 7250 -15034
rect 6850 -15204 7250 -15094
rect 3652 -15274 7250 -15204
rect 3652 -15384 4052 -15274
rect 3652 -15444 3662 -15384
rect 3722 -15444 3982 -15384
rect 4042 -15444 4052 -15384
rect 3652 -15454 4052 -15444
rect 4110 -15384 4510 -15274
rect 4110 -15444 4120 -15384
rect 4180 -15444 4440 -15384
rect 4500 -15444 4510 -15384
rect 4110 -15454 4510 -15444
rect 4566 -15384 4966 -15274
rect 4566 -15444 4576 -15384
rect 4636 -15444 4896 -15384
rect 4956 -15444 4966 -15384
rect 4566 -15454 4966 -15444
rect 5022 -15384 5422 -15274
rect 5022 -15444 5032 -15384
rect 5092 -15444 5352 -15384
rect 5412 -15444 5422 -15384
rect 5022 -15454 5422 -15444
rect 5480 -15384 5880 -15274
rect 5480 -15444 5490 -15384
rect 5550 -15444 5810 -15384
rect 5870 -15444 5880 -15384
rect 5480 -15454 5880 -15444
rect 5936 -15384 6336 -15274
rect 5936 -15444 5946 -15384
rect 6006 -15444 6266 -15384
rect 6326 -15444 6336 -15384
rect 5936 -15454 6336 -15444
rect 6392 -15384 6792 -15274
rect 6392 -15444 6402 -15384
rect 6462 -15444 6722 -15384
rect 6782 -15444 6792 -15384
rect 6392 -15454 6792 -15444
rect 6850 -15384 7250 -15274
rect 6850 -15444 6860 -15384
rect 6920 -15444 7180 -15384
rect 7240 -15444 7250 -15384
rect 6850 -15454 7250 -15444
rect 7306 -15034 7706 -15024
rect 7306 -15094 7316 -15034
rect 7376 -15094 7636 -15034
rect 7696 -15094 7706 -15034
rect 7306 -15204 7706 -15094
rect 7762 -15034 8162 -15024
rect 7762 -15094 7772 -15034
rect 7832 -15094 8092 -15034
rect 8152 -15094 8162 -15034
rect 7762 -15204 8162 -15094
rect 8236 -15034 8636 -15024
rect 8236 -15094 8246 -15034
rect 8306 -15094 8566 -15034
rect 8626 -15094 8636 -15034
rect 8236 -15204 8636 -15094
rect 8692 -15034 9092 -15024
rect 8692 -15094 8702 -15034
rect 8762 -15094 9022 -15034
rect 9082 -15094 9092 -15034
rect 8692 -15204 9092 -15094
rect 9150 -15034 9550 -15024
rect 9150 -15094 9160 -15034
rect 9220 -15094 9480 -15034
rect 9540 -15094 9550 -15034
rect 9150 -15204 9550 -15094
rect 9606 -15034 10006 -15024
rect 9606 -15094 9616 -15034
rect 9676 -15094 9936 -15034
rect 9996 -15094 10006 -15034
rect 9606 -15204 10006 -15094
rect 10062 -15034 10462 -15024
rect 10062 -15094 10072 -15034
rect 10132 -15094 10392 -15034
rect 10452 -15094 10462 -15034
rect 10062 -15204 10462 -15094
rect 10520 -15034 10920 -15024
rect 10520 -15094 10530 -15034
rect 10590 -15094 10850 -15034
rect 10910 -15094 10920 -15034
rect 10520 -15204 10920 -15094
rect 7306 -15274 9093 -15204
rect 9150 -15274 10920 -15204
rect 7306 -15384 7706 -15274
rect 7306 -15444 7316 -15384
rect 7376 -15444 7636 -15384
rect 7696 -15444 7706 -15384
rect 7306 -15454 7706 -15444
rect 7762 -15384 8162 -15274
rect 7762 -15444 7772 -15384
rect 7832 -15444 8092 -15384
rect 8152 -15444 8162 -15384
rect 7762 -15454 8162 -15444
rect 8236 -15384 8636 -15274
rect 8236 -15444 8246 -15384
rect 8306 -15444 8566 -15384
rect 8626 -15444 8636 -15384
rect 8236 -15454 8636 -15444
rect 8692 -15384 9092 -15274
rect 8692 -15444 8702 -15384
rect 8762 -15444 9022 -15384
rect 9082 -15444 9092 -15384
rect 8692 -15454 9092 -15444
rect 9150 -15384 9550 -15274
rect 9150 -15444 9160 -15384
rect 9220 -15444 9480 -15384
rect 9540 -15444 9550 -15384
rect 9150 -15454 9550 -15444
rect 9606 -15384 10006 -15274
rect 9606 -15444 9616 -15384
rect 9676 -15444 9936 -15384
rect 9996 -15444 10006 -15384
rect 9606 -15454 10006 -15444
rect 10062 -15384 10462 -15274
rect 10062 -15444 10072 -15384
rect 10132 -15444 10392 -15384
rect 10452 -15444 10462 -15384
rect 10062 -15454 10462 -15444
rect 10520 -15384 10920 -15274
rect 10520 -15444 10530 -15384
rect 10590 -15444 10850 -15384
rect 10910 -15444 10920 -15384
rect 10520 -15454 10920 -15444
rect 10976 -15034 11376 -15024
rect 10976 -15094 10986 -15034
rect 11046 -15094 11306 -15034
rect 11366 -15094 11376 -15034
rect 10976 -15204 11376 -15094
rect 11432 -15034 11832 -15024
rect 11432 -15094 11442 -15034
rect 11502 -15094 11762 -15034
rect 11822 -15094 11832 -15034
rect 11432 -15204 11832 -15094
rect 10976 -15274 11832 -15204
rect 10976 -15384 11376 -15274
rect 10976 -15444 10986 -15384
rect 11046 -15444 11306 -15384
rect 11366 -15444 11376 -15384
rect 10976 -15454 11376 -15444
rect 11432 -15384 11832 -15274
rect 11432 -15444 11442 -15384
rect 11502 -15444 11762 -15384
rect 11822 -15444 11832 -15384
rect 11432 -15454 11832 -15444
rect 11890 -15034 12290 -15024
rect 11890 -15094 11900 -15034
rect 11960 -15094 12220 -15034
rect 12280 -15094 12290 -15034
rect 11890 -15204 12290 -15094
rect 12346 -15034 12746 -15024
rect 12346 -15094 12356 -15034
rect 12416 -15094 12676 -15034
rect 12736 -15094 12746 -15034
rect 12346 -15204 12746 -15094
rect 12802 -15034 13202 -15024
rect 12802 -15094 12812 -15034
rect 12872 -15094 13132 -15034
rect 13192 -15094 13202 -15034
rect 12802 -15204 13202 -15094
rect 11890 -15274 13202 -15204
rect 11890 -15384 12290 -15274
rect 11890 -15444 11900 -15384
rect 11960 -15444 12220 -15384
rect 12280 -15444 12290 -15384
rect 11890 -15454 12290 -15444
rect 12346 -15384 12746 -15274
rect 12346 -15444 12356 -15384
rect 12416 -15444 12676 -15384
rect 12736 -15444 12746 -15384
rect 12346 -15454 12746 -15444
rect 12802 -15384 13202 -15274
rect 12802 -15444 12812 -15384
rect 12872 -15444 13132 -15384
rect 13192 -15444 13202 -15384
rect 12802 -15454 13202 -15444
rect 13260 -15034 13660 -15024
rect 13260 -15094 13270 -15034
rect 13330 -15094 13590 -15034
rect 13650 -15094 13660 -15034
rect 13260 -15384 13660 -15094
rect 13260 -15444 13270 -15384
rect 13330 -15444 13590 -15384
rect 13650 -15444 13660 -15384
rect 13260 -15454 13660 -15444
rect 13716 -15034 14116 -15024
rect 13716 -15094 13726 -15034
rect 13786 -15094 14046 -15034
rect 14106 -15094 14116 -15034
rect 13716 -15384 14116 -15094
rect 13716 -15444 13726 -15384
rect 13786 -15444 14046 -15384
rect 14106 -15444 14116 -15384
rect 13716 -15454 14116 -15444
rect 14172 -15034 14572 -15024
rect 14172 -15094 14182 -15034
rect 14242 -15094 14502 -15034
rect 14562 -15094 14572 -15034
rect 14172 -15200 14572 -15094
rect 14630 -15034 15030 -15024
rect 14630 -15094 14640 -15034
rect 14700 -15094 14960 -15034
rect 15020 -15094 15030 -15034
rect 14630 -15200 15030 -15094
rect 14172 -15204 15030 -15200
rect 15086 -15034 15486 -15024
rect 15086 -15094 15096 -15034
rect 15156 -15094 15416 -15034
rect 15476 -15094 15486 -15034
rect 15086 -15204 15486 -15094
rect 14172 -15205 15486 -15204
rect 14172 -15270 15720 -15205
rect 14172 -15275 14571 -15270
rect 14630 -15274 15720 -15270
rect 14172 -15384 14572 -15275
rect 14172 -15444 14182 -15384
rect 14242 -15444 14502 -15384
rect 14562 -15444 14572 -15384
rect 14172 -15454 14572 -15444
rect 14630 -15384 15030 -15274
rect 14630 -15444 14640 -15384
rect 14700 -15444 14960 -15384
rect 15020 -15444 15030 -15384
rect 14630 -15454 15030 -15444
rect 15086 -15276 15720 -15274
rect 15086 -15384 15486 -15276
rect 15086 -15444 15096 -15384
rect 15156 -15444 15416 -15384
rect 15476 -15444 15486 -15384
rect 15086 -15454 15486 -15444
rect 66 -15540 80 -15454
rect 456 -15540 526 -15454
rect 912 -15540 982 -15454
rect 1370 -15540 1440 -15454
rect 1826 -15540 1896 -15454
rect 2282 -15540 2352 -15454
rect 2740 -15540 2810 -15454
rect 3196 -15540 3266 -15454
rect 3652 -15540 3722 -15454
rect 4110 -15540 4180 -15454
rect 4566 -15540 4636 -15454
rect 5022 -15540 5092 -15454
rect 5480 -15540 5550 -15454
rect 5936 -15540 6006 -15454
rect 6392 -15540 6462 -15454
rect 7306 -15540 7376 -15454
rect 7762 -15540 7832 -15454
rect 8236 -15540 8306 -15454
rect 8692 -15540 8762 -15454
rect 9150 -15540 9220 -15454
rect 9606 -15540 9676 -15454
rect 10062 -15540 10132 -15454
rect 10976 -15540 11046 -15454
rect 11432 -15540 11502 -15454
rect 11890 -15540 11960 -15454
rect 12346 -15540 12416 -15454
rect 12802 -15540 12872 -15454
rect 13260 -15540 13330 -15454
rect 13716 -15540 13786 -15454
rect 66 -15550 400 -15540
rect 0 -15610 10 -15550
rect 70 -15610 330 -15550
rect 390 -15610 400 -15550
rect 0 -15900 14 -15610
rect 66 -15900 400 -15610
rect 0 -15960 10 -15900
rect 70 -15960 330 -15900
rect 390 -15960 400 -15900
rect 0 -16052 14 -15960
rect 66 -15970 400 -15960
rect 456 -15550 856 -15540
rect 456 -15610 466 -15550
rect 526 -15610 786 -15550
rect 846 -15610 856 -15550
rect 456 -15720 856 -15610
rect 912 -15550 1312 -15540
rect 912 -15610 922 -15550
rect 982 -15610 1242 -15550
rect 1302 -15610 1312 -15550
rect 912 -15720 1312 -15610
rect 1370 -15550 1770 -15540
rect 1370 -15610 1380 -15550
rect 1440 -15610 1700 -15550
rect 1760 -15610 1770 -15550
rect 1370 -15720 1770 -15610
rect 1826 -15550 2226 -15540
rect 1826 -15610 1836 -15550
rect 1896 -15610 2156 -15550
rect 2216 -15610 2226 -15550
rect 1826 -15720 2226 -15610
rect 2282 -15550 2682 -15540
rect 2282 -15610 2292 -15550
rect 2352 -15610 2612 -15550
rect 2672 -15610 2682 -15550
rect 2282 -15720 2682 -15610
rect 456 -15721 2682 -15720
rect 2740 -15550 3140 -15540
rect 2740 -15610 2750 -15550
rect 2810 -15610 3070 -15550
rect 3130 -15610 3140 -15550
rect 2740 -15720 3140 -15610
rect 3196 -15550 3596 -15540
rect 3196 -15610 3206 -15550
rect 3266 -15610 3526 -15550
rect 3586 -15610 3596 -15550
rect 3196 -15720 3596 -15610
rect 2740 -15721 3596 -15720
rect 456 -15791 3596 -15721
rect 456 -15900 856 -15791
rect 456 -15960 466 -15900
rect 526 -15960 786 -15900
rect 846 -15960 856 -15900
rect 456 -15970 856 -15960
rect 912 -15900 1312 -15791
rect 912 -15960 922 -15900
rect 982 -15960 1242 -15900
rect 1302 -15960 1312 -15900
rect 912 -15970 1312 -15960
rect 1370 -15900 1770 -15791
rect 1370 -15960 1380 -15900
rect 1440 -15960 1700 -15900
rect 1760 -15960 1770 -15900
rect 1370 -15970 1770 -15960
rect 1826 -15900 2226 -15791
rect 1826 -15960 1836 -15900
rect 1896 -15960 2156 -15900
rect 2216 -15960 2226 -15900
rect 1826 -15970 2226 -15960
rect 2282 -15900 2682 -15791
rect 2282 -15960 2292 -15900
rect 2352 -15960 2612 -15900
rect 2672 -15960 2682 -15900
rect 2282 -15970 2682 -15960
rect 2740 -15900 3140 -15791
rect 2740 -15960 2750 -15900
rect 2810 -15960 3070 -15900
rect 3130 -15960 3140 -15900
rect 2740 -15970 3140 -15960
rect 3196 -15900 3596 -15791
rect 3196 -15960 3206 -15900
rect 3266 -15960 3526 -15900
rect 3586 -15960 3596 -15900
rect 3196 -15970 3596 -15960
rect 3652 -15550 4052 -15540
rect 3652 -15610 3662 -15550
rect 3722 -15610 3982 -15550
rect 4042 -15610 4052 -15550
rect 3652 -15720 4052 -15610
rect 4110 -15550 4510 -15540
rect 4110 -15610 4120 -15550
rect 4180 -15610 4440 -15550
rect 4500 -15610 4510 -15550
rect 4110 -15720 4510 -15610
rect 4566 -15550 4966 -15540
rect 4566 -15610 4576 -15550
rect 4636 -15610 4896 -15550
rect 4956 -15610 4966 -15550
rect 4566 -15720 4966 -15610
rect 5022 -15550 5422 -15540
rect 5022 -15610 5032 -15550
rect 5092 -15610 5352 -15550
rect 5412 -15610 5422 -15550
rect 5022 -15720 5422 -15610
rect 5480 -15550 5880 -15540
rect 5480 -15610 5490 -15550
rect 5550 -15610 5810 -15550
rect 5870 -15610 5880 -15550
rect 5480 -15720 5880 -15610
rect 5936 -15550 6336 -15540
rect 5936 -15610 5946 -15550
rect 6006 -15610 6266 -15550
rect 6326 -15610 6336 -15550
rect 5936 -15720 6336 -15610
rect 6392 -15550 6792 -15540
rect 6392 -15610 6402 -15550
rect 6462 -15610 6722 -15550
rect 6782 -15610 6792 -15550
rect 6392 -15720 6792 -15610
rect 3652 -15791 6792 -15720
rect 3652 -15900 4052 -15791
rect 3652 -15960 3662 -15900
rect 3722 -15960 3982 -15900
rect 4042 -15960 4052 -15900
rect 3652 -15970 4052 -15960
rect 4110 -15900 4510 -15791
rect 4110 -15960 4120 -15900
rect 4180 -15960 4440 -15900
rect 4500 -15960 4510 -15900
rect 4110 -15970 4510 -15960
rect 4566 -15900 4966 -15791
rect 4566 -15960 4576 -15900
rect 4636 -15960 4896 -15900
rect 4956 -15960 4966 -15900
rect 4566 -15970 4966 -15960
rect 5022 -15900 5422 -15791
rect 5022 -15960 5032 -15900
rect 5092 -15960 5352 -15900
rect 5412 -15960 5422 -15900
rect 5022 -15970 5422 -15960
rect 5480 -15900 5880 -15791
rect 5480 -15960 5490 -15900
rect 5550 -15960 5810 -15900
rect 5870 -15960 5880 -15900
rect 5480 -15970 5880 -15960
rect 5936 -15900 6336 -15791
rect 5936 -15960 5946 -15900
rect 6006 -15960 6266 -15900
rect 6326 -15960 6336 -15900
rect 5936 -15970 6336 -15960
rect 6392 -15900 6792 -15791
rect 6392 -15960 6402 -15900
rect 6462 -15960 6722 -15900
rect 6782 -15960 6792 -15900
rect 6392 -15970 6792 -15960
rect 6850 -15550 7250 -15540
rect 6850 -15610 6860 -15550
rect 6920 -15610 7180 -15550
rect 7240 -15610 7250 -15550
rect 6850 -15720 7250 -15610
rect 7306 -15550 7706 -15540
rect 7306 -15610 7316 -15550
rect 7376 -15610 7636 -15550
rect 7696 -15610 7706 -15550
rect 7306 -15720 7706 -15610
rect 7762 -15550 8162 -15540
rect 7762 -15610 7772 -15550
rect 7832 -15610 8092 -15550
rect 8152 -15610 8162 -15550
rect 7762 -15720 8162 -15610
rect 8236 -15550 8636 -15540
rect 8236 -15610 8246 -15550
rect 8306 -15610 8566 -15550
rect 8626 -15610 8636 -15550
rect 8236 -15720 8636 -15610
rect 8692 -15550 9092 -15540
rect 8692 -15610 8702 -15550
rect 8762 -15610 9022 -15550
rect 9082 -15610 9092 -15550
rect 8692 -15720 9092 -15610
rect 9150 -15550 9550 -15540
rect 9150 -15610 9160 -15550
rect 9220 -15610 9480 -15550
rect 9540 -15610 9550 -15550
rect 9150 -15720 9550 -15610
rect 9606 -15550 10006 -15540
rect 9606 -15610 9616 -15550
rect 9676 -15610 9936 -15550
rect 9996 -15610 10006 -15550
rect 9606 -15720 10006 -15610
rect 10062 -15550 10462 -15540
rect 10062 -15610 10072 -15550
rect 10132 -15610 10392 -15550
rect 10452 -15610 10462 -15550
rect 10062 -15720 10462 -15610
rect 6850 -15791 9093 -15720
rect 9150 -15791 10462 -15720
rect 6850 -15900 7250 -15791
rect 6850 -15960 6860 -15900
rect 6920 -15960 7180 -15900
rect 7240 -15960 7250 -15900
rect 6850 -15970 7250 -15960
rect 7306 -15900 7706 -15791
rect 7306 -15960 7316 -15900
rect 7376 -15960 7636 -15900
rect 7696 -15960 7706 -15900
rect 7306 -15970 7706 -15960
rect 7762 -15900 8162 -15791
rect 7762 -15960 7772 -15900
rect 7832 -15960 8092 -15900
rect 8152 -15960 8162 -15900
rect 7762 -15970 8162 -15960
rect 8236 -15900 8636 -15791
rect 8236 -15960 8246 -15900
rect 8306 -15960 8566 -15900
rect 8626 -15960 8636 -15900
rect 8236 -15970 8636 -15960
rect 8692 -15900 9092 -15791
rect 8692 -15960 8702 -15900
rect 8762 -15960 9022 -15900
rect 9082 -15960 9092 -15900
rect 8692 -15970 9092 -15960
rect 9150 -15900 9550 -15791
rect 9150 -15960 9160 -15900
rect 9220 -15960 9480 -15900
rect 9540 -15960 9550 -15900
rect 9150 -15970 9550 -15960
rect 9606 -15900 10006 -15791
rect 9606 -15960 9616 -15900
rect 9676 -15960 9936 -15900
rect 9996 -15960 10006 -15900
rect 9606 -15970 10006 -15960
rect 10062 -15900 10462 -15791
rect 10062 -15960 10072 -15900
rect 10132 -15960 10392 -15900
rect 10452 -15960 10462 -15900
rect 10062 -15970 10462 -15960
rect 10520 -15550 10920 -15540
rect 10520 -15610 10530 -15550
rect 10590 -15610 10850 -15550
rect 10910 -15610 10920 -15550
rect 10520 -15720 10920 -15610
rect 10976 -15550 11376 -15540
rect 10976 -15610 10986 -15550
rect 11046 -15610 11306 -15550
rect 11366 -15610 11376 -15550
rect 10976 -15720 11376 -15610
rect 11432 -15550 11832 -15540
rect 11432 -15610 11442 -15550
rect 11502 -15610 11762 -15550
rect 11822 -15610 11832 -15550
rect 11432 -15720 11832 -15610
rect 10520 -15791 11832 -15720
rect 10520 -15900 10920 -15791
rect 10520 -15960 10530 -15900
rect 10590 -15960 10850 -15900
rect 10910 -15960 10920 -15900
rect 10520 -15970 10920 -15960
rect 10976 -15900 11376 -15791
rect 10976 -15960 10986 -15900
rect 11046 -15960 11306 -15900
rect 11366 -15960 11376 -15900
rect 10976 -15970 11376 -15960
rect 11432 -15900 11832 -15791
rect 11432 -15960 11442 -15900
rect 11502 -15960 11762 -15900
rect 11822 -15960 11832 -15900
rect 11432 -15970 11832 -15960
rect 11890 -15550 12290 -15540
rect 11890 -15610 11900 -15550
rect 11960 -15610 12220 -15550
rect 12280 -15610 12290 -15550
rect 11890 -15720 12290 -15610
rect 12346 -15550 12746 -15540
rect 12346 -15610 12356 -15550
rect 12416 -15610 12676 -15550
rect 12736 -15610 12746 -15550
rect 12346 -15720 12746 -15610
rect 12802 -15550 13202 -15540
rect 12802 -15610 12812 -15550
rect 12872 -15610 13132 -15550
rect 13192 -15610 13202 -15550
rect 12802 -15720 13202 -15610
rect 11890 -15791 13202 -15720
rect 11890 -15900 12290 -15791
rect 11890 -15960 11900 -15900
rect 11960 -15960 12220 -15900
rect 12280 -15960 12290 -15900
rect 11890 -15970 12290 -15960
rect 12346 -15900 12746 -15791
rect 12346 -15960 12356 -15900
rect 12416 -15960 12676 -15900
rect 12736 -15960 12746 -15900
rect 12346 -15970 12746 -15960
rect 12802 -15900 13202 -15791
rect 12802 -15960 12812 -15900
rect 12872 -15960 13132 -15900
rect 13192 -15960 13202 -15900
rect 12802 -15970 13202 -15960
rect 13260 -15550 13660 -15540
rect 13260 -15610 13270 -15550
rect 13330 -15610 13590 -15550
rect 13650 -15610 13660 -15550
rect 13260 -15900 13660 -15610
rect 13260 -15960 13270 -15900
rect 13330 -15960 13590 -15900
rect 13650 -15960 13660 -15900
rect 13260 -15970 13660 -15960
rect 13716 -15550 14116 -15540
rect 13716 -15610 13726 -15550
rect 13786 -15610 14046 -15550
rect 14106 -15610 14116 -15550
rect 13716 -15900 14116 -15610
rect 13716 -15960 13726 -15900
rect 13786 -15960 14046 -15900
rect 14106 -15960 14116 -15900
rect 13716 -15970 14116 -15960
rect 14172 -15550 14572 -15540
rect 14172 -15610 14182 -15550
rect 14242 -15610 14502 -15550
rect 14562 -15610 14572 -15550
rect 14172 -15900 14572 -15610
rect 14172 -15960 14182 -15900
rect 14242 -15960 14502 -15900
rect 14562 -15960 14572 -15900
rect 14172 -15970 14572 -15960
rect 14630 -15550 15030 -15540
rect 14630 -15610 14640 -15550
rect 14700 -15610 14960 -15550
rect 15020 -15610 15030 -15550
rect 14630 -15720 15030 -15610
rect 15086 -15550 15486 -15540
rect 15086 -15610 15096 -15550
rect 15156 -15610 15416 -15550
rect 15476 -15610 15486 -15550
rect 15086 -15719 15486 -15610
rect 15086 -15720 15720 -15719
rect 14630 -15790 15720 -15720
rect 14630 -15791 15486 -15790
rect 14630 -15900 15030 -15791
rect 14630 -15960 14640 -15900
rect 14700 -15960 14960 -15900
rect 15020 -15960 15030 -15900
rect 14630 -15970 15030 -15960
rect 15086 -15900 15486 -15791
rect 15086 -15960 15096 -15900
rect 15156 -15960 15416 -15900
rect 15476 -15960 15486 -15900
rect 15086 -15970 15486 -15960
rect 66 -16042 80 -15970
rect 456 -16042 526 -15970
rect 912 -16042 983 -15970
rect 1370 -16042 1441 -15970
rect 1826 -16042 1897 -15970
rect 2282 -16042 2353 -15970
rect 2740 -16042 2811 -15970
rect 3196 -16042 3267 -15970
rect 3652 -16042 3723 -15970
rect 4110 -16042 4181 -15970
rect 4566 -16042 4637 -15970
rect 5022 -16042 5093 -15970
rect 5480 -16042 5551 -15970
rect 5936 -16042 6007 -15970
rect 6392 -16042 6463 -15970
rect 6850 -16042 6921 -15970
rect 7306 -16042 7377 -15970
rect 7762 -16042 7833 -15970
rect 8236 -16042 8307 -15970
rect 8692 -16042 8763 -15970
rect 9150 -16042 9221 -15970
rect 9606 -16042 9677 -15970
rect 10062 -16042 10133 -15970
rect 10520 -16042 10591 -15970
rect 10976 -16042 11047 -15970
rect 11432 -16042 11503 -15970
rect 11890 -16042 11961 -15970
rect 12346 -16042 12417 -15970
rect 12802 -16042 12873 -15970
rect 13260 -16042 13331 -15970
rect 13716 -16042 13787 -15970
rect 14172 -16042 14243 -15970
rect 66 -16052 400 -16042
rect 0 -16112 10 -16052
rect 70 -16112 330 -16052
rect 390 -16112 400 -16052
rect 0 -16402 14 -16112
rect 66 -16402 400 -16112
rect 0 -16462 10 -16402
rect 70 -16462 330 -16402
rect 390 -16462 400 -16402
rect 0 -16544 14 -16462
rect 66 -16472 400 -16462
rect 456 -16052 856 -16042
rect 456 -16112 466 -16052
rect 526 -16112 786 -16052
rect 846 -16112 856 -16052
rect 456 -16221 856 -16112
rect 912 -16052 1312 -16042
rect 912 -16112 922 -16052
rect 982 -16112 1242 -16052
rect 1302 -16112 1312 -16052
rect 912 -16221 1312 -16112
rect 1370 -16052 1770 -16042
rect 1370 -16112 1380 -16052
rect 1440 -16112 1700 -16052
rect 1760 -16112 1770 -16052
rect 1370 -16221 1770 -16112
rect 1826 -16052 2226 -16042
rect 1826 -16112 1836 -16052
rect 1896 -16112 2156 -16052
rect 2216 -16112 2226 -16052
rect 1826 -16221 2226 -16112
rect 2282 -16052 2682 -16042
rect 2282 -16112 2292 -16052
rect 2352 -16112 2612 -16052
rect 2672 -16112 2682 -16052
rect 2282 -16221 2682 -16112
rect 2740 -16052 3140 -16042
rect 2740 -16112 2750 -16052
rect 2810 -16112 3070 -16052
rect 3130 -16112 3140 -16052
rect 2740 -16221 3140 -16112
rect 3196 -16052 3596 -16042
rect 3196 -16112 3206 -16052
rect 3266 -16112 3526 -16052
rect 3586 -16112 3596 -16052
rect 3196 -16221 3596 -16112
rect 456 -16291 3596 -16221
rect 456 -16292 2682 -16291
rect 456 -16402 856 -16292
rect 456 -16462 466 -16402
rect 526 -16462 786 -16402
rect 846 -16462 856 -16402
rect 456 -16472 856 -16462
rect 912 -16402 1312 -16292
rect 912 -16462 922 -16402
rect 982 -16462 1242 -16402
rect 1302 -16462 1312 -16402
rect 912 -16472 1312 -16462
rect 1370 -16402 1770 -16292
rect 1370 -16462 1380 -16402
rect 1440 -16462 1700 -16402
rect 1760 -16462 1770 -16402
rect 1370 -16472 1770 -16462
rect 1826 -16402 2226 -16292
rect 1826 -16462 1836 -16402
rect 1896 -16462 2156 -16402
rect 2216 -16462 2226 -16402
rect 1826 -16472 2226 -16462
rect 2282 -16402 2682 -16292
rect 2282 -16462 2292 -16402
rect 2352 -16462 2612 -16402
rect 2672 -16462 2682 -16402
rect 2282 -16472 2682 -16462
rect 2740 -16292 3596 -16291
rect 2740 -16402 3140 -16292
rect 2740 -16462 2750 -16402
rect 2810 -16462 3070 -16402
rect 3130 -16462 3140 -16402
rect 2740 -16472 3140 -16462
rect 3196 -16402 3596 -16292
rect 3196 -16462 3206 -16402
rect 3266 -16462 3526 -16402
rect 3586 -16462 3596 -16402
rect 3196 -16472 3596 -16462
rect 3652 -16052 4052 -16042
rect 3652 -16112 3662 -16052
rect 3722 -16112 3982 -16052
rect 4042 -16112 4052 -16052
rect 3652 -16221 4052 -16112
rect 4110 -16052 4510 -16042
rect 4110 -16112 4120 -16052
rect 4180 -16112 4440 -16052
rect 4500 -16112 4510 -16052
rect 4110 -16221 4510 -16112
rect 4566 -16052 4966 -16042
rect 4566 -16112 4576 -16052
rect 4636 -16112 4896 -16052
rect 4956 -16112 4966 -16052
rect 4566 -16221 4966 -16112
rect 5022 -16052 5422 -16042
rect 5022 -16112 5032 -16052
rect 5092 -16112 5352 -16052
rect 5412 -16112 5422 -16052
rect 5022 -16221 5422 -16112
rect 5480 -16052 5880 -16042
rect 5480 -16112 5490 -16052
rect 5550 -16112 5810 -16052
rect 5870 -16112 5880 -16052
rect 5480 -16221 5880 -16112
rect 5936 -16052 6336 -16042
rect 5936 -16112 5946 -16052
rect 6006 -16112 6266 -16052
rect 6326 -16112 6336 -16052
rect 5936 -16221 6336 -16112
rect 6392 -16052 6792 -16042
rect 6392 -16112 6402 -16052
rect 6462 -16112 6722 -16052
rect 6782 -16112 6792 -16052
rect 6392 -16221 6792 -16112
rect 3652 -16292 6792 -16221
rect 3652 -16402 4052 -16292
rect 3652 -16462 3662 -16402
rect 3722 -16462 3982 -16402
rect 4042 -16462 4052 -16402
rect 3652 -16472 4052 -16462
rect 4110 -16402 4510 -16292
rect 4110 -16462 4120 -16402
rect 4180 -16462 4440 -16402
rect 4500 -16462 4510 -16402
rect 4110 -16472 4510 -16462
rect 4566 -16402 4966 -16292
rect 4566 -16462 4576 -16402
rect 4636 -16462 4896 -16402
rect 4956 -16462 4966 -16402
rect 4566 -16472 4966 -16462
rect 5022 -16402 5422 -16292
rect 5022 -16462 5032 -16402
rect 5092 -16462 5352 -16402
rect 5412 -16462 5422 -16402
rect 5022 -16472 5422 -16462
rect 5480 -16402 5880 -16292
rect 5480 -16462 5490 -16402
rect 5550 -16462 5810 -16402
rect 5870 -16462 5880 -16402
rect 5480 -16472 5880 -16462
rect 5936 -16402 6336 -16292
rect 5936 -16462 5946 -16402
rect 6006 -16462 6266 -16402
rect 6326 -16462 6336 -16402
rect 5936 -16472 6336 -16462
rect 6392 -16402 6792 -16292
rect 6392 -16462 6402 -16402
rect 6462 -16462 6722 -16402
rect 6782 -16462 6792 -16402
rect 6392 -16472 6792 -16462
rect 6850 -16052 7250 -16042
rect 6850 -16112 6860 -16052
rect 6920 -16112 7180 -16052
rect 7240 -16112 7250 -16052
rect 6850 -16221 7250 -16112
rect 7306 -16052 7706 -16042
rect 7306 -16112 7316 -16052
rect 7376 -16112 7636 -16052
rect 7696 -16112 7706 -16052
rect 7306 -16221 7706 -16112
rect 7762 -16052 8162 -16042
rect 7762 -16112 7772 -16052
rect 7832 -16112 8092 -16052
rect 8152 -16112 8162 -16052
rect 7762 -16221 8162 -16112
rect 8236 -16052 8636 -16042
rect 8236 -16112 8246 -16052
rect 8306 -16112 8566 -16052
rect 8626 -16112 8636 -16052
rect 8236 -16221 8636 -16112
rect 8692 -16052 9092 -16042
rect 8692 -16112 8702 -16052
rect 8762 -16112 9022 -16052
rect 9082 -16112 9092 -16052
rect 8692 -16221 9092 -16112
rect 9150 -16052 9550 -16042
rect 9150 -16112 9160 -16052
rect 9220 -16112 9480 -16052
rect 9540 -16112 9550 -16052
rect 9150 -16221 9550 -16112
rect 9606 -16052 10006 -16042
rect 9606 -16112 9616 -16052
rect 9676 -16112 9936 -16052
rect 9996 -16112 10006 -16052
rect 9606 -16221 10006 -16112
rect 10062 -16052 10462 -16042
rect 10062 -16112 10072 -16052
rect 10132 -16112 10392 -16052
rect 10452 -16112 10462 -16052
rect 10062 -16221 10462 -16112
rect 6850 -16292 9093 -16221
rect 9150 -16292 10462 -16221
rect 6850 -16402 7250 -16292
rect 6850 -16462 6860 -16402
rect 6920 -16462 7180 -16402
rect 7240 -16462 7250 -16402
rect 6850 -16472 7250 -16462
rect 7306 -16402 7706 -16292
rect 7306 -16462 7316 -16402
rect 7376 -16462 7636 -16402
rect 7696 -16462 7706 -16402
rect 7306 -16472 7706 -16462
rect 7762 -16402 8162 -16292
rect 7762 -16462 7772 -16402
rect 7832 -16462 8092 -16402
rect 8152 -16462 8162 -16402
rect 7762 -16472 8162 -16462
rect 8236 -16402 8636 -16292
rect 8236 -16462 8246 -16402
rect 8306 -16462 8566 -16402
rect 8626 -16462 8636 -16402
rect 8236 -16472 8636 -16462
rect 8692 -16402 9092 -16292
rect 8692 -16462 8702 -16402
rect 8762 -16462 9022 -16402
rect 9082 -16462 9092 -16402
rect 8692 -16472 9092 -16462
rect 9150 -16402 9550 -16292
rect 9150 -16462 9160 -16402
rect 9220 -16462 9480 -16402
rect 9540 -16462 9550 -16402
rect 9150 -16472 9550 -16462
rect 9606 -16402 10006 -16292
rect 9606 -16462 9616 -16402
rect 9676 -16462 9936 -16402
rect 9996 -16462 10006 -16402
rect 9606 -16472 10006 -16462
rect 10062 -16402 10462 -16292
rect 10062 -16462 10072 -16402
rect 10132 -16462 10392 -16402
rect 10452 -16462 10462 -16402
rect 10062 -16472 10462 -16462
rect 10520 -16052 10920 -16042
rect 10520 -16112 10530 -16052
rect 10590 -16112 10850 -16052
rect 10910 -16112 10920 -16052
rect 10520 -16221 10920 -16112
rect 10976 -16052 11376 -16042
rect 10976 -16112 10986 -16052
rect 11046 -16112 11306 -16052
rect 11366 -16112 11376 -16052
rect 10976 -16221 11376 -16112
rect 11432 -16052 11832 -16042
rect 11432 -16112 11442 -16052
rect 11502 -16112 11762 -16052
rect 11822 -16112 11832 -16052
rect 11432 -16221 11832 -16112
rect 10520 -16292 11832 -16221
rect 10520 -16402 10920 -16292
rect 10520 -16462 10530 -16402
rect 10590 -16462 10850 -16402
rect 10910 -16462 10920 -16402
rect 10520 -16472 10920 -16462
rect 10976 -16402 11376 -16292
rect 10976 -16462 10986 -16402
rect 11046 -16462 11306 -16402
rect 11366 -16462 11376 -16402
rect 10976 -16472 11376 -16462
rect 11432 -16402 11832 -16292
rect 11432 -16462 11442 -16402
rect 11502 -16462 11762 -16402
rect 11822 -16462 11832 -16402
rect 11432 -16472 11832 -16462
rect 11890 -16052 12290 -16042
rect 11890 -16112 11900 -16052
rect 11960 -16112 12220 -16052
rect 12280 -16112 12290 -16052
rect 11890 -16221 12290 -16112
rect 12346 -16052 12746 -16042
rect 12346 -16112 12356 -16052
rect 12416 -16112 12676 -16052
rect 12736 -16112 12746 -16052
rect 12346 -16221 12746 -16112
rect 12802 -16052 13202 -16042
rect 12802 -16112 12812 -16052
rect 12872 -16112 13132 -16052
rect 13192 -16112 13202 -16052
rect 12802 -16221 13202 -16112
rect 11890 -16292 13202 -16221
rect 11890 -16402 12290 -16292
rect 11890 -16462 11900 -16402
rect 11960 -16462 12220 -16402
rect 12280 -16462 12290 -16402
rect 11890 -16472 12290 -16462
rect 12346 -16402 12746 -16292
rect 12346 -16462 12356 -16402
rect 12416 -16462 12676 -16402
rect 12736 -16462 12746 -16402
rect 12346 -16472 12746 -16462
rect 12802 -16402 13202 -16292
rect 12802 -16462 12812 -16402
rect 12872 -16462 13132 -16402
rect 13192 -16462 13202 -16402
rect 12802 -16472 13202 -16462
rect 13260 -16052 13660 -16042
rect 13260 -16112 13270 -16052
rect 13330 -16112 13590 -16052
rect 13650 -16112 13660 -16052
rect 13260 -16402 13660 -16112
rect 13260 -16462 13270 -16402
rect 13330 -16462 13590 -16402
rect 13650 -16462 13660 -16402
rect 13260 -16472 13660 -16462
rect 13716 -16052 14116 -16042
rect 13716 -16112 13726 -16052
rect 13786 -16112 14046 -16052
rect 14106 -16112 14116 -16052
rect 13716 -16402 14116 -16112
rect 13716 -16462 13726 -16402
rect 13786 -16462 14046 -16402
rect 14106 -16462 14116 -16402
rect 13716 -16472 14116 -16462
rect 14172 -16052 14572 -16042
rect 14172 -16112 14182 -16052
rect 14242 -16112 14502 -16052
rect 14562 -16112 14572 -16052
rect 14172 -16402 14572 -16112
rect 14172 -16462 14182 -16402
rect 14242 -16462 14502 -16402
rect 14562 -16462 14572 -16402
rect 14172 -16472 14572 -16462
rect 14630 -16052 15030 -16042
rect 14630 -16112 14640 -16052
rect 14700 -16112 14960 -16052
rect 15020 -16112 15030 -16052
rect 14630 -16221 15030 -16112
rect 15086 -16052 15486 -16042
rect 15086 -16112 15096 -16052
rect 15156 -16112 15416 -16052
rect 15476 -16112 15486 -16052
rect 15086 -16221 15486 -16112
rect 14630 -16222 15486 -16221
rect 14630 -16292 15720 -16222
rect 14630 -16402 15030 -16292
rect 14630 -16462 14640 -16402
rect 14700 -16462 14960 -16402
rect 15020 -16462 15030 -16402
rect 14630 -16472 15030 -16462
rect 15086 -16293 15720 -16292
rect 15086 -16402 15486 -16293
rect 15086 -16462 15096 -16402
rect 15156 -16462 15416 -16402
rect 15476 -16462 15486 -16402
rect 15086 -16472 15486 -16462
rect 66 -16534 80 -16472
rect 456 -16534 527 -16472
rect 912 -16534 983 -16472
rect 1370 -16534 1441 -16472
rect 1826 -16534 1897 -16472
rect 2282 -16534 2353 -16472
rect 2740 -16534 2810 -16472
rect 3196 -16534 3266 -16472
rect 3652 -16534 3722 -16472
rect 4110 -16534 4180 -16472
rect 4566 -16534 4636 -16472
rect 5022 -16534 5092 -16472
rect 5480 -16534 5550 -16472
rect 5936 -16534 6006 -16472
rect 6392 -16534 6462 -16472
rect 7306 -16534 7376 -16472
rect 7762 -16534 7832 -16472
rect 8236 -16534 8306 -16472
rect 8692 -16534 8762 -16472
rect 9150 -16534 9220 -16472
rect 9606 -16534 9676 -16472
rect 10062 -16534 10132 -16472
rect 10976 -16534 11046 -16472
rect 11432 -16534 11502 -16472
rect 11890 -16534 11960 -16472
rect 12346 -16534 12416 -16472
rect 12802 -16534 12872 -16472
rect 13260 -16534 13330 -16472
rect 13716 -16534 13786 -16472
rect 14172 -16534 14242 -16472
rect 66 -16544 400 -16534
rect 0 -16604 10 -16544
rect 70 -16604 330 -16544
rect 390 -16604 400 -16544
rect 0 -16894 14 -16604
rect 66 -16894 400 -16604
rect 0 -16954 10 -16894
rect 70 -16954 330 -16894
rect 390 -16954 400 -16894
rect 0 -17041 14 -16954
rect 66 -16964 400 -16954
rect 456 -16544 856 -16534
rect 456 -16604 466 -16544
rect 526 -16604 786 -16544
rect 846 -16604 856 -16544
rect 456 -16712 856 -16604
rect 912 -16544 1312 -16534
rect 912 -16604 922 -16544
rect 982 -16604 1242 -16544
rect 1302 -16604 1312 -16544
rect 912 -16712 1312 -16604
rect 1370 -16544 1770 -16534
rect 1370 -16604 1380 -16544
rect 1440 -16604 1700 -16544
rect 1760 -16604 1770 -16544
rect 1370 -16712 1770 -16604
rect 1826 -16544 2226 -16534
rect 1826 -16604 1836 -16544
rect 1896 -16604 2156 -16544
rect 2216 -16604 2226 -16544
rect 1826 -16712 2226 -16604
rect 2282 -16544 2682 -16534
rect 2282 -16604 2292 -16544
rect 2352 -16604 2612 -16544
rect 2672 -16604 2682 -16544
rect 2282 -16712 2682 -16604
rect 2740 -16544 3140 -16534
rect 2740 -16604 2750 -16544
rect 2810 -16604 3070 -16544
rect 3130 -16604 3140 -16544
rect 2740 -16712 3140 -16604
rect 3196 -16544 3596 -16534
rect 3196 -16604 3206 -16544
rect 3266 -16604 3526 -16544
rect 3586 -16604 3596 -16544
rect 3196 -16712 3596 -16604
rect 456 -16782 3596 -16712
rect 456 -16784 2682 -16782
rect 456 -16894 856 -16784
rect 456 -16954 466 -16894
rect 526 -16954 786 -16894
rect 846 -16954 856 -16894
rect 456 -16964 856 -16954
rect 912 -16894 1312 -16784
rect 912 -16954 922 -16894
rect 982 -16954 1242 -16894
rect 1302 -16954 1312 -16894
rect 912 -16964 1312 -16954
rect 1370 -16894 1770 -16784
rect 1370 -16954 1380 -16894
rect 1440 -16954 1700 -16894
rect 1760 -16954 1770 -16894
rect 1370 -16964 1770 -16954
rect 1826 -16894 2226 -16784
rect 1826 -16954 1836 -16894
rect 1896 -16954 2156 -16894
rect 2216 -16954 2226 -16894
rect 1826 -16964 2226 -16954
rect 2282 -16894 2682 -16784
rect 2282 -16954 2292 -16894
rect 2352 -16954 2612 -16894
rect 2672 -16954 2682 -16894
rect 2282 -16964 2682 -16954
rect 2740 -16784 3596 -16782
rect 2740 -16894 3140 -16784
rect 2740 -16954 2750 -16894
rect 2810 -16954 3070 -16894
rect 3130 -16954 3140 -16894
rect 2740 -16964 3140 -16954
rect 3196 -16894 3596 -16784
rect 3196 -16954 3206 -16894
rect 3266 -16954 3526 -16894
rect 3586 -16954 3596 -16894
rect 3196 -16964 3596 -16954
rect 3652 -16544 4052 -16534
rect 3652 -16604 3662 -16544
rect 3722 -16604 3982 -16544
rect 4042 -16604 4052 -16544
rect 3652 -16712 4052 -16604
rect 4110 -16544 4510 -16534
rect 4110 -16604 4120 -16544
rect 4180 -16604 4440 -16544
rect 4500 -16604 4510 -16544
rect 4110 -16712 4510 -16604
rect 4566 -16544 4966 -16534
rect 4566 -16604 4576 -16544
rect 4636 -16604 4896 -16544
rect 4956 -16604 4966 -16544
rect 4566 -16712 4966 -16604
rect 5022 -16544 5422 -16534
rect 5022 -16604 5032 -16544
rect 5092 -16604 5352 -16544
rect 5412 -16604 5422 -16544
rect 5022 -16712 5422 -16604
rect 5480 -16544 5880 -16534
rect 5480 -16604 5490 -16544
rect 5550 -16604 5810 -16544
rect 5870 -16604 5880 -16544
rect 5480 -16712 5880 -16604
rect 5936 -16544 6336 -16534
rect 5936 -16604 5946 -16544
rect 6006 -16604 6266 -16544
rect 6326 -16604 6336 -16544
rect 5936 -16712 6336 -16604
rect 6392 -16544 6792 -16534
rect 6392 -16604 6402 -16544
rect 6462 -16604 6722 -16544
rect 6782 -16604 6792 -16544
rect 6392 -16712 6792 -16604
rect 6850 -16544 7250 -16534
rect 6850 -16604 6860 -16544
rect 6920 -16604 7180 -16544
rect 7240 -16604 7250 -16544
rect 6850 -16712 7250 -16604
rect 3652 -16784 7250 -16712
rect 3652 -16894 4052 -16784
rect 3652 -16954 3662 -16894
rect 3722 -16954 3982 -16894
rect 4042 -16954 4052 -16894
rect 3652 -16964 4052 -16954
rect 4110 -16894 4510 -16784
rect 4110 -16954 4120 -16894
rect 4180 -16954 4440 -16894
rect 4500 -16954 4510 -16894
rect 4110 -16964 4510 -16954
rect 4566 -16894 4966 -16784
rect 4566 -16954 4576 -16894
rect 4636 -16954 4896 -16894
rect 4956 -16954 4966 -16894
rect 4566 -16964 4966 -16954
rect 5022 -16894 5422 -16784
rect 5022 -16954 5032 -16894
rect 5092 -16954 5352 -16894
rect 5412 -16954 5422 -16894
rect 5022 -16964 5422 -16954
rect 5480 -16894 5880 -16784
rect 5480 -16954 5490 -16894
rect 5550 -16954 5810 -16894
rect 5870 -16954 5880 -16894
rect 5480 -16964 5880 -16954
rect 5936 -16894 6336 -16784
rect 5936 -16954 5946 -16894
rect 6006 -16954 6266 -16894
rect 6326 -16954 6336 -16894
rect 5936 -16964 6336 -16954
rect 6392 -16894 6792 -16784
rect 6392 -16954 6402 -16894
rect 6462 -16954 6722 -16894
rect 6782 -16954 6792 -16894
rect 6392 -16964 6792 -16954
rect 6850 -16894 7250 -16784
rect 6850 -16954 6860 -16894
rect 6920 -16954 7180 -16894
rect 7240 -16954 7250 -16894
rect 6850 -16964 7250 -16954
rect 7306 -16544 7706 -16534
rect 7306 -16604 7316 -16544
rect 7376 -16604 7636 -16544
rect 7696 -16604 7706 -16544
rect 7306 -16712 7706 -16604
rect 7762 -16544 8162 -16534
rect 7762 -16604 7772 -16544
rect 7832 -16604 8092 -16544
rect 8152 -16604 8162 -16544
rect 7762 -16712 8162 -16604
rect 8236 -16544 8636 -16534
rect 8236 -16604 8246 -16544
rect 8306 -16604 8566 -16544
rect 8626 -16604 8636 -16544
rect 8236 -16712 8636 -16604
rect 8692 -16544 9092 -16534
rect 8692 -16604 8702 -16544
rect 8762 -16604 9022 -16544
rect 9082 -16604 9092 -16544
rect 8692 -16712 9092 -16604
rect 9150 -16544 9550 -16534
rect 9150 -16604 9160 -16544
rect 9220 -16604 9480 -16544
rect 9540 -16604 9550 -16544
rect 9150 -16712 9550 -16604
rect 9606 -16544 10006 -16534
rect 9606 -16604 9616 -16544
rect 9676 -16604 9936 -16544
rect 9996 -16604 10006 -16544
rect 9606 -16712 10006 -16604
rect 10062 -16544 10462 -16534
rect 10062 -16604 10072 -16544
rect 10132 -16604 10392 -16544
rect 10452 -16604 10462 -16544
rect 10062 -16712 10462 -16604
rect 10520 -16544 10920 -16534
rect 10520 -16604 10530 -16544
rect 10590 -16604 10850 -16544
rect 10910 -16604 10920 -16544
rect 10520 -16712 10920 -16604
rect 7306 -16784 9093 -16712
rect 9150 -16782 10920 -16712
rect 9150 -16784 10462 -16782
rect 7306 -16894 7706 -16784
rect 7306 -16954 7316 -16894
rect 7376 -16954 7636 -16894
rect 7696 -16954 7706 -16894
rect 7306 -16964 7706 -16954
rect 7762 -16894 8162 -16784
rect 7762 -16954 7772 -16894
rect 7832 -16954 8092 -16894
rect 8152 -16954 8162 -16894
rect 7762 -16964 8162 -16954
rect 8236 -16894 8636 -16784
rect 8236 -16954 8246 -16894
rect 8306 -16954 8566 -16894
rect 8626 -16954 8636 -16894
rect 8236 -16964 8636 -16954
rect 8692 -16894 9092 -16784
rect 8692 -16954 8702 -16894
rect 8762 -16954 9022 -16894
rect 9082 -16954 9092 -16894
rect 8692 -16964 9092 -16954
rect 9150 -16894 9550 -16784
rect 9150 -16954 9160 -16894
rect 9220 -16954 9480 -16894
rect 9540 -16954 9550 -16894
rect 9150 -16964 9550 -16954
rect 9606 -16894 10006 -16784
rect 9606 -16954 9616 -16894
rect 9676 -16954 9936 -16894
rect 9996 -16954 10006 -16894
rect 9606 -16964 10006 -16954
rect 10062 -16894 10462 -16784
rect 10062 -16954 10072 -16894
rect 10132 -16954 10392 -16894
rect 10452 -16954 10462 -16894
rect 10062 -16964 10462 -16954
rect 10520 -16894 10920 -16782
rect 10520 -16954 10530 -16894
rect 10590 -16954 10850 -16894
rect 10910 -16954 10920 -16894
rect 10520 -16964 10920 -16954
rect 10976 -16544 11376 -16534
rect 10976 -16604 10986 -16544
rect 11046 -16604 11306 -16544
rect 11366 -16604 11376 -16544
rect 10976 -16712 11376 -16604
rect 11432 -16544 11832 -16534
rect 11432 -16604 11442 -16544
rect 11502 -16604 11762 -16544
rect 11822 -16604 11832 -16544
rect 11432 -16712 11832 -16604
rect 10976 -16784 11832 -16712
rect 10976 -16894 11376 -16784
rect 10976 -16954 10986 -16894
rect 11046 -16954 11306 -16894
rect 11366 -16954 11376 -16894
rect 10976 -16964 11376 -16954
rect 11432 -16894 11832 -16784
rect 11432 -16954 11442 -16894
rect 11502 -16954 11762 -16894
rect 11822 -16954 11832 -16894
rect 11432 -16964 11832 -16954
rect 11890 -16544 12290 -16534
rect 11890 -16604 11900 -16544
rect 11960 -16604 12220 -16544
rect 12280 -16604 12290 -16544
rect 11890 -16712 12290 -16604
rect 12346 -16544 12746 -16534
rect 12346 -16604 12356 -16544
rect 12416 -16604 12676 -16544
rect 12736 -16604 12746 -16544
rect 12346 -16712 12746 -16604
rect 12802 -16544 13202 -16534
rect 12802 -16604 12812 -16544
rect 12872 -16604 13132 -16544
rect 13192 -16604 13202 -16544
rect 12802 -16712 13202 -16604
rect 11890 -16784 13202 -16712
rect 11890 -16894 12290 -16784
rect 11890 -16954 11900 -16894
rect 11960 -16954 12220 -16894
rect 12280 -16954 12290 -16894
rect 11890 -16964 12290 -16954
rect 12346 -16894 12746 -16784
rect 12346 -16954 12356 -16894
rect 12416 -16954 12676 -16894
rect 12736 -16954 12746 -16894
rect 12346 -16964 12746 -16954
rect 12802 -16894 13202 -16784
rect 12802 -16954 12812 -16894
rect 12872 -16954 13132 -16894
rect 13192 -16954 13202 -16894
rect 12802 -16964 13202 -16954
rect 13260 -16544 13660 -16534
rect 13260 -16604 13270 -16544
rect 13330 -16604 13590 -16544
rect 13650 -16604 13660 -16544
rect 13260 -16894 13660 -16604
rect 13260 -16954 13270 -16894
rect 13330 -16954 13590 -16894
rect 13650 -16954 13660 -16894
rect 13260 -16964 13660 -16954
rect 13716 -16544 14116 -16534
rect 13716 -16604 13726 -16544
rect 13786 -16604 14046 -16544
rect 14106 -16604 14116 -16544
rect 13716 -16894 14116 -16604
rect 13716 -16954 13726 -16894
rect 13786 -16954 14046 -16894
rect 14106 -16954 14116 -16894
rect 13716 -16964 14116 -16954
rect 14172 -16544 14572 -16534
rect 14172 -16604 14182 -16544
rect 14242 -16604 14502 -16544
rect 14562 -16604 14572 -16544
rect 14172 -16714 14572 -16604
rect 14630 -16544 15030 -16534
rect 14630 -16604 14640 -16544
rect 14700 -16604 14960 -16544
rect 15020 -16604 15030 -16544
rect 14630 -16712 15030 -16604
rect 15086 -16544 15486 -16534
rect 15086 -16604 15096 -16544
rect 15156 -16604 15416 -16544
rect 15476 -16604 15486 -16544
rect 15086 -16712 15486 -16604
rect 14630 -16713 15486 -16712
rect 14630 -16714 15720 -16713
rect 14172 -16778 15720 -16714
rect 14172 -16894 14572 -16778
rect 14172 -16954 14182 -16894
rect 14242 -16954 14502 -16894
rect 14562 -16954 14572 -16894
rect 14172 -16964 14572 -16954
rect 14630 -16784 15720 -16778
rect 14630 -16894 15030 -16784
rect 14630 -16954 14640 -16894
rect 14700 -16954 14960 -16894
rect 15020 -16954 15030 -16894
rect 14630 -16964 15030 -16954
rect 15086 -16894 15486 -16784
rect 15086 -16954 15096 -16894
rect 15156 -16954 15416 -16894
rect 15476 -16954 15486 -16894
rect 15086 -16964 15486 -16954
rect 66 -17031 80 -16964
rect 456 -16965 527 -16964
rect 457 -17031 527 -16965
rect 913 -17031 984 -16964
rect 1371 -17031 1442 -16964
rect 1827 -17031 1898 -16964
rect 2283 -17031 2354 -16964
rect 2741 -17031 2812 -16964
rect 3197 -17031 3268 -16964
rect 3653 -17031 3724 -16964
rect 4111 -17031 4182 -16964
rect 4567 -17031 4638 -16964
rect 5023 -17031 5094 -16964
rect 5481 -17031 5552 -16964
rect 5937 -17031 6008 -16964
rect 6393 -17031 6464 -16964
rect 6851 -17031 6922 -16964
rect 7307 -17031 7378 -16964
rect 7763 -17031 7834 -16964
rect 8237 -17031 8308 -16964
rect 8693 -17031 8764 -16964
rect 9151 -17031 9222 -16964
rect 9607 -17031 9678 -16964
rect 10063 -17031 10134 -16964
rect 10521 -17031 10592 -16964
rect 10977 -17031 11048 -16964
rect 11433 -17031 11504 -16964
rect 12347 -17031 12418 -16964
rect 12803 -17031 12874 -16964
rect 13261 -17031 13332 -16964
rect 13717 -17031 13788 -16964
rect 66 -17041 400 -17031
rect 0 -17101 11 -17041
rect 71 -17101 331 -17041
rect 391 -17101 400 -17041
rect 0 -17391 14 -17101
rect 66 -17391 400 -17101
rect 0 -17451 11 -17391
rect 71 -17451 331 -17391
rect 391 -17451 400 -17391
rect 0 -17533 14 -17451
rect 66 -17461 400 -17451
rect 457 -17041 857 -17031
rect 457 -17101 467 -17041
rect 527 -17101 787 -17041
rect 847 -17101 857 -17041
rect 457 -17211 857 -17101
rect 913 -17041 1313 -17031
rect 913 -17101 923 -17041
rect 983 -17101 1243 -17041
rect 1303 -17101 1313 -17041
rect 913 -17211 1313 -17101
rect 1371 -17041 1771 -17031
rect 1371 -17101 1381 -17041
rect 1441 -17101 1701 -17041
rect 1761 -17101 1771 -17041
rect 1371 -17211 1771 -17101
rect 1827 -17041 2227 -17031
rect 1827 -17101 1837 -17041
rect 1897 -17101 2157 -17041
rect 2217 -17101 2227 -17041
rect 1827 -17211 2227 -17101
rect 2283 -17041 2683 -17031
rect 2283 -17101 2293 -17041
rect 2353 -17101 2613 -17041
rect 2673 -17101 2683 -17041
rect 2283 -17211 2683 -17101
rect 2741 -17041 3141 -17031
rect 2741 -17101 2751 -17041
rect 2811 -17101 3071 -17041
rect 3131 -17101 3141 -17041
rect 2741 -17211 3141 -17101
rect 3197 -17041 3597 -17031
rect 3197 -17101 3207 -17041
rect 3267 -17101 3527 -17041
rect 3587 -17101 3597 -17041
rect 3197 -17211 3597 -17101
rect 457 -17281 3597 -17211
rect 457 -17391 857 -17281
rect 457 -17451 467 -17391
rect 527 -17451 787 -17391
rect 847 -17451 857 -17391
rect 457 -17461 857 -17451
rect 913 -17391 1313 -17281
rect 913 -17451 923 -17391
rect 983 -17451 1243 -17391
rect 1303 -17451 1313 -17391
rect 913 -17461 1313 -17451
rect 1371 -17391 1771 -17281
rect 1371 -17451 1381 -17391
rect 1441 -17451 1701 -17391
rect 1761 -17451 1771 -17391
rect 1371 -17461 1771 -17451
rect 1827 -17391 2227 -17281
rect 1827 -17451 1837 -17391
rect 1897 -17451 2157 -17391
rect 2217 -17451 2227 -17391
rect 1827 -17461 2227 -17451
rect 2283 -17391 2683 -17281
rect 2283 -17451 2293 -17391
rect 2353 -17451 2613 -17391
rect 2673 -17451 2683 -17391
rect 2283 -17461 2683 -17451
rect 2741 -17391 3141 -17281
rect 2741 -17451 2751 -17391
rect 2811 -17451 3071 -17391
rect 3131 -17451 3141 -17391
rect 2741 -17461 3141 -17451
rect 3197 -17391 3597 -17281
rect 3197 -17451 3207 -17391
rect 3267 -17451 3527 -17391
rect 3587 -17451 3597 -17391
rect 3197 -17461 3597 -17451
rect 3653 -17041 4053 -17031
rect 3653 -17101 3663 -17041
rect 3723 -17101 3983 -17041
rect 4043 -17101 4053 -17041
rect 3653 -17211 4053 -17101
rect 4111 -17041 4511 -17031
rect 4111 -17101 4121 -17041
rect 4181 -17101 4441 -17041
rect 4501 -17101 4511 -17041
rect 4111 -17211 4511 -17101
rect 4567 -17041 4967 -17031
rect 4567 -17101 4577 -17041
rect 4637 -17101 4897 -17041
rect 4957 -17101 4967 -17041
rect 4567 -17211 4967 -17101
rect 5023 -17041 5423 -17031
rect 5023 -17101 5033 -17041
rect 5093 -17101 5353 -17041
rect 5413 -17101 5423 -17041
rect 5023 -17211 5423 -17101
rect 5481 -17041 5881 -17031
rect 5481 -17101 5491 -17041
rect 5551 -17101 5811 -17041
rect 5871 -17101 5881 -17041
rect 5481 -17211 5881 -17101
rect 5937 -17041 6337 -17031
rect 5937 -17101 5947 -17041
rect 6007 -17101 6267 -17041
rect 6327 -17101 6337 -17041
rect 5937 -17211 6337 -17101
rect 6393 -17041 6793 -17031
rect 6393 -17101 6403 -17041
rect 6463 -17101 6723 -17041
rect 6783 -17101 6793 -17041
rect 6393 -17211 6793 -17101
rect 6851 -17041 7251 -17031
rect 6851 -17101 6861 -17041
rect 6921 -17101 7181 -17041
rect 7241 -17101 7251 -17041
rect 6851 -17211 7251 -17101
rect 3653 -17281 7251 -17211
rect 3653 -17391 4053 -17281
rect 3653 -17451 3663 -17391
rect 3723 -17451 3983 -17391
rect 4043 -17451 4053 -17391
rect 3653 -17461 4053 -17451
rect 4111 -17391 4511 -17281
rect 4111 -17451 4121 -17391
rect 4181 -17451 4441 -17391
rect 4501 -17451 4511 -17391
rect 4111 -17461 4511 -17451
rect 4567 -17391 4967 -17281
rect 4567 -17451 4577 -17391
rect 4637 -17451 4897 -17391
rect 4957 -17451 4967 -17391
rect 4567 -17461 4967 -17451
rect 5023 -17391 5423 -17281
rect 5023 -17451 5033 -17391
rect 5093 -17451 5353 -17391
rect 5413 -17451 5423 -17391
rect 5023 -17461 5423 -17451
rect 5481 -17391 5881 -17281
rect 5481 -17451 5491 -17391
rect 5551 -17451 5811 -17391
rect 5871 -17451 5881 -17391
rect 5481 -17461 5881 -17451
rect 5937 -17391 6337 -17281
rect 5937 -17451 5947 -17391
rect 6007 -17451 6267 -17391
rect 6327 -17451 6337 -17391
rect 5937 -17461 6337 -17451
rect 6393 -17391 6793 -17281
rect 6393 -17451 6403 -17391
rect 6463 -17451 6723 -17391
rect 6783 -17451 6793 -17391
rect 6393 -17461 6793 -17451
rect 6851 -17391 7251 -17281
rect 6851 -17451 6861 -17391
rect 6921 -17451 7181 -17391
rect 7241 -17451 7251 -17391
rect 6851 -17461 7251 -17451
rect 7307 -17041 7707 -17031
rect 7307 -17101 7317 -17041
rect 7377 -17101 7637 -17041
rect 7697 -17101 7707 -17041
rect 7307 -17211 7707 -17101
rect 7763 -17041 8163 -17031
rect 7763 -17101 7773 -17041
rect 7833 -17101 8093 -17041
rect 8153 -17101 8163 -17041
rect 7763 -17211 8163 -17101
rect 8237 -17041 8637 -17031
rect 8237 -17101 8247 -17041
rect 8307 -17101 8567 -17041
rect 8627 -17101 8637 -17041
rect 8237 -17211 8637 -17101
rect 8693 -17041 9093 -17031
rect 8693 -17101 8703 -17041
rect 8763 -17101 9023 -17041
rect 9083 -17101 9093 -17041
rect 8693 -17211 9093 -17101
rect 9151 -17041 9551 -17031
rect 9151 -17101 9161 -17041
rect 9221 -17101 9481 -17041
rect 9541 -17101 9551 -17041
rect 9151 -17211 9551 -17101
rect 9607 -17041 10007 -17031
rect 9607 -17101 9617 -17041
rect 9677 -17101 9937 -17041
rect 9997 -17101 10007 -17041
rect 9607 -17211 10007 -17101
rect 10063 -17041 10463 -17031
rect 10063 -17101 10073 -17041
rect 10133 -17101 10393 -17041
rect 10453 -17101 10463 -17041
rect 10063 -17211 10463 -17101
rect 10521 -17041 10921 -17031
rect 10521 -17101 10531 -17041
rect 10591 -17101 10851 -17041
rect 10911 -17101 10921 -17041
rect 10521 -17211 10921 -17101
rect 7307 -17281 9093 -17211
rect 9150 -17281 10921 -17211
rect 7307 -17391 7707 -17281
rect 7307 -17451 7317 -17391
rect 7377 -17451 7637 -17391
rect 7697 -17451 7707 -17391
rect 7307 -17461 7707 -17451
rect 7763 -17391 8163 -17281
rect 7763 -17451 7773 -17391
rect 7833 -17451 8093 -17391
rect 8153 -17451 8163 -17391
rect 7763 -17461 8163 -17451
rect 8237 -17391 8637 -17281
rect 8237 -17451 8247 -17391
rect 8307 -17451 8567 -17391
rect 8627 -17451 8637 -17391
rect 8237 -17461 8637 -17451
rect 8693 -17391 9093 -17281
rect 8693 -17451 8703 -17391
rect 8763 -17451 9023 -17391
rect 9083 -17451 9093 -17391
rect 8693 -17461 9093 -17451
rect 9151 -17391 9551 -17281
rect 9151 -17451 9161 -17391
rect 9221 -17451 9481 -17391
rect 9541 -17451 9551 -17391
rect 9151 -17461 9551 -17451
rect 9607 -17391 10007 -17281
rect 9607 -17451 9617 -17391
rect 9677 -17451 9937 -17391
rect 9997 -17451 10007 -17391
rect 9607 -17461 10007 -17451
rect 10063 -17391 10463 -17281
rect 10063 -17451 10073 -17391
rect 10133 -17451 10393 -17391
rect 10453 -17451 10463 -17391
rect 10063 -17461 10463 -17451
rect 10521 -17391 10921 -17281
rect 10521 -17451 10531 -17391
rect 10591 -17451 10851 -17391
rect 10911 -17451 10921 -17391
rect 10521 -17461 10921 -17451
rect 10977 -17041 11377 -17031
rect 10977 -17101 10987 -17041
rect 11047 -17101 11307 -17041
rect 11367 -17101 11377 -17041
rect 10977 -17211 11377 -17101
rect 11433 -17041 11833 -17031
rect 11433 -17101 11443 -17041
rect 11503 -17101 11763 -17041
rect 11823 -17101 11833 -17041
rect 11433 -17211 11833 -17101
rect 11891 -17041 12291 -17031
rect 11891 -17101 11901 -17041
rect 11961 -17101 12221 -17041
rect 12281 -17101 12291 -17041
rect 11891 -17211 12291 -17101
rect 10977 -17281 12291 -17211
rect 10977 -17391 11377 -17281
rect 10977 -17451 10987 -17391
rect 11047 -17451 11307 -17391
rect 11367 -17451 11377 -17391
rect 10977 -17461 11377 -17451
rect 11433 -17391 11833 -17281
rect 11433 -17451 11443 -17391
rect 11503 -17451 11763 -17391
rect 11823 -17451 11833 -17391
rect 11433 -17461 11833 -17451
rect 11891 -17391 12291 -17281
rect 11891 -17451 11901 -17391
rect 11961 -17451 12221 -17391
rect 12281 -17451 12291 -17391
rect 11891 -17461 12291 -17451
rect 12347 -17041 12747 -17031
rect 12347 -17101 12357 -17041
rect 12417 -17101 12677 -17041
rect 12737 -17101 12747 -17041
rect 12347 -17211 12747 -17101
rect 12803 -17041 13203 -17031
rect 12803 -17101 12813 -17041
rect 12873 -17101 13133 -17041
rect 13193 -17101 13203 -17041
rect 12803 -17211 13203 -17101
rect 12347 -17281 13203 -17211
rect 12347 -17391 12747 -17281
rect 12347 -17451 12357 -17391
rect 12417 -17451 12677 -17391
rect 12737 -17451 12747 -17391
rect 12347 -17461 12747 -17451
rect 12803 -17391 13203 -17281
rect 12803 -17451 12813 -17391
rect 12873 -17451 13133 -17391
rect 13193 -17451 13203 -17391
rect 12803 -17461 13203 -17451
rect 13261 -17041 13661 -17031
rect 13261 -17101 13271 -17041
rect 13331 -17101 13591 -17041
rect 13651 -17101 13661 -17041
rect 13261 -17391 13661 -17101
rect 13261 -17451 13271 -17391
rect 13331 -17451 13591 -17391
rect 13651 -17451 13661 -17391
rect 13261 -17461 13661 -17451
rect 13717 -17041 14117 -17031
rect 13717 -17101 13727 -17041
rect 13787 -17101 14047 -17041
rect 14107 -17101 14117 -17041
rect 13717 -17391 14117 -17101
rect 13717 -17451 13727 -17391
rect 13787 -17451 14047 -17391
rect 14107 -17451 14117 -17391
rect 13717 -17461 14117 -17451
rect 14173 -17041 14573 -17031
rect 14173 -17101 14183 -17041
rect 14243 -17101 14503 -17041
rect 14563 -17101 14573 -17041
rect 14173 -17211 14573 -17101
rect 14631 -17041 15031 -17031
rect 14631 -17101 14641 -17041
rect 14701 -17101 14961 -17041
rect 15021 -17101 15031 -17041
rect 14631 -17211 15031 -17101
rect 15087 -17041 15487 -17031
rect 15087 -17101 15097 -17041
rect 15157 -17101 15417 -17041
rect 15477 -17101 15487 -17041
rect 15087 -17210 15487 -17101
rect 15087 -17211 15720 -17210
rect 14173 -17281 15720 -17211
rect 14173 -17391 14573 -17281
rect 14173 -17451 14183 -17391
rect 14243 -17451 14503 -17391
rect 14563 -17451 14573 -17391
rect 14173 -17461 14573 -17451
rect 14631 -17391 15031 -17281
rect 14631 -17451 14641 -17391
rect 14701 -17451 14961 -17391
rect 15021 -17451 15031 -17391
rect 14631 -17461 15031 -17451
rect 15087 -17391 15487 -17281
rect 15087 -17451 15097 -17391
rect 15157 -17451 15417 -17391
rect 15477 -17451 15487 -17391
rect 15087 -17461 15487 -17451
rect 66 -17523 80 -17461
rect 457 -17523 528 -17461
rect 913 -17523 984 -17461
rect 1371 -17523 1442 -17461
rect 1827 -17523 1898 -17461
rect 2283 -17523 2354 -17461
rect 2741 -17523 2811 -17461
rect 3197 -17523 3267 -17461
rect 3653 -17523 3723 -17461
rect 4111 -17523 4181 -17461
rect 4567 -17523 4637 -17461
rect 5023 -17523 5093 -17461
rect 5481 -17523 5551 -17461
rect 5937 -17523 6007 -17461
rect 6393 -17523 6463 -17461
rect 6851 -17523 6921 -17461
rect 7307 -17523 7377 -17461
rect 7763 -17523 7833 -17461
rect 8237 -17523 8307 -17461
rect 8693 -17523 8763 -17461
rect 9151 -17523 9221 -17461
rect 9607 -17523 9677 -17461
rect 10063 -17523 10133 -17461
rect 10521 -17523 10591 -17461
rect 10977 -17523 11047 -17461
rect 11433 -17523 11503 -17461
rect 11891 -17523 11961 -17461
rect 12347 -17523 12417 -17461
rect 12803 -17523 12873 -17461
rect 13261 -17523 13331 -17461
rect 14173 -17523 14243 -17461
rect 14631 -17523 14701 -17461
rect 66 -17533 400 -17523
rect 0 -17593 11 -17533
rect 71 -17593 331 -17533
rect 391 -17593 400 -17533
rect 0 -17883 14 -17593
rect 66 -17883 400 -17593
rect 0 -17943 11 -17883
rect 71 -17943 331 -17883
rect 391 -17943 400 -17883
rect 0 -18049 14 -17943
rect 66 -17953 400 -17943
rect 457 -17533 857 -17523
rect 457 -17593 467 -17533
rect 527 -17593 787 -17533
rect 847 -17593 857 -17533
rect 457 -17700 857 -17593
rect 913 -17533 1313 -17523
rect 913 -17593 923 -17533
rect 983 -17593 1243 -17533
rect 1303 -17593 1313 -17533
rect 913 -17700 1313 -17593
rect 1371 -17533 1771 -17523
rect 1371 -17593 1381 -17533
rect 1441 -17593 1701 -17533
rect 1761 -17593 1771 -17533
rect 1371 -17700 1771 -17593
rect 1827 -17533 2227 -17523
rect 1827 -17593 1837 -17533
rect 1897 -17593 2157 -17533
rect 2217 -17593 2227 -17533
rect 1827 -17700 2227 -17593
rect 2283 -17533 2683 -17523
rect 2283 -17593 2293 -17533
rect 2353 -17593 2613 -17533
rect 2673 -17593 2683 -17533
rect 2283 -17700 2683 -17593
rect 2741 -17533 3141 -17523
rect 2741 -17593 2751 -17533
rect 2811 -17593 3071 -17533
rect 3131 -17593 3141 -17533
rect 2741 -17700 3141 -17593
rect 3197 -17533 3597 -17523
rect 3197 -17593 3207 -17533
rect 3267 -17593 3527 -17533
rect 3587 -17593 3597 -17533
rect 3197 -17700 3597 -17593
rect 457 -17770 3597 -17700
rect 457 -17773 2683 -17770
rect 457 -17883 857 -17773
rect 457 -17943 467 -17883
rect 527 -17943 787 -17883
rect 847 -17943 857 -17883
rect 457 -17953 857 -17943
rect 913 -17883 1313 -17773
rect 913 -17943 923 -17883
rect 983 -17943 1243 -17883
rect 1303 -17943 1313 -17883
rect 913 -17953 1313 -17943
rect 1371 -17883 1771 -17773
rect 1371 -17943 1381 -17883
rect 1441 -17943 1701 -17883
rect 1761 -17943 1771 -17883
rect 1371 -17953 1771 -17943
rect 1827 -17883 2227 -17773
rect 1827 -17943 1837 -17883
rect 1897 -17943 2157 -17883
rect 2217 -17943 2227 -17883
rect 1827 -17953 2227 -17943
rect 2283 -17883 2683 -17773
rect 2283 -17943 2293 -17883
rect 2353 -17943 2613 -17883
rect 2673 -17943 2683 -17883
rect 2283 -17953 2683 -17943
rect 2741 -17773 3597 -17770
rect 2741 -17883 3141 -17773
rect 2741 -17943 2751 -17883
rect 2811 -17943 3071 -17883
rect 3131 -17943 3141 -17883
rect 2741 -17953 3141 -17943
rect 3197 -17883 3597 -17773
rect 3197 -17943 3207 -17883
rect 3267 -17943 3527 -17883
rect 3587 -17943 3597 -17883
rect 3197 -17953 3597 -17943
rect 3653 -17533 4053 -17523
rect 3653 -17593 3663 -17533
rect 3723 -17593 3983 -17533
rect 4043 -17593 4053 -17533
rect 3653 -17700 4053 -17593
rect 4111 -17533 4511 -17523
rect 4111 -17593 4121 -17533
rect 4181 -17593 4441 -17533
rect 4501 -17593 4511 -17533
rect 4111 -17700 4511 -17593
rect 4567 -17533 4967 -17523
rect 4567 -17593 4577 -17533
rect 4637 -17593 4897 -17533
rect 4957 -17593 4967 -17533
rect 4567 -17700 4967 -17593
rect 5023 -17533 5423 -17523
rect 5023 -17593 5033 -17533
rect 5093 -17593 5353 -17533
rect 5413 -17593 5423 -17533
rect 5023 -17700 5423 -17593
rect 5481 -17533 5881 -17523
rect 5481 -17593 5491 -17533
rect 5551 -17593 5811 -17533
rect 5871 -17593 5881 -17533
rect 5481 -17700 5881 -17593
rect 5937 -17533 6337 -17523
rect 5937 -17593 5947 -17533
rect 6007 -17593 6267 -17533
rect 6327 -17593 6337 -17533
rect 5937 -17700 6337 -17593
rect 6393 -17533 6793 -17523
rect 6393 -17593 6403 -17533
rect 6463 -17593 6723 -17533
rect 6783 -17593 6793 -17533
rect 6393 -17700 6793 -17593
rect 6851 -17533 7251 -17523
rect 6851 -17593 6861 -17533
rect 6921 -17593 7181 -17533
rect 7241 -17593 7251 -17533
rect 6851 -17700 7251 -17593
rect 3653 -17773 7251 -17700
rect 3653 -17883 4053 -17773
rect 3653 -17943 3663 -17883
rect 3723 -17943 3983 -17883
rect 4043 -17943 4053 -17883
rect 3653 -17953 4053 -17943
rect 4111 -17883 4511 -17773
rect 4111 -17943 4121 -17883
rect 4181 -17943 4441 -17883
rect 4501 -17943 4511 -17883
rect 4111 -17953 4511 -17943
rect 4567 -17883 4967 -17773
rect 4567 -17943 4577 -17883
rect 4637 -17943 4897 -17883
rect 4957 -17943 4967 -17883
rect 4567 -17953 4967 -17943
rect 5023 -17883 5423 -17773
rect 5023 -17943 5033 -17883
rect 5093 -17943 5353 -17883
rect 5413 -17943 5423 -17883
rect 5023 -17953 5423 -17943
rect 5481 -17883 5881 -17773
rect 5481 -17943 5491 -17883
rect 5551 -17943 5811 -17883
rect 5871 -17943 5881 -17883
rect 5481 -17953 5881 -17943
rect 5937 -17883 6337 -17773
rect 5937 -17943 5947 -17883
rect 6007 -17943 6267 -17883
rect 6327 -17943 6337 -17883
rect 5937 -17953 6337 -17943
rect 6393 -17883 6793 -17773
rect 6393 -17943 6403 -17883
rect 6463 -17943 6723 -17883
rect 6783 -17943 6793 -17883
rect 6393 -17953 6793 -17943
rect 6851 -17883 7251 -17773
rect 6851 -17943 6861 -17883
rect 6921 -17943 7181 -17883
rect 7241 -17943 7251 -17883
rect 6851 -17953 7251 -17943
rect 7307 -17533 7707 -17523
rect 7307 -17593 7317 -17533
rect 7377 -17593 7637 -17533
rect 7697 -17593 7707 -17533
rect 7307 -17700 7707 -17593
rect 7763 -17533 8163 -17523
rect 7763 -17593 7773 -17533
rect 7833 -17593 8093 -17533
rect 8153 -17593 8163 -17533
rect 7763 -17700 8163 -17593
rect 8237 -17533 8637 -17523
rect 8237 -17593 8247 -17533
rect 8307 -17593 8567 -17533
rect 8627 -17593 8637 -17533
rect 8237 -17700 8637 -17593
rect 8693 -17533 9093 -17523
rect 8693 -17593 8703 -17533
rect 8763 -17593 9023 -17533
rect 9083 -17593 9093 -17533
rect 8693 -17700 9093 -17593
rect 9151 -17533 9551 -17523
rect 9151 -17593 9161 -17533
rect 9221 -17593 9481 -17533
rect 9541 -17593 9551 -17533
rect 9151 -17700 9551 -17593
rect 9607 -17533 10007 -17523
rect 9607 -17593 9617 -17533
rect 9677 -17593 9937 -17533
rect 9997 -17593 10007 -17533
rect 9607 -17700 10007 -17593
rect 10063 -17533 10463 -17523
rect 10063 -17593 10073 -17533
rect 10133 -17593 10393 -17533
rect 10453 -17593 10463 -17533
rect 10063 -17700 10463 -17593
rect 10521 -17533 10921 -17523
rect 10521 -17593 10531 -17533
rect 10591 -17593 10851 -17533
rect 10911 -17593 10921 -17533
rect 10521 -17700 10921 -17593
rect 7307 -17773 9093 -17700
rect 9150 -17770 10921 -17700
rect 9150 -17773 10463 -17770
rect 7307 -17883 7707 -17773
rect 7307 -17943 7317 -17883
rect 7377 -17943 7637 -17883
rect 7697 -17943 7707 -17883
rect 7307 -17953 7707 -17943
rect 7763 -17883 8163 -17773
rect 7763 -17943 7773 -17883
rect 7833 -17943 8093 -17883
rect 8153 -17943 8163 -17883
rect 7763 -17953 8163 -17943
rect 8237 -17883 8637 -17773
rect 8237 -17943 8247 -17883
rect 8307 -17943 8567 -17883
rect 8627 -17943 8637 -17883
rect 8237 -17953 8637 -17943
rect 8693 -17883 9093 -17773
rect 8693 -17943 8703 -17883
rect 8763 -17943 9023 -17883
rect 9083 -17943 9093 -17883
rect 8693 -17953 9093 -17943
rect 9151 -17883 9551 -17773
rect 9151 -17943 9161 -17883
rect 9221 -17943 9481 -17883
rect 9541 -17943 9551 -17883
rect 9151 -17953 9551 -17943
rect 9607 -17883 10007 -17773
rect 9607 -17943 9617 -17883
rect 9677 -17943 9937 -17883
rect 9997 -17943 10007 -17883
rect 9607 -17953 10007 -17943
rect 10063 -17883 10463 -17773
rect 10063 -17943 10073 -17883
rect 10133 -17943 10393 -17883
rect 10453 -17943 10463 -17883
rect 10063 -17953 10463 -17943
rect 10521 -17883 10921 -17770
rect 10521 -17943 10531 -17883
rect 10591 -17943 10851 -17883
rect 10911 -17943 10921 -17883
rect 10521 -17953 10921 -17943
rect 10977 -17533 11377 -17523
rect 10977 -17593 10987 -17533
rect 11047 -17593 11307 -17533
rect 11367 -17593 11377 -17533
rect 10977 -17700 11377 -17593
rect 11433 -17533 11833 -17523
rect 11433 -17593 11443 -17533
rect 11503 -17593 11763 -17533
rect 11823 -17593 11833 -17533
rect 11433 -17700 11833 -17593
rect 11891 -17533 12291 -17523
rect 11891 -17593 11901 -17533
rect 11961 -17593 12221 -17533
rect 12281 -17593 12291 -17533
rect 11891 -17700 12291 -17593
rect 10977 -17773 12291 -17700
rect 10977 -17883 11377 -17773
rect 10977 -17943 10987 -17883
rect 11047 -17943 11307 -17883
rect 11367 -17943 11377 -17883
rect 10977 -17953 11377 -17943
rect 11433 -17883 11833 -17773
rect 11433 -17943 11443 -17883
rect 11503 -17943 11763 -17883
rect 11823 -17943 11833 -17883
rect 11433 -17953 11833 -17943
rect 11891 -17883 12291 -17773
rect 11891 -17943 11901 -17883
rect 11961 -17943 12221 -17883
rect 12281 -17943 12291 -17883
rect 11891 -17953 12291 -17943
rect 12347 -17533 12747 -17523
rect 12347 -17593 12357 -17533
rect 12417 -17593 12677 -17533
rect 12737 -17593 12747 -17533
rect 12347 -17700 12747 -17593
rect 12803 -17533 13203 -17523
rect 12803 -17593 12813 -17533
rect 12873 -17593 13133 -17533
rect 13193 -17593 13203 -17533
rect 12803 -17700 13203 -17593
rect 12347 -17773 13203 -17700
rect 12347 -17883 12747 -17773
rect 12347 -17943 12357 -17883
rect 12417 -17943 12677 -17883
rect 12737 -17943 12747 -17883
rect 12347 -17953 12747 -17943
rect 12803 -17883 13203 -17773
rect 12803 -17943 12813 -17883
rect 12873 -17943 13133 -17883
rect 13193 -17943 13203 -17883
rect 12803 -17953 13203 -17943
rect 13261 -17533 13661 -17523
rect 13261 -17593 13271 -17533
rect 13331 -17593 13591 -17533
rect 13651 -17593 13661 -17533
rect 13261 -17700 13661 -17593
rect 13717 -17533 14117 -17523
rect 13717 -17593 13727 -17533
rect 13787 -17593 14047 -17533
rect 14107 -17593 14117 -17533
rect 13717 -17700 14117 -17593
rect 14173 -17533 14573 -17523
rect 14173 -17593 14183 -17533
rect 14243 -17593 14503 -17533
rect 14563 -17593 14573 -17533
rect 14173 -17700 14573 -17593
rect 14631 -17533 15031 -17523
rect 14631 -17593 14641 -17533
rect 14701 -17593 14961 -17533
rect 15021 -17593 15031 -17533
rect 14631 -17700 15031 -17593
rect 15087 -17533 15487 -17523
rect 15087 -17593 15097 -17533
rect 15157 -17593 15417 -17533
rect 15477 -17593 15487 -17533
rect 15087 -17700 15487 -17593
rect 13261 -17773 15487 -17700
rect 13261 -17883 13661 -17773
rect 13261 -17943 13271 -17883
rect 13331 -17943 13591 -17883
rect 13651 -17943 13661 -17883
rect 13261 -17953 13661 -17943
rect 13717 -17883 14117 -17773
rect 13717 -17943 13727 -17883
rect 13787 -17943 14047 -17883
rect 14107 -17943 14117 -17883
rect 13717 -17953 14117 -17943
rect 14173 -17883 14573 -17773
rect 14173 -17943 14183 -17883
rect 14243 -17943 14503 -17883
rect 14563 -17943 14573 -17883
rect 14173 -17953 14573 -17943
rect 14631 -17883 15031 -17773
rect 14631 -17943 14641 -17883
rect 14701 -17943 14961 -17883
rect 15021 -17943 15031 -17883
rect 14631 -17953 15031 -17943
rect 15087 -17883 15487 -17773
rect 15087 -17943 15097 -17883
rect 15157 -17943 15417 -17883
rect 15477 -17943 15487 -17883
rect 15087 -17953 15487 -17943
rect 66 -18039 80 -17953
rect 457 -18039 527 -17953
rect 913 -18039 983 -17953
rect 1371 -18039 1441 -17953
rect 1827 -18039 1897 -17953
rect 2283 -18039 2353 -17953
rect 2741 -18039 2811 -17953
rect 3197 -18039 3267 -17953
rect 3653 -18039 3723 -17953
rect 4111 -18039 4181 -17953
rect 4567 -18039 4637 -17953
rect 5023 -18039 5093 -17953
rect 5481 -18039 5551 -17953
rect 5937 -18039 6007 -17953
rect 6393 -18039 6463 -17953
rect 6851 -18039 6921 -17953
rect 7307 -18039 7377 -17953
rect 7763 -18039 7833 -17953
rect 8237 -18039 8307 -17953
rect 8693 -18039 8763 -17953
rect 9151 -18039 9221 -17953
rect 9607 -18039 9677 -17953
rect 10063 -18039 10133 -17953
rect 10521 -18039 10591 -17953
rect 10977 -18039 11047 -17953
rect 11433 -18039 11503 -17953
rect 11891 -18039 11961 -17953
rect 12347 -18039 12417 -17953
rect 12803 -18039 12873 -17953
rect 66 -18049 400 -18039
rect 0 -18109 11 -18049
rect 71 -18109 331 -18049
rect 391 -18109 400 -18049
rect 0 -18399 14 -18109
rect 66 -18399 400 -18109
rect 0 -18459 11 -18399
rect 71 -18459 331 -18399
rect 391 -18459 400 -18399
rect 0 -18551 14 -18459
rect 66 -18469 400 -18459
rect 457 -18049 857 -18039
rect 457 -18109 467 -18049
rect 527 -18109 787 -18049
rect 847 -18109 857 -18049
rect 457 -18219 857 -18109
rect 913 -18049 1313 -18039
rect 913 -18109 923 -18049
rect 983 -18109 1243 -18049
rect 1303 -18109 1313 -18049
rect 913 -18219 1313 -18109
rect 1371 -18049 1771 -18039
rect 1371 -18109 1381 -18049
rect 1441 -18109 1701 -18049
rect 1761 -18109 1771 -18049
rect 1371 -18219 1771 -18109
rect 1827 -18049 2227 -18039
rect 1827 -18109 1837 -18049
rect 1897 -18109 2157 -18049
rect 2217 -18109 2227 -18049
rect 1827 -18219 2227 -18109
rect 2283 -18049 2683 -18039
rect 2283 -18109 2293 -18049
rect 2353 -18109 2613 -18049
rect 2673 -18109 2683 -18049
rect 2283 -18219 2683 -18109
rect 457 -18220 2683 -18219
rect 2741 -18049 3141 -18039
rect 2741 -18109 2751 -18049
rect 2811 -18109 3071 -18049
rect 3131 -18109 3141 -18049
rect 2741 -18219 3141 -18109
rect 3197 -18049 3597 -18039
rect 3197 -18109 3207 -18049
rect 3267 -18109 3527 -18049
rect 3587 -18109 3597 -18049
rect 3197 -18219 3597 -18109
rect 2741 -18220 3597 -18219
rect 457 -18290 3597 -18220
rect 457 -18399 857 -18290
rect 457 -18459 467 -18399
rect 527 -18459 787 -18399
rect 847 -18459 857 -18399
rect 457 -18469 857 -18459
rect 913 -18399 1313 -18290
rect 913 -18459 923 -18399
rect 983 -18459 1243 -18399
rect 1303 -18459 1313 -18399
rect 913 -18469 1313 -18459
rect 1371 -18399 1771 -18290
rect 1371 -18459 1381 -18399
rect 1441 -18459 1701 -18399
rect 1761 -18459 1771 -18399
rect 1371 -18469 1771 -18459
rect 1827 -18399 2227 -18290
rect 1827 -18459 1837 -18399
rect 1897 -18459 2157 -18399
rect 2217 -18459 2227 -18399
rect 1827 -18469 2227 -18459
rect 2283 -18399 2683 -18290
rect 2283 -18459 2293 -18399
rect 2353 -18459 2613 -18399
rect 2673 -18459 2683 -18399
rect 2283 -18469 2683 -18459
rect 2741 -18399 3141 -18290
rect 2741 -18459 2751 -18399
rect 2811 -18459 3071 -18399
rect 3131 -18459 3141 -18399
rect 2741 -18469 3141 -18459
rect 3197 -18399 3597 -18290
rect 3197 -18459 3207 -18399
rect 3267 -18459 3527 -18399
rect 3587 -18459 3597 -18399
rect 3197 -18469 3597 -18459
rect 3653 -18049 4053 -18039
rect 3653 -18109 3663 -18049
rect 3723 -18109 3983 -18049
rect 4043 -18109 4053 -18049
rect 3653 -18219 4053 -18109
rect 4111 -18049 4511 -18039
rect 4111 -18109 4121 -18049
rect 4181 -18109 4441 -18049
rect 4501 -18109 4511 -18049
rect 4111 -18219 4511 -18109
rect 4567 -18049 4967 -18039
rect 4567 -18109 4577 -18049
rect 4637 -18109 4897 -18049
rect 4957 -18109 4967 -18049
rect 4567 -18219 4967 -18109
rect 5023 -18049 5423 -18039
rect 5023 -18109 5033 -18049
rect 5093 -18109 5353 -18049
rect 5413 -18109 5423 -18049
rect 5023 -18219 5423 -18109
rect 5481 -18049 5881 -18039
rect 5481 -18109 5491 -18049
rect 5551 -18109 5811 -18049
rect 5871 -18109 5881 -18049
rect 5481 -18219 5881 -18109
rect 5937 -18049 6337 -18039
rect 5937 -18109 5947 -18049
rect 6007 -18109 6267 -18049
rect 6327 -18109 6337 -18049
rect 5937 -18219 6337 -18109
rect 6393 -18049 6793 -18039
rect 6393 -18109 6403 -18049
rect 6463 -18109 6723 -18049
rect 6783 -18109 6793 -18049
rect 6393 -18219 6793 -18109
rect 6851 -18049 7251 -18039
rect 6851 -18109 6861 -18049
rect 6921 -18109 7181 -18049
rect 7241 -18109 7251 -18049
rect 6851 -18219 7251 -18109
rect 3653 -18290 7251 -18219
rect 3653 -18399 4053 -18290
rect 3653 -18459 3663 -18399
rect 3723 -18459 3983 -18399
rect 4043 -18459 4053 -18399
rect 3653 -18469 4053 -18459
rect 4111 -18399 4511 -18290
rect 4111 -18459 4121 -18399
rect 4181 -18459 4441 -18399
rect 4501 -18459 4511 -18399
rect 4111 -18469 4511 -18459
rect 4567 -18399 4967 -18290
rect 4567 -18459 4577 -18399
rect 4637 -18459 4897 -18399
rect 4957 -18459 4967 -18399
rect 4567 -18469 4967 -18459
rect 5023 -18399 5423 -18290
rect 5023 -18459 5033 -18399
rect 5093 -18459 5353 -18399
rect 5413 -18459 5423 -18399
rect 5023 -18469 5423 -18459
rect 5481 -18399 5881 -18290
rect 5481 -18459 5491 -18399
rect 5551 -18459 5811 -18399
rect 5871 -18459 5881 -18399
rect 5481 -18469 5881 -18459
rect 5937 -18399 6337 -18290
rect 5937 -18459 5947 -18399
rect 6007 -18459 6267 -18399
rect 6327 -18459 6337 -18399
rect 5937 -18469 6337 -18459
rect 6393 -18399 6793 -18290
rect 6393 -18459 6403 -18399
rect 6463 -18459 6723 -18399
rect 6783 -18459 6793 -18399
rect 6393 -18469 6793 -18459
rect 6851 -18399 7251 -18290
rect 6851 -18459 6861 -18399
rect 6921 -18459 7181 -18399
rect 7241 -18459 7251 -18399
rect 6851 -18469 7251 -18459
rect 7307 -18049 7707 -18039
rect 7307 -18109 7317 -18049
rect 7377 -18109 7637 -18049
rect 7697 -18109 7707 -18049
rect 7307 -18219 7707 -18109
rect 7763 -18049 8163 -18039
rect 7763 -18109 7773 -18049
rect 7833 -18109 8093 -18049
rect 8153 -18109 8163 -18049
rect 7763 -18219 8163 -18109
rect 8237 -18049 8637 -18039
rect 8237 -18109 8247 -18049
rect 8307 -18109 8567 -18049
rect 8627 -18109 8637 -18049
rect 8237 -18219 8637 -18109
rect 8693 -18049 9093 -18039
rect 8693 -18109 8703 -18049
rect 8763 -18109 9023 -18049
rect 9083 -18109 9093 -18049
rect 8693 -18219 9093 -18109
rect 9151 -18049 9551 -18039
rect 9151 -18109 9161 -18049
rect 9221 -18109 9481 -18049
rect 9541 -18109 9551 -18049
rect 9151 -18219 9551 -18109
rect 9607 -18049 10007 -18039
rect 9607 -18109 9617 -18049
rect 9677 -18109 9937 -18049
rect 9997 -18109 10007 -18049
rect 9607 -18219 10007 -18109
rect 10063 -18049 10463 -18039
rect 10063 -18109 10073 -18049
rect 10133 -18109 10393 -18049
rect 10453 -18109 10463 -18049
rect 10063 -18219 10463 -18109
rect 7307 -18290 9093 -18219
rect 9150 -18220 10463 -18219
rect 10521 -18049 10921 -18039
rect 10521 -18109 10531 -18049
rect 10591 -18109 10851 -18049
rect 10911 -18109 10921 -18049
rect 10521 -18220 10921 -18109
rect 9150 -18290 10921 -18220
rect 7307 -18399 7707 -18290
rect 7307 -18459 7317 -18399
rect 7377 -18459 7637 -18399
rect 7697 -18459 7707 -18399
rect 7307 -18469 7707 -18459
rect 7763 -18399 8163 -18290
rect 7763 -18459 7773 -18399
rect 7833 -18459 8093 -18399
rect 8153 -18459 8163 -18399
rect 7763 -18469 8163 -18459
rect 8237 -18399 8637 -18290
rect 8237 -18459 8247 -18399
rect 8307 -18459 8567 -18399
rect 8627 -18459 8637 -18399
rect 8237 -18469 8637 -18459
rect 8693 -18399 9093 -18290
rect 8693 -18459 8703 -18399
rect 8763 -18459 9023 -18399
rect 9083 -18459 9093 -18399
rect 8693 -18469 9093 -18459
rect 9151 -18399 9551 -18290
rect 9151 -18459 9161 -18399
rect 9221 -18459 9481 -18399
rect 9541 -18459 9551 -18399
rect 9151 -18469 9551 -18459
rect 9607 -18399 10007 -18290
rect 9607 -18459 9617 -18399
rect 9677 -18459 9937 -18399
rect 9997 -18459 10007 -18399
rect 9607 -18469 10007 -18459
rect 10063 -18399 10463 -18290
rect 10063 -18459 10073 -18399
rect 10133 -18459 10393 -18399
rect 10453 -18459 10463 -18399
rect 10063 -18469 10463 -18459
rect 10521 -18399 10921 -18290
rect 10521 -18459 10531 -18399
rect 10591 -18459 10851 -18399
rect 10911 -18459 10921 -18399
rect 10521 -18469 10921 -18459
rect 10977 -18049 11377 -18039
rect 10977 -18109 10987 -18049
rect 11047 -18109 11307 -18049
rect 11367 -18109 11377 -18049
rect 10977 -18219 11377 -18109
rect 11433 -18049 11833 -18039
rect 11433 -18109 11443 -18049
rect 11503 -18109 11763 -18049
rect 11823 -18109 11833 -18049
rect 11433 -18219 11833 -18109
rect 11891 -18049 12291 -18039
rect 11891 -18109 11901 -18049
rect 11961 -18109 12221 -18049
rect 12281 -18109 12291 -18049
rect 11891 -18219 12291 -18109
rect 10977 -18290 12291 -18219
rect 10977 -18399 11377 -18290
rect 10977 -18459 10987 -18399
rect 11047 -18459 11307 -18399
rect 11367 -18459 11377 -18399
rect 10977 -18469 11377 -18459
rect 11433 -18399 11833 -18290
rect 11433 -18459 11443 -18399
rect 11503 -18459 11763 -18399
rect 11823 -18459 11833 -18399
rect 11433 -18469 11833 -18459
rect 11891 -18399 12291 -18290
rect 11891 -18459 11901 -18399
rect 11961 -18459 12221 -18399
rect 12281 -18459 12291 -18399
rect 11891 -18469 12291 -18459
rect 12347 -18049 12747 -18039
rect 12347 -18109 12357 -18049
rect 12417 -18109 12677 -18049
rect 12737 -18109 12747 -18049
rect 12347 -18219 12747 -18109
rect 12803 -18049 13203 -18039
rect 12803 -18109 12813 -18049
rect 12873 -18109 13133 -18049
rect 13193 -18109 13203 -18049
rect 12803 -18219 13203 -18109
rect 13261 -18049 13661 -18039
rect 13261 -18109 13271 -18049
rect 13331 -18109 13591 -18049
rect 13651 -18109 13661 -18049
rect 13261 -18219 13661 -18109
rect 13717 -18049 14117 -18039
rect 13717 -18109 13727 -18049
rect 13787 -18109 14047 -18049
rect 14107 -18109 14117 -18049
rect 13717 -18219 14117 -18109
rect 14173 -18049 14573 -18039
rect 14173 -18109 14183 -18049
rect 14243 -18109 14503 -18049
rect 14563 -18109 14573 -18049
rect 14173 -18219 14573 -18109
rect 14631 -18049 15031 -18039
rect 14631 -18109 14641 -18049
rect 14701 -18109 14961 -18049
rect 15021 -18109 15031 -18049
rect 14631 -18219 15031 -18109
rect 15087 -18049 15487 -18039
rect 15087 -18109 15097 -18049
rect 15157 -18109 15417 -18049
rect 15477 -18109 15487 -18049
rect 15087 -18219 15487 -18109
rect 12347 -18290 15720 -18219
rect 12347 -18399 12747 -18290
rect 12347 -18459 12357 -18399
rect 12417 -18459 12677 -18399
rect 12737 -18459 12747 -18399
rect 12347 -18469 12747 -18459
rect 12803 -18399 13203 -18290
rect 12803 -18459 12813 -18399
rect 12873 -18459 13133 -18399
rect 13193 -18459 13203 -18399
rect 12803 -18469 13203 -18459
rect 13261 -18399 13661 -18290
rect 13261 -18459 13271 -18399
rect 13331 -18459 13591 -18399
rect 13651 -18459 13661 -18399
rect 13261 -18469 13661 -18459
rect 13717 -18399 14117 -18290
rect 13717 -18459 13727 -18399
rect 13787 -18459 14047 -18399
rect 14107 -18459 14117 -18399
rect 13717 -18469 14117 -18459
rect 14173 -18399 14573 -18290
rect 14173 -18459 14183 -18399
rect 14243 -18459 14503 -18399
rect 14563 -18459 14573 -18399
rect 14173 -18469 14573 -18459
rect 14631 -18399 15031 -18290
rect 14631 -18459 14641 -18399
rect 14701 -18459 14961 -18399
rect 15021 -18459 15031 -18399
rect 14631 -18469 15031 -18459
rect 15087 -18399 15487 -18290
rect 15087 -18459 15097 -18399
rect 15157 -18459 15417 -18399
rect 15477 -18459 15487 -18399
rect 15087 -18469 15487 -18459
rect 66 -18541 80 -18469
rect 457 -18541 527 -18469
rect 913 -18541 984 -18469
rect 1371 -18541 1442 -18469
rect 1827 -18541 1898 -18469
rect 2283 -18541 2354 -18469
rect 2741 -18541 2812 -18469
rect 3197 -18541 3268 -18469
rect 3653 -18541 3724 -18469
rect 4111 -18541 4182 -18469
rect 4567 -18541 4638 -18469
rect 5023 -18541 5094 -18469
rect 5481 -18541 5552 -18469
rect 5937 -18541 6008 -18469
rect 6393 -18541 6464 -18469
rect 6851 -18541 6922 -18469
rect 7307 -18541 7378 -18469
rect 7763 -18541 7834 -18469
rect 8237 -18541 8308 -18469
rect 8693 -18541 8764 -18469
rect 9151 -18541 9222 -18469
rect 9607 -18541 9678 -18469
rect 10063 -18541 10134 -18469
rect 10521 -18541 10592 -18469
rect 10977 -18541 11048 -18469
rect 11433 -18541 11504 -18469
rect 11891 -18541 11962 -18469
rect 13717 -18470 13788 -18469
rect 14173 -18470 14244 -18469
rect 13261 -18541 13332 -18540
rect 14631 -18541 14702 -18540
rect 66 -18551 400 -18541
rect 0 -18611 11 -18551
rect 71 -18611 331 -18551
rect 391 -18611 400 -18551
rect 0 -18901 14 -18611
rect 66 -18901 400 -18611
rect 0 -18961 11 -18901
rect 71 -18961 331 -18901
rect 391 -18961 400 -18901
rect 0 -19043 14 -18961
rect 66 -18971 400 -18961
rect 457 -18551 857 -18541
rect 457 -18611 467 -18551
rect 527 -18611 787 -18551
rect 847 -18611 857 -18551
rect 457 -18721 857 -18611
rect 913 -18551 1313 -18541
rect 913 -18611 923 -18551
rect 983 -18611 1243 -18551
rect 1303 -18611 1313 -18551
rect 913 -18721 1313 -18611
rect 1371 -18551 1771 -18541
rect 1371 -18611 1381 -18551
rect 1441 -18611 1701 -18551
rect 1761 -18611 1771 -18551
rect 1371 -18721 1771 -18611
rect 1827 -18551 2227 -18541
rect 1827 -18611 1837 -18551
rect 1897 -18611 2157 -18551
rect 2217 -18611 2227 -18551
rect 1827 -18721 2227 -18611
rect 2283 -18551 2683 -18541
rect 2283 -18611 2293 -18551
rect 2353 -18611 2613 -18551
rect 2673 -18611 2683 -18551
rect 2283 -18721 2683 -18611
rect 2741 -18551 3141 -18541
rect 2741 -18611 2751 -18551
rect 2811 -18611 3071 -18551
rect 3131 -18611 3141 -18551
rect 2741 -18721 3141 -18611
rect 3197 -18551 3597 -18541
rect 3197 -18611 3207 -18551
rect 3267 -18611 3527 -18551
rect 3587 -18611 3597 -18551
rect 3197 -18721 3597 -18611
rect 457 -18791 3597 -18721
rect 457 -18901 857 -18791
rect 457 -18961 467 -18901
rect 527 -18961 787 -18901
rect 847 -18961 857 -18901
rect 457 -18971 857 -18961
rect 913 -18901 1313 -18791
rect 913 -18961 923 -18901
rect 983 -18961 1243 -18901
rect 1303 -18961 1313 -18901
rect 913 -18971 1313 -18961
rect 1371 -18901 1771 -18791
rect 1371 -18961 1381 -18901
rect 1441 -18961 1701 -18901
rect 1761 -18961 1771 -18901
rect 1371 -18971 1771 -18961
rect 1827 -18901 2227 -18791
rect 1827 -18961 1837 -18901
rect 1897 -18961 2157 -18901
rect 2217 -18961 2227 -18901
rect 1827 -18971 2227 -18961
rect 2283 -18901 2683 -18791
rect 2283 -18961 2293 -18901
rect 2353 -18961 2613 -18901
rect 2673 -18961 2683 -18901
rect 2283 -18971 2683 -18961
rect 2741 -18901 3141 -18791
rect 2741 -18961 2751 -18901
rect 2811 -18961 3071 -18901
rect 3131 -18961 3141 -18901
rect 2741 -18971 3141 -18961
rect 3197 -18901 3597 -18791
rect 3197 -18961 3207 -18901
rect 3267 -18961 3527 -18901
rect 3587 -18961 3597 -18901
rect 3197 -18971 3597 -18961
rect 3653 -18551 4053 -18541
rect 3653 -18611 3663 -18551
rect 3723 -18611 3983 -18551
rect 4043 -18611 4053 -18551
rect 3653 -18721 4053 -18611
rect 4111 -18551 4511 -18541
rect 4111 -18611 4121 -18551
rect 4181 -18611 4441 -18551
rect 4501 -18611 4511 -18551
rect 4111 -18721 4511 -18611
rect 4567 -18551 4967 -18541
rect 4567 -18611 4577 -18551
rect 4637 -18611 4897 -18551
rect 4957 -18611 4967 -18551
rect 4567 -18721 4967 -18611
rect 5023 -18551 5423 -18541
rect 5023 -18611 5033 -18551
rect 5093 -18611 5353 -18551
rect 5413 -18611 5423 -18551
rect 5023 -18721 5423 -18611
rect 5481 -18551 5881 -18541
rect 5481 -18611 5491 -18551
rect 5551 -18611 5811 -18551
rect 5871 -18611 5881 -18551
rect 5481 -18721 5881 -18611
rect 5937 -18551 6337 -18541
rect 5937 -18611 5947 -18551
rect 6007 -18611 6267 -18551
rect 6327 -18611 6337 -18551
rect 5937 -18721 6337 -18611
rect 6393 -18551 6793 -18541
rect 6393 -18611 6403 -18551
rect 6463 -18611 6723 -18551
rect 6783 -18611 6793 -18551
rect 6393 -18721 6793 -18611
rect 6851 -18551 7251 -18541
rect 6851 -18611 6861 -18551
rect 6921 -18611 7181 -18551
rect 7241 -18611 7251 -18551
rect 6851 -18721 7251 -18611
rect 3653 -18791 7251 -18721
rect 3653 -18901 4053 -18791
rect 3653 -18961 3663 -18901
rect 3723 -18961 3983 -18901
rect 4043 -18961 4053 -18901
rect 3653 -18971 4053 -18961
rect 4111 -18901 4511 -18791
rect 4111 -18961 4121 -18901
rect 4181 -18961 4441 -18901
rect 4501 -18961 4511 -18901
rect 4111 -18971 4511 -18961
rect 4567 -18901 4967 -18791
rect 4567 -18961 4577 -18901
rect 4637 -18961 4897 -18901
rect 4957 -18961 4967 -18901
rect 4567 -18971 4967 -18961
rect 5023 -18901 5423 -18791
rect 5023 -18961 5033 -18901
rect 5093 -18961 5353 -18901
rect 5413 -18961 5423 -18901
rect 5023 -18971 5423 -18961
rect 5481 -18901 5881 -18791
rect 5481 -18961 5491 -18901
rect 5551 -18961 5811 -18901
rect 5871 -18961 5881 -18901
rect 5481 -18971 5881 -18961
rect 5937 -18901 6337 -18791
rect 5937 -18961 5947 -18901
rect 6007 -18961 6267 -18901
rect 6327 -18961 6337 -18901
rect 5937 -18971 6337 -18961
rect 6393 -18901 6793 -18791
rect 6393 -18961 6403 -18901
rect 6463 -18961 6723 -18901
rect 6783 -18961 6793 -18901
rect 6393 -18971 6793 -18961
rect 6851 -18901 7251 -18791
rect 6851 -18961 6861 -18901
rect 6921 -18961 7181 -18901
rect 7241 -18961 7251 -18901
rect 6851 -18971 7251 -18961
rect 7307 -18551 7707 -18541
rect 7307 -18611 7317 -18551
rect 7377 -18611 7637 -18551
rect 7697 -18611 7707 -18551
rect 7307 -18721 7707 -18611
rect 7763 -18551 8163 -18541
rect 7763 -18611 7773 -18551
rect 7833 -18611 8093 -18551
rect 8153 -18611 8163 -18551
rect 7763 -18721 8163 -18611
rect 8237 -18551 8637 -18541
rect 8237 -18611 8247 -18551
rect 8307 -18611 8567 -18551
rect 8627 -18611 8637 -18551
rect 8237 -18721 8637 -18611
rect 8693 -18551 9093 -18541
rect 8693 -18611 8703 -18551
rect 8763 -18611 9023 -18551
rect 9083 -18611 9093 -18551
rect 8693 -18721 9093 -18611
rect 9151 -18551 9551 -18541
rect 9151 -18611 9161 -18551
rect 9221 -18611 9481 -18551
rect 9541 -18611 9551 -18551
rect 9151 -18721 9551 -18611
rect 9607 -18551 10007 -18541
rect 9607 -18611 9617 -18551
rect 9677 -18611 9937 -18551
rect 9997 -18611 10007 -18551
rect 9607 -18721 10007 -18611
rect 10063 -18551 10463 -18541
rect 10063 -18611 10073 -18551
rect 10133 -18611 10393 -18551
rect 10453 -18611 10463 -18551
rect 10063 -18721 10463 -18611
rect 10521 -18551 10921 -18541
rect 10521 -18611 10531 -18551
rect 10591 -18611 10851 -18551
rect 10911 -18611 10921 -18551
rect 10521 -18721 10921 -18611
rect 7307 -18791 9093 -18721
rect 9150 -18791 10921 -18721
rect 7307 -18901 7707 -18791
rect 7307 -18961 7317 -18901
rect 7377 -18961 7637 -18901
rect 7697 -18961 7707 -18901
rect 7307 -18971 7707 -18961
rect 7763 -18901 8163 -18791
rect 7763 -18961 7773 -18901
rect 7833 -18961 8093 -18901
rect 8153 -18961 8163 -18901
rect 7763 -18971 8163 -18961
rect 8237 -18901 8637 -18791
rect 8237 -18961 8247 -18901
rect 8307 -18961 8567 -18901
rect 8627 -18961 8637 -18901
rect 8237 -18971 8637 -18961
rect 8693 -18901 9093 -18791
rect 8693 -18961 8703 -18901
rect 8763 -18961 9023 -18901
rect 9083 -18961 9093 -18901
rect 8693 -18971 9093 -18961
rect 9151 -18901 9551 -18791
rect 9151 -18961 9161 -18901
rect 9221 -18961 9481 -18901
rect 9541 -18961 9551 -18901
rect 9151 -18971 9551 -18961
rect 9607 -18901 10007 -18791
rect 9607 -18961 9617 -18901
rect 9677 -18961 9937 -18901
rect 9997 -18961 10007 -18901
rect 9607 -18971 10007 -18961
rect 10063 -18901 10463 -18791
rect 10063 -18961 10073 -18901
rect 10133 -18961 10393 -18901
rect 10453 -18961 10463 -18901
rect 10063 -18971 10463 -18961
rect 10521 -18901 10921 -18791
rect 10521 -18961 10531 -18901
rect 10591 -18961 10851 -18901
rect 10911 -18961 10921 -18901
rect 10521 -18971 10921 -18961
rect 10977 -18551 11377 -18541
rect 10977 -18611 10987 -18551
rect 11047 -18611 11307 -18551
rect 11367 -18611 11377 -18551
rect 10977 -18721 11377 -18611
rect 11433 -18551 11833 -18541
rect 11433 -18611 11443 -18551
rect 11503 -18611 11763 -18551
rect 11823 -18611 11833 -18551
rect 11433 -18721 11833 -18611
rect 11891 -18551 12291 -18541
rect 11891 -18611 11901 -18551
rect 11961 -18611 12221 -18551
rect 12281 -18611 12291 -18551
rect 11891 -18721 12291 -18611
rect 12347 -18551 12747 -18541
rect 12347 -18611 12357 -18551
rect 12417 -18611 12677 -18551
rect 12737 -18611 12747 -18551
rect 12347 -18721 12747 -18611
rect 12803 -18551 13203 -18541
rect 12803 -18611 12813 -18551
rect 12873 -18611 13133 -18551
rect 13193 -18611 13203 -18551
rect 12803 -18721 13203 -18611
rect 13261 -18551 13661 -18541
rect 13261 -18611 13271 -18551
rect 13331 -18611 13591 -18551
rect 13651 -18611 13661 -18551
rect 13261 -18721 13661 -18611
rect 13717 -18551 14117 -18541
rect 13717 -18611 13727 -18551
rect 13787 -18611 14047 -18551
rect 14107 -18611 14117 -18551
rect 13717 -18721 14117 -18611
rect 14173 -18551 14573 -18541
rect 14173 -18611 14183 -18551
rect 14243 -18611 14503 -18551
rect 14563 -18611 14573 -18551
rect 14173 -18721 14573 -18611
rect 14631 -18551 15031 -18541
rect 14631 -18611 14641 -18551
rect 14701 -18611 14961 -18551
rect 15021 -18611 15031 -18551
rect 14631 -18721 15031 -18611
rect 15087 -18551 15487 -18541
rect 15087 -18611 15097 -18551
rect 15157 -18611 15417 -18551
rect 15477 -18611 15487 -18551
rect 15087 -18720 15487 -18611
rect 15087 -18721 15721 -18720
rect 10977 -18791 15721 -18721
rect 10977 -18901 11377 -18791
rect 10977 -18961 10987 -18901
rect 11047 -18961 11307 -18901
rect 11367 -18961 11377 -18901
rect 10977 -18971 11377 -18961
rect 11433 -18901 11833 -18791
rect 11433 -18961 11443 -18901
rect 11503 -18961 11763 -18901
rect 11823 -18961 11833 -18901
rect 11433 -18971 11833 -18961
rect 11891 -18901 12291 -18791
rect 11891 -18961 11901 -18901
rect 11961 -18961 12221 -18901
rect 12281 -18961 12291 -18901
rect 11891 -18971 12291 -18961
rect 12347 -18901 12747 -18791
rect 12347 -18961 12357 -18901
rect 12417 -18961 12677 -18901
rect 12737 -18961 12747 -18901
rect 12347 -18971 12747 -18961
rect 12803 -18901 13203 -18791
rect 12803 -18961 12813 -18901
rect 12873 -18961 13133 -18901
rect 13193 -18961 13203 -18901
rect 12803 -18971 13203 -18961
rect 13261 -18901 13661 -18791
rect 13261 -18961 13271 -18901
rect 13331 -18961 13591 -18901
rect 13651 -18961 13661 -18901
rect 13261 -18971 13661 -18961
rect 13717 -18901 14117 -18791
rect 13717 -18961 13727 -18901
rect 13787 -18961 14047 -18901
rect 14107 -18961 14117 -18901
rect 13717 -18971 14117 -18961
rect 14173 -18901 14573 -18791
rect 14173 -18961 14183 -18901
rect 14243 -18961 14503 -18901
rect 14563 -18961 14573 -18901
rect 14173 -18971 14573 -18961
rect 14631 -18901 15031 -18791
rect 14631 -18961 14641 -18901
rect 14701 -18961 14961 -18901
rect 15021 -18961 15031 -18901
rect 14631 -18971 15031 -18961
rect 15087 -18901 15487 -18791
rect 15087 -18961 15097 -18901
rect 15157 -18961 15417 -18901
rect 15477 -18961 15487 -18901
rect 15087 -18971 15487 -18961
rect 66 -19033 80 -18971
rect 457 -19033 528 -18971
rect 913 -19033 984 -18971
rect 1371 -19033 1442 -18971
rect 1827 -19033 1898 -18971
rect 2283 -19033 2354 -18971
rect 2741 -19033 2811 -18971
rect 3197 -19033 3267 -18971
rect 3653 -19033 3723 -18971
rect 4111 -19033 4181 -18971
rect 4567 -19033 4637 -18971
rect 5023 -19033 5093 -18971
rect 5481 -19033 5551 -18971
rect 5937 -19033 6007 -18971
rect 6393 -19033 6463 -18971
rect 6851 -19033 6921 -18971
rect 7307 -19033 7377 -18971
rect 7763 -19033 7833 -18971
rect 8237 -19033 8307 -18971
rect 8693 -19033 8763 -18971
rect 9151 -19033 9221 -18971
rect 9607 -19033 9677 -18971
rect 10063 -19033 10133 -18971
rect 10521 -19033 10591 -18971
rect 10977 -19033 11047 -18971
rect 11433 -19033 11503 -18971
rect 11891 -19033 11961 -18971
rect 12347 -19033 12417 -18971
rect 12803 -19033 12873 -18971
rect 13261 -19033 13331 -18971
rect 13717 -19033 13787 -18971
rect 14173 -19033 14243 -18971
rect 14631 -19033 14701 -18971
rect 66 -19043 400 -19033
rect 0 -19103 11 -19043
rect 71 -19103 331 -19043
rect 391 -19103 400 -19043
rect 0 -19393 14 -19103
rect 66 -19393 400 -19103
rect 0 -19453 11 -19393
rect 71 -19453 331 -19393
rect 391 -19453 400 -19393
rect 0 -19537 14 -19453
rect 66 -19463 400 -19453
rect 457 -19043 857 -19033
rect 457 -19103 467 -19043
rect 527 -19103 787 -19043
rect 847 -19103 857 -19043
rect 457 -19211 857 -19103
rect 913 -19043 1313 -19033
rect 913 -19103 923 -19043
rect 983 -19103 1243 -19043
rect 1303 -19103 1313 -19043
rect 913 -19211 1313 -19103
rect 1371 -19043 1771 -19033
rect 1371 -19103 1381 -19043
rect 1441 -19103 1701 -19043
rect 1761 -19103 1771 -19043
rect 1371 -19211 1771 -19103
rect 1827 -19043 2227 -19033
rect 1827 -19103 1837 -19043
rect 1897 -19103 2157 -19043
rect 2217 -19103 2227 -19043
rect 1827 -19211 2227 -19103
rect 2283 -19043 2683 -19033
rect 2283 -19103 2293 -19043
rect 2353 -19103 2613 -19043
rect 2673 -19103 2683 -19043
rect 2283 -19211 2683 -19103
rect 2741 -19043 3141 -19033
rect 2741 -19103 2751 -19043
rect 2811 -19103 3071 -19043
rect 3131 -19103 3141 -19043
rect 2741 -19211 3141 -19103
rect 3197 -19043 3597 -19033
rect 3197 -19103 3207 -19043
rect 3267 -19103 3527 -19043
rect 3587 -19103 3597 -19043
rect 3197 -19211 3597 -19103
rect 457 -19281 3597 -19211
rect 457 -19283 2683 -19281
rect 457 -19393 857 -19283
rect 457 -19453 467 -19393
rect 527 -19453 787 -19393
rect 847 -19453 857 -19393
rect 457 -19463 857 -19453
rect 913 -19393 1313 -19283
rect 913 -19453 923 -19393
rect 983 -19453 1243 -19393
rect 1303 -19453 1313 -19393
rect 913 -19463 1313 -19453
rect 1371 -19393 1771 -19283
rect 1371 -19453 1381 -19393
rect 1441 -19453 1701 -19393
rect 1761 -19453 1771 -19393
rect 1371 -19463 1771 -19453
rect 1827 -19393 2227 -19283
rect 1827 -19453 1837 -19393
rect 1897 -19453 2157 -19393
rect 2217 -19453 2227 -19393
rect 1827 -19463 2227 -19453
rect 2283 -19393 2683 -19283
rect 2283 -19453 2293 -19393
rect 2353 -19453 2613 -19393
rect 2673 -19453 2683 -19393
rect 2283 -19463 2683 -19453
rect 2741 -19283 3597 -19281
rect 2741 -19393 3141 -19283
rect 2741 -19453 2751 -19393
rect 2811 -19453 3071 -19393
rect 3131 -19453 3141 -19393
rect 2741 -19463 3141 -19453
rect 3197 -19393 3597 -19283
rect 3197 -19453 3207 -19393
rect 3267 -19453 3527 -19393
rect 3587 -19453 3597 -19393
rect 3197 -19463 3597 -19453
rect 3653 -19043 4053 -19033
rect 3653 -19103 3663 -19043
rect 3723 -19103 3983 -19043
rect 4043 -19103 4053 -19043
rect 3653 -19211 4053 -19103
rect 4111 -19043 4511 -19033
rect 4111 -19103 4121 -19043
rect 4181 -19103 4441 -19043
rect 4501 -19103 4511 -19043
rect 4111 -19211 4511 -19103
rect 4567 -19043 4967 -19033
rect 4567 -19103 4577 -19043
rect 4637 -19103 4897 -19043
rect 4957 -19103 4967 -19043
rect 4567 -19211 4967 -19103
rect 5023 -19043 5423 -19033
rect 5023 -19103 5033 -19043
rect 5093 -19103 5353 -19043
rect 5413 -19103 5423 -19043
rect 5023 -19211 5423 -19103
rect 5481 -19043 5881 -19033
rect 5481 -19103 5491 -19043
rect 5551 -19103 5811 -19043
rect 5871 -19103 5881 -19043
rect 5481 -19211 5881 -19103
rect 5937 -19043 6337 -19033
rect 5937 -19103 5947 -19043
rect 6007 -19103 6267 -19043
rect 6327 -19103 6337 -19043
rect 5937 -19211 6337 -19103
rect 6393 -19043 6793 -19033
rect 6393 -19103 6403 -19043
rect 6463 -19103 6723 -19043
rect 6783 -19103 6793 -19043
rect 6393 -19211 6793 -19103
rect 6851 -19043 7251 -19033
rect 6851 -19103 6861 -19043
rect 6921 -19103 7181 -19043
rect 7241 -19103 7251 -19043
rect 6851 -19211 7251 -19103
rect 3653 -19283 7251 -19211
rect 3653 -19393 4053 -19283
rect 3653 -19453 3663 -19393
rect 3723 -19453 3983 -19393
rect 4043 -19453 4053 -19393
rect 3653 -19463 4053 -19453
rect 4111 -19393 4511 -19283
rect 4111 -19453 4121 -19393
rect 4181 -19453 4441 -19393
rect 4501 -19453 4511 -19393
rect 4111 -19463 4511 -19453
rect 4567 -19393 4967 -19283
rect 4567 -19453 4577 -19393
rect 4637 -19453 4897 -19393
rect 4957 -19453 4967 -19393
rect 4567 -19463 4967 -19453
rect 5023 -19393 5423 -19283
rect 5023 -19453 5033 -19393
rect 5093 -19453 5353 -19393
rect 5413 -19453 5423 -19393
rect 5023 -19463 5423 -19453
rect 5481 -19393 5881 -19283
rect 5481 -19453 5491 -19393
rect 5551 -19453 5811 -19393
rect 5871 -19453 5881 -19393
rect 5481 -19463 5881 -19453
rect 5937 -19393 6337 -19283
rect 5937 -19453 5947 -19393
rect 6007 -19453 6267 -19393
rect 6327 -19453 6337 -19393
rect 5937 -19463 6337 -19453
rect 6393 -19393 6793 -19283
rect 6393 -19453 6403 -19393
rect 6463 -19453 6723 -19393
rect 6783 -19453 6793 -19393
rect 6393 -19463 6793 -19453
rect 6851 -19393 7251 -19283
rect 6851 -19453 6861 -19393
rect 6921 -19453 7181 -19393
rect 7241 -19453 7251 -19393
rect 6851 -19463 7251 -19453
rect 7307 -19043 7707 -19033
rect 7307 -19103 7317 -19043
rect 7377 -19103 7637 -19043
rect 7697 -19103 7707 -19043
rect 7307 -19211 7707 -19103
rect 7763 -19043 8163 -19033
rect 7763 -19103 7773 -19043
rect 7833 -19103 8093 -19043
rect 8153 -19103 8163 -19043
rect 7763 -19211 8163 -19103
rect 8237 -19043 8637 -19033
rect 8237 -19103 8247 -19043
rect 8307 -19103 8567 -19043
rect 8627 -19103 8637 -19043
rect 8237 -19211 8637 -19103
rect 8693 -19043 9093 -19033
rect 8693 -19103 8703 -19043
rect 8763 -19103 9023 -19043
rect 9083 -19103 9093 -19043
rect 8693 -19211 9093 -19103
rect 9151 -19043 9551 -19033
rect 9151 -19103 9161 -19043
rect 9221 -19103 9481 -19043
rect 9541 -19103 9551 -19043
rect 9151 -19211 9551 -19103
rect 9607 -19043 10007 -19033
rect 9607 -19103 9617 -19043
rect 9677 -19103 9937 -19043
rect 9997 -19103 10007 -19043
rect 9607 -19211 10007 -19103
rect 10063 -19043 10463 -19033
rect 10063 -19103 10073 -19043
rect 10133 -19103 10393 -19043
rect 10453 -19103 10463 -19043
rect 10063 -19211 10463 -19103
rect 10521 -19043 10921 -19033
rect 10521 -19103 10531 -19043
rect 10591 -19103 10851 -19043
rect 10911 -19103 10921 -19043
rect 10521 -19211 10921 -19103
rect 7307 -19283 9093 -19211
rect 9150 -19281 10921 -19211
rect 9150 -19283 10463 -19281
rect 7307 -19393 7707 -19283
rect 7307 -19453 7317 -19393
rect 7377 -19453 7637 -19393
rect 7697 -19453 7707 -19393
rect 7307 -19463 7707 -19453
rect 7763 -19393 8163 -19283
rect 7763 -19453 7773 -19393
rect 7833 -19453 8093 -19393
rect 8153 -19453 8163 -19393
rect 7763 -19463 8163 -19453
rect 8237 -19393 8637 -19283
rect 8237 -19453 8247 -19393
rect 8307 -19453 8567 -19393
rect 8627 -19453 8637 -19393
rect 8237 -19463 8637 -19453
rect 8693 -19393 9093 -19283
rect 8693 -19453 8703 -19393
rect 8763 -19453 9023 -19393
rect 9083 -19453 9093 -19393
rect 8693 -19463 9093 -19453
rect 9151 -19393 9551 -19283
rect 9151 -19453 9161 -19393
rect 9221 -19453 9481 -19393
rect 9541 -19453 9551 -19393
rect 9151 -19463 9551 -19453
rect 9607 -19393 10007 -19283
rect 9607 -19453 9617 -19393
rect 9677 -19453 9937 -19393
rect 9997 -19453 10007 -19393
rect 9607 -19463 10007 -19453
rect 10063 -19393 10463 -19283
rect 10063 -19453 10073 -19393
rect 10133 -19453 10393 -19393
rect 10453 -19453 10463 -19393
rect 10063 -19463 10463 -19453
rect 10521 -19393 10921 -19281
rect 10521 -19453 10531 -19393
rect 10591 -19453 10851 -19393
rect 10911 -19453 10921 -19393
rect 10521 -19463 10921 -19453
rect 10977 -19043 11377 -19033
rect 10977 -19103 10987 -19043
rect 11047 -19103 11307 -19043
rect 11367 -19103 11377 -19043
rect 10977 -19211 11377 -19103
rect 11433 -19043 11833 -19033
rect 11433 -19103 11443 -19043
rect 11503 -19103 11763 -19043
rect 11823 -19103 11833 -19043
rect 11433 -19211 11833 -19103
rect 11891 -19043 12291 -19033
rect 11891 -19103 11901 -19043
rect 11961 -19103 12221 -19043
rect 12281 -19103 12291 -19043
rect 11891 -19211 12291 -19103
rect 12347 -19043 12747 -19033
rect 12347 -19103 12357 -19043
rect 12417 -19103 12677 -19043
rect 12737 -19103 12747 -19043
rect 12347 -19211 12747 -19103
rect 12803 -19043 13203 -19033
rect 12803 -19103 12813 -19043
rect 12873 -19103 13133 -19043
rect 13193 -19103 13203 -19043
rect 12803 -19211 13203 -19103
rect 13261 -19043 13661 -19033
rect 13261 -19103 13271 -19043
rect 13331 -19103 13591 -19043
rect 13651 -19103 13661 -19043
rect 13261 -19211 13661 -19103
rect 13717 -19043 14117 -19033
rect 13717 -19103 13727 -19043
rect 13787 -19103 14047 -19043
rect 14107 -19103 14117 -19043
rect 13717 -19211 14117 -19103
rect 14173 -19043 14573 -19033
rect 14173 -19103 14183 -19043
rect 14243 -19103 14503 -19043
rect 14563 -19103 14573 -19043
rect 14173 -19211 14573 -19103
rect 14631 -19043 15031 -19033
rect 14631 -19103 14641 -19043
rect 14701 -19103 14961 -19043
rect 15021 -19103 15031 -19043
rect 14631 -19211 15031 -19103
rect 15087 -19043 15487 -19033
rect 15087 -19103 15097 -19043
rect 15157 -19103 15417 -19043
rect 15477 -19103 15487 -19043
rect 15087 -19211 15487 -19103
rect 10977 -19283 15487 -19211
rect 10977 -19393 11377 -19283
rect 10977 -19453 10987 -19393
rect 11047 -19453 11307 -19393
rect 11367 -19453 11377 -19393
rect 10977 -19463 11377 -19453
rect 11433 -19393 11833 -19283
rect 11433 -19453 11443 -19393
rect 11503 -19453 11763 -19393
rect 11823 -19453 11833 -19393
rect 11433 -19463 11833 -19453
rect 11891 -19393 12291 -19283
rect 11891 -19453 11901 -19393
rect 11961 -19453 12221 -19393
rect 12281 -19453 12291 -19393
rect 11891 -19463 12291 -19453
rect 12347 -19393 12747 -19283
rect 12347 -19453 12357 -19393
rect 12417 -19453 12677 -19393
rect 12737 -19453 12747 -19393
rect 12347 -19463 12747 -19453
rect 12803 -19393 13203 -19283
rect 12803 -19453 12813 -19393
rect 12873 -19453 13133 -19393
rect 13193 -19453 13203 -19393
rect 12803 -19463 13203 -19453
rect 13261 -19393 13661 -19283
rect 13261 -19453 13271 -19393
rect 13331 -19453 13591 -19393
rect 13651 -19453 13661 -19393
rect 13261 -19463 13661 -19453
rect 13717 -19393 14117 -19283
rect 13717 -19453 13727 -19393
rect 13787 -19453 14047 -19393
rect 14107 -19453 14117 -19393
rect 13717 -19463 14117 -19453
rect 14173 -19393 14573 -19283
rect 14173 -19453 14183 -19393
rect 14243 -19453 14503 -19393
rect 14563 -19453 14573 -19393
rect 14173 -19463 14573 -19453
rect 14631 -19393 15031 -19283
rect 14631 -19453 14641 -19393
rect 14701 -19453 14961 -19393
rect 15021 -19453 15031 -19393
rect 14631 -19463 15031 -19453
rect 15087 -19393 15487 -19283
rect 15087 -19453 15097 -19393
rect 15157 -19453 15417 -19393
rect 15477 -19453 15487 -19393
rect 15087 -19463 15487 -19453
rect 66 -19527 80 -19463
rect 457 -19527 527 -19463
rect 913 -19527 983 -19463
rect 1371 -19527 1441 -19463
rect 1827 -19527 1897 -19463
rect 2283 -19527 2353 -19463
rect 2741 -19527 2811 -19463
rect 3197 -19527 3267 -19463
rect 3653 -19527 3723 -19463
rect 4111 -19527 4181 -19463
rect 4567 -19527 4637 -19463
rect 5023 -19527 5093 -19463
rect 5481 -19527 5551 -19463
rect 5937 -19527 6007 -19463
rect 6393 -19527 6463 -19463
rect 6851 -19527 6921 -19463
rect 7307 -19527 7377 -19463
rect 7763 -19527 7833 -19463
rect 8237 -19527 8307 -19463
rect 8693 -19527 8763 -19463
rect 9151 -19527 9221 -19463
rect 9607 -19527 9677 -19463
rect 10063 -19527 10133 -19463
rect 10521 -19527 10591 -19463
rect 66 -19537 400 -19527
rect 0 -19597 11 -19537
rect 71 -19597 331 -19537
rect 391 -19597 400 -19537
rect 0 -19887 14 -19597
rect 66 -19887 400 -19597
rect 0 -19947 11 -19887
rect 71 -19947 331 -19887
rect 391 -19947 400 -19887
rect 0 -20039 14 -19947
rect 66 -19957 400 -19947
rect 457 -19537 857 -19527
rect 457 -19597 467 -19537
rect 527 -19597 787 -19537
rect 847 -19597 857 -19537
rect 457 -19706 857 -19597
rect 913 -19537 1313 -19527
rect 913 -19597 923 -19537
rect 983 -19597 1243 -19537
rect 1303 -19597 1313 -19537
rect 913 -19706 1313 -19597
rect 1371 -19537 1771 -19527
rect 1371 -19597 1381 -19537
rect 1441 -19597 1701 -19537
rect 1761 -19597 1771 -19537
rect 1371 -19706 1771 -19597
rect 1827 -19537 2227 -19527
rect 1827 -19597 1837 -19537
rect 1897 -19597 2157 -19537
rect 2217 -19597 2227 -19537
rect 1827 -19706 2227 -19597
rect 2283 -19537 2683 -19527
rect 2283 -19597 2293 -19537
rect 2353 -19597 2613 -19537
rect 2673 -19597 2683 -19537
rect 2283 -19706 2683 -19597
rect 2741 -19537 3141 -19527
rect 2741 -19597 2751 -19537
rect 2811 -19597 3071 -19537
rect 3131 -19597 3141 -19537
rect 2741 -19706 3141 -19597
rect 3197 -19537 3597 -19527
rect 3197 -19597 3207 -19537
rect 3267 -19597 3527 -19537
rect 3587 -19597 3597 -19537
rect 3197 -19706 3597 -19597
rect 457 -19776 3597 -19706
rect 457 -19887 857 -19776
rect 457 -19947 467 -19887
rect 527 -19947 787 -19887
rect 847 -19947 857 -19887
rect 457 -19957 857 -19947
rect 913 -19887 1313 -19776
rect 913 -19947 923 -19887
rect 983 -19947 1243 -19887
rect 1303 -19947 1313 -19887
rect 913 -19957 1313 -19947
rect 1371 -19887 1771 -19776
rect 1371 -19947 1381 -19887
rect 1441 -19947 1701 -19887
rect 1761 -19947 1771 -19887
rect 1371 -19957 1771 -19947
rect 1827 -19887 2227 -19776
rect 1827 -19947 1837 -19887
rect 1897 -19947 2157 -19887
rect 2217 -19947 2227 -19887
rect 1827 -19957 2227 -19947
rect 2283 -19887 2683 -19776
rect 2283 -19947 2293 -19887
rect 2353 -19947 2613 -19887
rect 2673 -19947 2683 -19887
rect 2283 -19957 2683 -19947
rect 2741 -19887 3141 -19776
rect 2741 -19947 2751 -19887
rect 2811 -19947 3071 -19887
rect 3131 -19947 3141 -19887
rect 2741 -19957 3141 -19947
rect 3197 -19887 3597 -19776
rect 3197 -19947 3207 -19887
rect 3267 -19947 3527 -19887
rect 3587 -19947 3597 -19887
rect 3197 -19957 3597 -19947
rect 3653 -19537 4053 -19527
rect 3653 -19597 3663 -19537
rect 3723 -19597 3983 -19537
rect 4043 -19597 4053 -19537
rect 3653 -19706 4053 -19597
rect 4111 -19537 4511 -19527
rect 4111 -19597 4121 -19537
rect 4181 -19597 4441 -19537
rect 4501 -19597 4511 -19537
rect 4111 -19706 4511 -19597
rect 4567 -19537 4967 -19527
rect 4567 -19597 4577 -19537
rect 4637 -19597 4897 -19537
rect 4957 -19597 4967 -19537
rect 4567 -19706 4967 -19597
rect 5023 -19537 5423 -19527
rect 5023 -19597 5033 -19537
rect 5093 -19597 5353 -19537
rect 5413 -19597 5423 -19537
rect 5023 -19706 5423 -19597
rect 5481 -19537 5881 -19527
rect 5481 -19597 5491 -19537
rect 5551 -19597 5811 -19537
rect 5871 -19597 5881 -19537
rect 5481 -19706 5881 -19597
rect 5937 -19537 6337 -19527
rect 5937 -19597 5947 -19537
rect 6007 -19597 6267 -19537
rect 6327 -19597 6337 -19537
rect 5937 -19706 6337 -19597
rect 6393 -19537 6793 -19527
rect 6393 -19597 6403 -19537
rect 6463 -19597 6723 -19537
rect 6783 -19597 6793 -19537
rect 6393 -19706 6793 -19597
rect 6851 -19537 7251 -19527
rect 6851 -19597 6861 -19537
rect 6921 -19597 7181 -19537
rect 7241 -19597 7251 -19537
rect 6851 -19706 7251 -19597
rect 3653 -19776 7251 -19706
rect 3653 -19887 4053 -19776
rect 3653 -19947 3663 -19887
rect 3723 -19947 3983 -19887
rect 4043 -19947 4053 -19887
rect 3653 -19957 4053 -19947
rect 4111 -19887 4511 -19776
rect 4111 -19947 4121 -19887
rect 4181 -19947 4441 -19887
rect 4501 -19947 4511 -19887
rect 4111 -19957 4511 -19947
rect 4567 -19887 4967 -19776
rect 4567 -19947 4577 -19887
rect 4637 -19947 4897 -19887
rect 4957 -19947 4967 -19887
rect 4567 -19957 4967 -19947
rect 5023 -19887 5423 -19776
rect 5023 -19947 5033 -19887
rect 5093 -19947 5353 -19887
rect 5413 -19947 5423 -19887
rect 5023 -19957 5423 -19947
rect 5481 -19887 5881 -19776
rect 5481 -19947 5491 -19887
rect 5551 -19947 5811 -19887
rect 5871 -19947 5881 -19887
rect 5481 -19957 5881 -19947
rect 5937 -19887 6337 -19776
rect 5937 -19947 5947 -19887
rect 6007 -19947 6267 -19887
rect 6327 -19947 6337 -19887
rect 5937 -19957 6337 -19947
rect 6393 -19887 6793 -19776
rect 6393 -19947 6403 -19887
rect 6463 -19947 6723 -19887
rect 6783 -19947 6793 -19887
rect 6393 -19957 6793 -19947
rect 6851 -19887 7251 -19776
rect 6851 -19947 6861 -19887
rect 6921 -19947 7181 -19887
rect 7241 -19947 7251 -19887
rect 6851 -19957 7251 -19947
rect 7307 -19537 7707 -19527
rect 7307 -19597 7317 -19537
rect 7377 -19597 7637 -19537
rect 7697 -19597 7707 -19537
rect 7307 -19706 7707 -19597
rect 7763 -19537 8163 -19527
rect 7763 -19597 7773 -19537
rect 7833 -19597 8093 -19537
rect 8153 -19597 8163 -19537
rect 7763 -19706 8163 -19597
rect 8237 -19537 8637 -19527
rect 8237 -19597 8247 -19537
rect 8307 -19597 8567 -19537
rect 8627 -19597 8637 -19537
rect 8237 -19706 8637 -19597
rect 8693 -19537 9093 -19527
rect 8693 -19597 8703 -19537
rect 8763 -19597 9023 -19537
rect 9083 -19597 9093 -19537
rect 8693 -19706 9093 -19597
rect 9151 -19537 9551 -19527
rect 9151 -19597 9161 -19537
rect 9221 -19597 9481 -19537
rect 9541 -19597 9551 -19537
rect 9151 -19706 9551 -19597
rect 9607 -19537 10007 -19527
rect 9607 -19597 9617 -19537
rect 9677 -19597 9937 -19537
rect 9997 -19597 10007 -19537
rect 9607 -19706 10007 -19597
rect 10063 -19537 10463 -19527
rect 10063 -19597 10073 -19537
rect 10133 -19597 10393 -19537
rect 10453 -19597 10463 -19537
rect 10063 -19706 10463 -19597
rect 10521 -19537 10921 -19527
rect 10521 -19597 10531 -19537
rect 10591 -19597 10851 -19537
rect 10911 -19597 10921 -19537
rect 10521 -19706 10921 -19597
rect 10977 -19537 11377 -19527
rect 10977 -19597 10987 -19537
rect 11047 -19597 11307 -19537
rect 11367 -19597 11377 -19537
rect 10977 -19706 11377 -19597
rect 11433 -19537 11833 -19527
rect 11433 -19597 11443 -19537
rect 11503 -19597 11763 -19537
rect 11823 -19597 11833 -19537
rect 11433 -19706 11833 -19597
rect 11891 -19537 12291 -19527
rect 11891 -19597 11901 -19537
rect 11961 -19597 12221 -19537
rect 12281 -19597 12291 -19537
rect 11891 -19706 12291 -19597
rect 12347 -19537 12747 -19527
rect 12347 -19597 12357 -19537
rect 12417 -19597 12677 -19537
rect 12737 -19597 12747 -19537
rect 12347 -19706 12747 -19597
rect 12803 -19537 13203 -19527
rect 12803 -19597 12813 -19537
rect 12873 -19597 13133 -19537
rect 13193 -19597 13203 -19537
rect 12803 -19706 13203 -19597
rect 13261 -19537 13661 -19527
rect 13261 -19597 13271 -19537
rect 13331 -19597 13591 -19537
rect 13651 -19597 13661 -19537
rect 13261 -19706 13661 -19597
rect 13717 -19537 14117 -19527
rect 13717 -19597 13727 -19537
rect 13787 -19597 14047 -19537
rect 14107 -19597 14117 -19537
rect 13717 -19706 14117 -19597
rect 14173 -19537 14573 -19527
rect 14173 -19597 14183 -19537
rect 14243 -19597 14503 -19537
rect 14563 -19597 14573 -19537
rect 14173 -19706 14573 -19597
rect 14631 -19537 15031 -19527
rect 14631 -19597 14641 -19537
rect 14701 -19597 14961 -19537
rect 15021 -19597 15031 -19537
rect 14631 -19706 15031 -19597
rect 15087 -19537 15487 -19527
rect 15087 -19597 15097 -19537
rect 15157 -19597 15417 -19537
rect 15477 -19597 15487 -19537
rect 15087 -19706 15487 -19597
rect 7307 -19776 9093 -19706
rect 9150 -19708 15487 -19706
rect 9150 -19776 15721 -19708
rect 7307 -19887 7707 -19776
rect 7307 -19947 7317 -19887
rect 7377 -19947 7637 -19887
rect 7697 -19947 7707 -19887
rect 7307 -19957 7707 -19947
rect 7763 -19887 8163 -19776
rect 7763 -19947 7773 -19887
rect 7833 -19947 8093 -19887
rect 8153 -19947 8163 -19887
rect 7763 -19957 8163 -19947
rect 8237 -19887 8637 -19776
rect 8237 -19947 8247 -19887
rect 8307 -19947 8567 -19887
rect 8627 -19947 8637 -19887
rect 8237 -19957 8637 -19947
rect 8693 -19887 9093 -19776
rect 8693 -19947 8703 -19887
rect 8763 -19947 9023 -19887
rect 9083 -19947 9093 -19887
rect 8693 -19957 9093 -19947
rect 9151 -19887 9551 -19776
rect 9151 -19947 9161 -19887
rect 9221 -19947 9481 -19887
rect 9541 -19947 9551 -19887
rect 9151 -19957 9551 -19947
rect 9607 -19887 10007 -19776
rect 9607 -19947 9617 -19887
rect 9677 -19947 9937 -19887
rect 9997 -19947 10007 -19887
rect 9607 -19957 10007 -19947
rect 10063 -19887 10463 -19776
rect 10063 -19947 10073 -19887
rect 10133 -19947 10393 -19887
rect 10453 -19947 10463 -19887
rect 10063 -19957 10463 -19947
rect 10521 -19887 10921 -19776
rect 10521 -19947 10531 -19887
rect 10591 -19947 10851 -19887
rect 10911 -19947 10921 -19887
rect 10521 -19957 10921 -19947
rect 10977 -19887 11377 -19776
rect 10977 -19947 10987 -19887
rect 11047 -19947 11307 -19887
rect 11367 -19947 11377 -19887
rect 10977 -19957 11377 -19947
rect 11433 -19887 11833 -19776
rect 11433 -19947 11443 -19887
rect 11503 -19947 11763 -19887
rect 11823 -19947 11833 -19887
rect 11433 -19957 11833 -19947
rect 11891 -19887 12291 -19776
rect 11891 -19947 11901 -19887
rect 11961 -19947 12221 -19887
rect 12281 -19947 12291 -19887
rect 11891 -19957 12291 -19947
rect 12347 -19887 12747 -19776
rect 12347 -19947 12357 -19887
rect 12417 -19947 12677 -19887
rect 12737 -19947 12747 -19887
rect 12347 -19957 12747 -19947
rect 12803 -19887 13203 -19776
rect 12803 -19947 12813 -19887
rect 12873 -19947 13133 -19887
rect 13193 -19947 13203 -19887
rect 12803 -19957 13203 -19947
rect 13261 -19887 13661 -19776
rect 13261 -19947 13271 -19887
rect 13331 -19947 13591 -19887
rect 13651 -19947 13661 -19887
rect 13261 -19957 13661 -19947
rect 13717 -19887 14117 -19776
rect 13717 -19947 13727 -19887
rect 13787 -19947 14047 -19887
rect 14107 -19947 14117 -19887
rect 13717 -19957 14117 -19947
rect 14173 -19887 14573 -19776
rect 14173 -19947 14183 -19887
rect 14243 -19947 14503 -19887
rect 14563 -19947 14573 -19887
rect 14173 -19957 14573 -19947
rect 14631 -19887 15031 -19776
rect 14631 -19947 14641 -19887
rect 14701 -19947 14961 -19887
rect 15021 -19947 15031 -19887
rect 14631 -19957 15031 -19947
rect 15087 -19779 15721 -19776
rect 15087 -19887 15487 -19779
rect 15087 -19947 15097 -19887
rect 15157 -19947 15417 -19887
rect 15477 -19947 15487 -19887
rect 15087 -19957 15487 -19947
rect 66 -20029 80 -19957
rect 457 -20029 527 -19957
rect 913 -20029 984 -19957
rect 1371 -20029 1442 -19957
rect 1827 -20029 1898 -19957
rect 2283 -20029 2354 -19957
rect 2741 -20029 2812 -19957
rect 3197 -20029 3268 -19957
rect 4111 -20029 4182 -19957
rect 4567 -20029 4638 -19957
rect 5023 -20029 5094 -19957
rect 5481 -20029 5552 -19957
rect 5937 -20029 6008 -19957
rect 6393 -20029 6464 -19957
rect 6851 -20029 6922 -19957
rect 7307 -20029 7378 -19957
rect 7763 -20029 7834 -19957
rect 8237 -20029 8308 -19957
rect 8693 -20029 8764 -19957
rect 9607 -20029 9678 -19957
rect 10063 -20029 10134 -19957
rect 10521 -20029 10592 -19957
rect 10977 -20029 11048 -19957
rect 11433 -20029 11504 -19957
rect 11891 -20029 11962 -19957
rect 12347 -20029 12418 -19957
rect 12803 -20029 12874 -19957
rect 13261 -20029 13332 -19957
rect 13717 -20029 13788 -19957
rect 14173 -20029 14244 -19957
rect 14631 -20029 14702 -19957
rect 66 -20039 400 -20029
rect 0 -20099 11 -20039
rect 71 -20099 331 -20039
rect 391 -20099 400 -20039
rect 0 -20389 14 -20099
rect 66 -20389 400 -20099
rect 0 -20449 11 -20389
rect 71 -20449 331 -20389
rect 391 -20449 400 -20389
rect 0 -20531 14 -20449
rect 66 -20459 400 -20449
rect 457 -20039 857 -20029
rect 457 -20099 467 -20039
rect 527 -20099 787 -20039
rect 847 -20099 857 -20039
rect 457 -20209 857 -20099
rect 913 -20039 1313 -20029
rect 913 -20099 923 -20039
rect 983 -20099 1243 -20039
rect 1303 -20099 1313 -20039
rect 913 -20209 1313 -20099
rect 1371 -20039 1771 -20029
rect 1371 -20099 1381 -20039
rect 1441 -20099 1701 -20039
rect 1761 -20099 1771 -20039
rect 1371 -20209 1771 -20099
rect 1827 -20039 2227 -20029
rect 1827 -20099 1837 -20039
rect 1897 -20099 2157 -20039
rect 2217 -20099 2227 -20039
rect 1827 -20209 2227 -20099
rect 2283 -20039 2683 -20029
rect 2283 -20099 2293 -20039
rect 2353 -20099 2613 -20039
rect 2673 -20099 2683 -20039
rect 2283 -20209 2683 -20099
rect 457 -20210 2683 -20209
rect 2741 -20039 3141 -20029
rect 2741 -20099 2751 -20039
rect 2811 -20099 3071 -20039
rect 3131 -20099 3141 -20039
rect 2741 -20209 3141 -20099
rect 3197 -20039 3597 -20029
rect 3197 -20099 3207 -20039
rect 3267 -20099 3527 -20039
rect 3587 -20099 3597 -20039
rect 3197 -20209 3597 -20099
rect 3653 -20039 4053 -20029
rect 3653 -20099 3663 -20039
rect 3723 -20099 3983 -20039
rect 4043 -20099 4053 -20039
rect 3653 -20209 4053 -20099
rect 2741 -20210 4053 -20209
rect 457 -20280 4053 -20210
rect 457 -20389 857 -20280
rect 457 -20449 467 -20389
rect 527 -20449 787 -20389
rect 847 -20449 857 -20389
rect 457 -20459 857 -20449
rect 913 -20389 1313 -20280
rect 913 -20449 923 -20389
rect 983 -20449 1243 -20389
rect 1303 -20449 1313 -20389
rect 913 -20459 1313 -20449
rect 1371 -20389 1771 -20280
rect 1371 -20449 1381 -20389
rect 1441 -20449 1701 -20389
rect 1761 -20449 1771 -20389
rect 1371 -20459 1771 -20449
rect 1827 -20389 2227 -20280
rect 1827 -20449 1837 -20389
rect 1897 -20449 2157 -20389
rect 2217 -20449 2227 -20389
rect 1827 -20459 2227 -20449
rect 2283 -20389 2683 -20280
rect 2283 -20449 2293 -20389
rect 2353 -20449 2613 -20389
rect 2673 -20449 2683 -20389
rect 2283 -20459 2683 -20449
rect 2741 -20389 3141 -20280
rect 2741 -20449 2751 -20389
rect 2811 -20449 3071 -20389
rect 3131 -20449 3141 -20389
rect 2741 -20459 3141 -20449
rect 3197 -20389 3597 -20280
rect 3197 -20449 3207 -20389
rect 3267 -20449 3527 -20389
rect 3587 -20449 3597 -20389
rect 3197 -20459 3597 -20449
rect 3653 -20389 4053 -20280
rect 3653 -20449 3663 -20389
rect 3723 -20449 3983 -20389
rect 4043 -20449 4053 -20389
rect 3653 -20459 4053 -20449
rect 4111 -20039 4511 -20029
rect 4111 -20099 4121 -20039
rect 4181 -20099 4441 -20039
rect 4501 -20099 4511 -20039
rect 4111 -20209 4511 -20099
rect 4567 -20039 4967 -20029
rect 4567 -20099 4577 -20039
rect 4637 -20099 4897 -20039
rect 4957 -20099 4967 -20039
rect 4567 -20209 4967 -20099
rect 5023 -20039 5423 -20029
rect 5023 -20099 5033 -20039
rect 5093 -20099 5353 -20039
rect 5413 -20099 5423 -20039
rect 5023 -20209 5423 -20099
rect 5481 -20039 5881 -20029
rect 5481 -20099 5491 -20039
rect 5551 -20099 5811 -20039
rect 5871 -20099 5881 -20039
rect 5481 -20209 5881 -20099
rect 5937 -20039 6337 -20029
rect 5937 -20099 5947 -20039
rect 6007 -20099 6267 -20039
rect 6327 -20099 6337 -20039
rect 5937 -20209 6337 -20099
rect 6393 -20039 6793 -20029
rect 6393 -20099 6403 -20039
rect 6463 -20099 6723 -20039
rect 6783 -20099 6793 -20039
rect 6393 -20209 6793 -20099
rect 6851 -20039 7251 -20029
rect 6851 -20099 6861 -20039
rect 6921 -20099 7181 -20039
rect 7241 -20099 7251 -20039
rect 6851 -20209 7251 -20099
rect 4111 -20280 7251 -20209
rect 4111 -20389 4511 -20280
rect 4111 -20449 4121 -20389
rect 4181 -20449 4441 -20389
rect 4501 -20449 4511 -20389
rect 4111 -20459 4511 -20449
rect 4567 -20389 4967 -20280
rect 4567 -20449 4577 -20389
rect 4637 -20449 4897 -20389
rect 4957 -20449 4967 -20389
rect 4567 -20459 4967 -20449
rect 5023 -20389 5423 -20280
rect 5023 -20449 5033 -20389
rect 5093 -20449 5353 -20389
rect 5413 -20449 5423 -20389
rect 5023 -20459 5423 -20449
rect 5481 -20389 5881 -20280
rect 5481 -20449 5491 -20389
rect 5551 -20449 5811 -20389
rect 5871 -20449 5881 -20389
rect 5481 -20459 5881 -20449
rect 5937 -20389 6337 -20280
rect 5937 -20449 5947 -20389
rect 6007 -20449 6267 -20389
rect 6327 -20449 6337 -20389
rect 5937 -20459 6337 -20449
rect 6393 -20389 6793 -20280
rect 6393 -20449 6403 -20389
rect 6463 -20449 6723 -20389
rect 6783 -20449 6793 -20389
rect 6393 -20459 6793 -20449
rect 6851 -20389 7251 -20280
rect 6851 -20449 6861 -20389
rect 6921 -20449 7181 -20389
rect 7241 -20449 7251 -20389
rect 6851 -20459 7251 -20449
rect 7307 -20039 7707 -20029
rect 7307 -20099 7317 -20039
rect 7377 -20099 7637 -20039
rect 7697 -20099 7707 -20039
rect 7307 -20209 7707 -20099
rect 7763 -20039 8163 -20029
rect 7763 -20099 7773 -20039
rect 7833 -20099 8093 -20039
rect 8153 -20099 8163 -20039
rect 7763 -20209 8163 -20099
rect 8237 -20039 8637 -20029
rect 8237 -20099 8247 -20039
rect 8307 -20099 8567 -20039
rect 8627 -20099 8637 -20039
rect 8237 -20209 8637 -20099
rect 8693 -20039 9093 -20029
rect 8693 -20099 8703 -20039
rect 8763 -20099 9023 -20039
rect 9083 -20099 9093 -20039
rect 8693 -20209 9093 -20099
rect 9151 -20039 9551 -20029
rect 9151 -20099 9161 -20039
rect 9221 -20099 9481 -20039
rect 9541 -20099 9551 -20039
rect 9151 -20209 9551 -20099
rect 7307 -20280 9551 -20209
rect 7307 -20389 7707 -20280
rect 7307 -20449 7317 -20389
rect 7377 -20449 7637 -20389
rect 7697 -20449 7707 -20389
rect 7307 -20459 7707 -20449
rect 7763 -20389 8163 -20280
rect 7763 -20449 7773 -20389
rect 7833 -20449 8093 -20389
rect 8153 -20449 8163 -20389
rect 7763 -20459 8163 -20449
rect 8237 -20389 8637 -20280
rect 8237 -20449 8247 -20389
rect 8307 -20449 8567 -20389
rect 8627 -20449 8637 -20389
rect 8237 -20459 8637 -20449
rect 8693 -20389 9093 -20280
rect 8693 -20449 8703 -20389
rect 8763 -20449 9023 -20389
rect 9083 -20449 9093 -20389
rect 8693 -20459 9093 -20449
rect 9151 -20389 9551 -20280
rect 9151 -20449 9161 -20389
rect 9221 -20449 9481 -20389
rect 9541 -20449 9551 -20389
rect 9151 -20459 9551 -20449
rect 9607 -20039 10007 -20029
rect 9607 -20099 9617 -20039
rect 9677 -20099 9937 -20039
rect 9997 -20099 10007 -20039
rect 9607 -20209 10007 -20099
rect 10063 -20039 10463 -20029
rect 10063 -20099 10073 -20039
rect 10133 -20099 10393 -20039
rect 10453 -20099 10463 -20039
rect 10063 -20209 10463 -20099
rect 9607 -20210 10463 -20209
rect 10521 -20039 10921 -20029
rect 10521 -20099 10531 -20039
rect 10591 -20099 10851 -20039
rect 10911 -20099 10921 -20039
rect 10521 -20209 10921 -20099
rect 10977 -20039 11377 -20029
rect 10977 -20099 10987 -20039
rect 11047 -20099 11307 -20039
rect 11367 -20099 11377 -20039
rect 10977 -20209 11377 -20099
rect 11433 -20039 11833 -20029
rect 11433 -20099 11443 -20039
rect 11503 -20099 11763 -20039
rect 11823 -20099 11833 -20039
rect 11433 -20209 11833 -20099
rect 11891 -20039 12291 -20029
rect 11891 -20099 11901 -20039
rect 11961 -20099 12221 -20039
rect 12281 -20099 12291 -20039
rect 11891 -20209 12291 -20099
rect 12347 -20039 12747 -20029
rect 12347 -20099 12357 -20039
rect 12417 -20099 12677 -20039
rect 12737 -20099 12747 -20039
rect 12347 -20209 12747 -20099
rect 12803 -20039 13203 -20029
rect 12803 -20099 12813 -20039
rect 12873 -20099 13133 -20039
rect 13193 -20099 13203 -20039
rect 12803 -20209 13203 -20099
rect 13261 -20039 13661 -20029
rect 13261 -20099 13271 -20039
rect 13331 -20099 13591 -20039
rect 13651 -20099 13661 -20039
rect 13261 -20209 13661 -20099
rect 13717 -20039 14117 -20029
rect 13717 -20099 13727 -20039
rect 13787 -20099 14047 -20039
rect 14107 -20099 14117 -20039
rect 13717 -20209 14117 -20099
rect 14173 -20039 14573 -20029
rect 14173 -20099 14183 -20039
rect 14243 -20099 14503 -20039
rect 14563 -20099 14573 -20039
rect 14173 -20209 14573 -20099
rect 14631 -20039 15031 -20029
rect 14631 -20099 14641 -20039
rect 14701 -20099 14961 -20039
rect 15021 -20099 15031 -20039
rect 14631 -20209 15031 -20099
rect 15087 -20039 15487 -20029
rect 15087 -20099 15097 -20039
rect 15157 -20099 15417 -20039
rect 15477 -20099 15487 -20039
rect 15087 -20209 15487 -20099
rect 10521 -20210 15487 -20209
rect 9607 -20280 15487 -20210
rect 9607 -20389 10007 -20280
rect 9607 -20449 9617 -20389
rect 9677 -20449 9937 -20389
rect 9997 -20449 10007 -20389
rect 9607 -20459 10007 -20449
rect 10063 -20389 10463 -20280
rect 10063 -20449 10073 -20389
rect 10133 -20449 10393 -20389
rect 10453 -20449 10463 -20389
rect 10063 -20459 10463 -20449
rect 10521 -20389 10921 -20280
rect 10521 -20449 10531 -20389
rect 10591 -20449 10851 -20389
rect 10911 -20449 10921 -20389
rect 10521 -20459 10921 -20449
rect 10977 -20389 11377 -20280
rect 10977 -20449 10987 -20389
rect 11047 -20449 11307 -20389
rect 11367 -20449 11377 -20389
rect 10977 -20459 11377 -20449
rect 11433 -20389 11833 -20280
rect 11433 -20449 11443 -20389
rect 11503 -20449 11763 -20389
rect 11823 -20449 11833 -20389
rect 11433 -20459 11833 -20449
rect 11891 -20389 12291 -20280
rect 11891 -20449 11901 -20389
rect 11961 -20449 12221 -20389
rect 12281 -20449 12291 -20389
rect 11891 -20459 12291 -20449
rect 12347 -20389 12747 -20280
rect 12347 -20449 12357 -20389
rect 12417 -20449 12677 -20389
rect 12737 -20449 12747 -20389
rect 12347 -20459 12747 -20449
rect 12803 -20389 13203 -20280
rect 12803 -20449 12813 -20389
rect 12873 -20449 13133 -20389
rect 13193 -20449 13203 -20389
rect 12803 -20459 13203 -20449
rect 13261 -20389 13661 -20280
rect 13261 -20449 13271 -20389
rect 13331 -20449 13591 -20389
rect 13651 -20449 13661 -20389
rect 13261 -20459 13661 -20449
rect 13717 -20389 14117 -20280
rect 13717 -20449 13727 -20389
rect 13787 -20449 14047 -20389
rect 14107 -20449 14117 -20389
rect 13717 -20459 14117 -20449
rect 14173 -20389 14573 -20280
rect 14173 -20449 14183 -20389
rect 14243 -20449 14503 -20389
rect 14563 -20449 14573 -20389
rect 14173 -20459 14573 -20449
rect 14631 -20389 15031 -20280
rect 14631 -20449 14641 -20389
rect 14701 -20449 14961 -20389
rect 15021 -20449 15031 -20389
rect 14631 -20459 15031 -20449
rect 15087 -20389 15487 -20280
rect 15087 -20449 15097 -20389
rect 15157 -20449 15417 -20389
rect 15477 -20449 15487 -20389
rect 15087 -20459 15487 -20449
rect 66 -20521 80 -20459
rect 457 -20521 528 -20459
rect 913 -20521 984 -20459
rect 1371 -20521 1442 -20459
rect 1827 -20521 1898 -20459
rect 2283 -20521 2354 -20459
rect 2741 -20521 2811 -20459
rect 3197 -20521 3267 -20459
rect 3653 -20521 3723 -20459
rect 4111 -20521 4181 -20459
rect 4567 -20521 4637 -20459
rect 5023 -20521 5093 -20459
rect 5481 -20521 5551 -20459
rect 5937 -20521 6007 -20459
rect 6393 -20521 6463 -20459
rect 6851 -20521 6921 -20459
rect 7307 -20521 7377 -20459
rect 7763 -20521 7833 -20459
rect 8237 -20521 8307 -20459
rect 8693 -20521 8763 -20459
rect 9151 -20521 9221 -20459
rect 9607 -20521 9677 -20459
rect 10063 -20521 10133 -20459
rect 10521 -20521 10591 -20459
rect 10977 -20521 11047 -20459
rect 11433 -20521 11503 -20459
rect 11891 -20521 11961 -20459
rect 12347 -20521 12417 -20459
rect 12803 -20521 12873 -20459
rect 13261 -20521 13331 -20459
rect 13717 -20521 13787 -20459
rect 14173 -20521 14243 -20459
rect 14631 -20521 14701 -20459
rect 66 -20531 400 -20521
rect 0 -20591 11 -20531
rect 71 -20591 331 -20531
rect 391 -20591 400 -20531
rect 0 -20881 14 -20591
rect 66 -20881 400 -20591
rect 0 -20941 11 -20881
rect 71 -20941 331 -20881
rect 391 -20941 400 -20881
rect 0 -21047 14 -20941
rect 66 -20951 400 -20941
rect 457 -20531 857 -20521
rect 457 -20591 467 -20531
rect 527 -20591 787 -20531
rect 847 -20591 857 -20531
rect 457 -20699 857 -20591
rect 913 -20531 1313 -20521
rect 913 -20591 923 -20531
rect 983 -20591 1243 -20531
rect 1303 -20591 1313 -20531
rect 913 -20699 1313 -20591
rect 1371 -20531 1771 -20521
rect 1371 -20591 1381 -20531
rect 1441 -20591 1701 -20531
rect 1761 -20591 1771 -20531
rect 1371 -20699 1771 -20591
rect 1827 -20531 2227 -20521
rect 1827 -20591 1837 -20531
rect 1897 -20591 2157 -20531
rect 2217 -20591 2227 -20531
rect 1827 -20699 2227 -20591
rect 2283 -20531 2683 -20521
rect 2283 -20591 2293 -20531
rect 2353 -20591 2613 -20531
rect 2673 -20591 2683 -20531
rect 2283 -20699 2683 -20591
rect 2741 -20531 3141 -20521
rect 2741 -20591 2751 -20531
rect 2811 -20591 3071 -20531
rect 3131 -20591 3141 -20531
rect 2741 -20699 3141 -20591
rect 3197 -20531 3597 -20521
rect 3197 -20591 3207 -20531
rect 3267 -20591 3527 -20531
rect 3587 -20591 3597 -20531
rect 3197 -20699 3597 -20591
rect 3653 -20531 4053 -20521
rect 3653 -20591 3663 -20531
rect 3723 -20591 3983 -20531
rect 4043 -20591 4053 -20531
rect 3653 -20699 4053 -20591
rect 457 -20769 4053 -20699
rect 457 -20771 2683 -20769
rect 457 -20881 857 -20771
rect 457 -20941 467 -20881
rect 527 -20941 787 -20881
rect 847 -20941 857 -20881
rect 457 -20951 857 -20941
rect 913 -20881 1313 -20771
rect 913 -20941 923 -20881
rect 983 -20941 1243 -20881
rect 1303 -20941 1313 -20881
rect 913 -20951 1313 -20941
rect 1371 -20881 1771 -20771
rect 1371 -20941 1381 -20881
rect 1441 -20941 1701 -20881
rect 1761 -20941 1771 -20881
rect 1371 -20951 1771 -20941
rect 1827 -20881 2227 -20771
rect 1827 -20941 1837 -20881
rect 1897 -20941 2157 -20881
rect 2217 -20941 2227 -20881
rect 1827 -20951 2227 -20941
rect 2283 -20881 2683 -20771
rect 2283 -20941 2293 -20881
rect 2353 -20941 2613 -20881
rect 2673 -20941 2683 -20881
rect 2283 -20951 2683 -20941
rect 2741 -20771 4053 -20769
rect 2741 -20881 3141 -20771
rect 2741 -20941 2751 -20881
rect 2811 -20941 3071 -20881
rect 3131 -20941 3141 -20881
rect 2741 -20951 3141 -20941
rect 3197 -20881 3597 -20771
rect 3197 -20941 3207 -20881
rect 3267 -20941 3527 -20881
rect 3587 -20941 3597 -20881
rect 3197 -20951 3597 -20941
rect 3653 -20881 4053 -20771
rect 3653 -20941 3663 -20881
rect 3723 -20941 3983 -20881
rect 4043 -20941 4053 -20881
rect 3653 -20951 4053 -20941
rect 4111 -20531 4511 -20521
rect 4111 -20591 4121 -20531
rect 4181 -20591 4441 -20531
rect 4501 -20591 4511 -20531
rect 4111 -20699 4511 -20591
rect 4567 -20531 4967 -20521
rect 4567 -20591 4577 -20531
rect 4637 -20591 4897 -20531
rect 4957 -20591 4967 -20531
rect 4567 -20699 4967 -20591
rect 5023 -20531 5423 -20521
rect 5023 -20591 5033 -20531
rect 5093 -20591 5353 -20531
rect 5413 -20591 5423 -20531
rect 5023 -20699 5423 -20591
rect 5481 -20531 5881 -20521
rect 5481 -20591 5491 -20531
rect 5551 -20591 5811 -20531
rect 5871 -20591 5881 -20531
rect 5481 -20699 5881 -20591
rect 5937 -20531 6337 -20521
rect 5937 -20591 5947 -20531
rect 6007 -20591 6267 -20531
rect 6327 -20591 6337 -20531
rect 5937 -20699 6337 -20591
rect 6393 -20531 6793 -20521
rect 6393 -20591 6403 -20531
rect 6463 -20591 6723 -20531
rect 6783 -20591 6793 -20531
rect 6393 -20699 6793 -20591
rect 6851 -20531 7251 -20521
rect 6851 -20591 6861 -20531
rect 6921 -20591 7181 -20531
rect 7241 -20591 7251 -20531
rect 6851 -20699 7251 -20591
rect 4111 -20771 7251 -20699
rect 4111 -20881 4511 -20771
rect 4111 -20941 4121 -20881
rect 4181 -20941 4441 -20881
rect 4501 -20941 4511 -20881
rect 4111 -20951 4511 -20941
rect 4567 -20881 4967 -20771
rect 4567 -20941 4577 -20881
rect 4637 -20941 4897 -20881
rect 4957 -20941 4967 -20881
rect 4567 -20951 4967 -20941
rect 5023 -20881 5423 -20771
rect 5023 -20941 5033 -20881
rect 5093 -20941 5353 -20881
rect 5413 -20941 5423 -20881
rect 5023 -20951 5423 -20941
rect 5481 -20881 5881 -20771
rect 5481 -20941 5491 -20881
rect 5551 -20941 5811 -20881
rect 5871 -20941 5881 -20881
rect 5481 -20951 5881 -20941
rect 5937 -20881 6337 -20771
rect 5937 -20941 5947 -20881
rect 6007 -20941 6267 -20881
rect 6327 -20941 6337 -20881
rect 5937 -20951 6337 -20941
rect 6393 -20881 6793 -20771
rect 6393 -20941 6403 -20881
rect 6463 -20941 6723 -20881
rect 6783 -20941 6793 -20881
rect 6393 -20951 6793 -20941
rect 6851 -20881 7251 -20771
rect 6851 -20941 6861 -20881
rect 6921 -20941 7181 -20881
rect 7241 -20941 7251 -20881
rect 6851 -20951 7251 -20941
rect 7307 -20531 7707 -20521
rect 7307 -20591 7317 -20531
rect 7377 -20591 7637 -20531
rect 7697 -20591 7707 -20531
rect 7307 -20699 7707 -20591
rect 7763 -20531 8163 -20521
rect 7763 -20591 7773 -20531
rect 7833 -20591 8093 -20531
rect 8153 -20591 8163 -20531
rect 7763 -20699 8163 -20591
rect 8237 -20531 8637 -20521
rect 8237 -20591 8247 -20531
rect 8307 -20591 8567 -20531
rect 8627 -20591 8637 -20531
rect 8237 -20699 8637 -20591
rect 8693 -20531 9093 -20521
rect 8693 -20591 8703 -20531
rect 8763 -20591 9023 -20531
rect 9083 -20591 9093 -20531
rect 8693 -20699 9093 -20591
rect 9151 -20531 9551 -20521
rect 9151 -20591 9161 -20531
rect 9221 -20591 9481 -20531
rect 9541 -20591 9551 -20531
rect 9151 -20699 9551 -20591
rect 7307 -20771 9551 -20699
rect 7307 -20881 7707 -20771
rect 7307 -20941 7317 -20881
rect 7377 -20941 7637 -20881
rect 7697 -20941 7707 -20881
rect 7307 -20951 7707 -20941
rect 7763 -20881 8163 -20771
rect 7763 -20941 7773 -20881
rect 7833 -20941 8093 -20881
rect 8153 -20941 8163 -20881
rect 7763 -20951 8163 -20941
rect 8237 -20881 8637 -20771
rect 8237 -20941 8247 -20881
rect 8307 -20941 8567 -20881
rect 8627 -20941 8637 -20881
rect 8237 -20951 8637 -20941
rect 8693 -20881 9093 -20771
rect 8693 -20941 8703 -20881
rect 8763 -20941 9023 -20881
rect 9083 -20941 9093 -20881
rect 8693 -20951 9093 -20941
rect 9151 -20881 9551 -20771
rect 9151 -20941 9161 -20881
rect 9221 -20941 9481 -20881
rect 9541 -20941 9551 -20881
rect 9151 -20951 9551 -20941
rect 9607 -20531 10007 -20521
rect 9607 -20591 9617 -20531
rect 9677 -20591 9937 -20531
rect 9997 -20591 10007 -20531
rect 9607 -20699 10007 -20591
rect 10063 -20531 10463 -20521
rect 10063 -20591 10073 -20531
rect 10133 -20591 10393 -20531
rect 10453 -20591 10463 -20531
rect 10063 -20699 10463 -20591
rect 10521 -20531 10921 -20521
rect 10521 -20591 10531 -20531
rect 10591 -20591 10851 -20531
rect 10911 -20591 10921 -20531
rect 10521 -20699 10921 -20591
rect 10977 -20531 11377 -20521
rect 10977 -20591 10987 -20531
rect 11047 -20591 11307 -20531
rect 11367 -20591 11377 -20531
rect 10977 -20699 11377 -20591
rect 11433 -20531 11833 -20521
rect 11433 -20591 11443 -20531
rect 11503 -20591 11763 -20531
rect 11823 -20591 11833 -20531
rect 11433 -20699 11833 -20591
rect 11891 -20531 12291 -20521
rect 11891 -20591 11901 -20531
rect 11961 -20591 12221 -20531
rect 12281 -20591 12291 -20531
rect 11891 -20699 12291 -20591
rect 12347 -20531 12747 -20521
rect 12347 -20591 12357 -20531
rect 12417 -20591 12677 -20531
rect 12737 -20591 12747 -20531
rect 12347 -20699 12747 -20591
rect 12803 -20531 13203 -20521
rect 12803 -20591 12813 -20531
rect 12873 -20591 13133 -20531
rect 13193 -20591 13203 -20531
rect 12803 -20699 13203 -20591
rect 13261 -20531 13661 -20521
rect 13261 -20591 13271 -20531
rect 13331 -20591 13591 -20531
rect 13651 -20591 13661 -20531
rect 13261 -20699 13661 -20591
rect 13717 -20531 14117 -20521
rect 13717 -20591 13727 -20531
rect 13787 -20591 14047 -20531
rect 14107 -20591 14117 -20531
rect 13717 -20699 14117 -20591
rect 14173 -20531 14573 -20521
rect 14173 -20591 14183 -20531
rect 14243 -20591 14503 -20531
rect 14563 -20591 14573 -20531
rect 14173 -20699 14573 -20591
rect 14631 -20531 15031 -20521
rect 14631 -20591 14641 -20531
rect 14701 -20591 14961 -20531
rect 15021 -20591 15031 -20531
rect 14631 -20699 15031 -20591
rect 15087 -20531 15487 -20521
rect 15087 -20591 15097 -20531
rect 15157 -20591 15417 -20531
rect 15477 -20591 15487 -20531
rect 15087 -20699 15487 -20591
rect 9607 -20769 15487 -20699
rect 9607 -20771 10463 -20769
rect 9607 -20881 10007 -20771
rect 9607 -20941 9617 -20881
rect 9677 -20941 9937 -20881
rect 9997 -20941 10007 -20881
rect 9607 -20951 10007 -20941
rect 10063 -20881 10463 -20771
rect 10063 -20941 10073 -20881
rect 10133 -20941 10393 -20881
rect 10453 -20941 10463 -20881
rect 10063 -20951 10463 -20941
rect 10521 -20771 15487 -20769
rect 10521 -20881 10921 -20771
rect 10521 -20941 10531 -20881
rect 10591 -20941 10851 -20881
rect 10911 -20941 10921 -20881
rect 10521 -20951 10921 -20941
rect 10977 -20881 11377 -20771
rect 10977 -20941 10987 -20881
rect 11047 -20941 11307 -20881
rect 11367 -20941 11377 -20881
rect 10977 -20951 11377 -20941
rect 11433 -20881 11833 -20771
rect 11433 -20941 11443 -20881
rect 11503 -20941 11763 -20881
rect 11823 -20941 11833 -20881
rect 11433 -20951 11833 -20941
rect 11891 -20881 12291 -20771
rect 11891 -20941 11901 -20881
rect 11961 -20941 12221 -20881
rect 12281 -20941 12291 -20881
rect 11891 -20951 12291 -20941
rect 12347 -20881 12747 -20771
rect 12347 -20941 12357 -20881
rect 12417 -20941 12677 -20881
rect 12737 -20941 12747 -20881
rect 12347 -20951 12747 -20941
rect 12803 -20881 13203 -20771
rect 12803 -20941 12813 -20881
rect 12873 -20941 13133 -20881
rect 13193 -20941 13203 -20881
rect 12803 -20951 13203 -20941
rect 13261 -20881 13661 -20771
rect 13261 -20941 13271 -20881
rect 13331 -20941 13591 -20881
rect 13651 -20941 13661 -20881
rect 13261 -20951 13661 -20941
rect 13717 -20881 14117 -20771
rect 13717 -20941 13727 -20881
rect 13787 -20941 14047 -20881
rect 14107 -20941 14117 -20881
rect 13717 -20951 14117 -20941
rect 14173 -20881 14573 -20771
rect 14173 -20941 14183 -20881
rect 14243 -20941 14503 -20881
rect 14563 -20941 14573 -20881
rect 14173 -20951 14573 -20941
rect 14631 -20881 15031 -20771
rect 14631 -20941 14641 -20881
rect 14701 -20941 14961 -20881
rect 15021 -20941 15031 -20881
rect 14631 -20951 15031 -20941
rect 15087 -20881 15487 -20771
rect 15087 -20941 15097 -20881
rect 15157 -20941 15417 -20881
rect 15477 -20941 15487 -20881
rect 15087 -20951 15487 -20941
rect 66 -21037 80 -20951
rect 457 -21037 527 -20951
rect 913 -21037 983 -20951
rect 1371 -21037 1441 -20951
rect 1827 -21037 1897 -20951
rect 2283 -21037 2353 -20951
rect 2741 -21037 2811 -20951
rect 3197 -21037 3267 -20951
rect 3653 -21037 3723 -20951
rect 4111 -21037 4181 -20951
rect 4567 -21037 4637 -20951
rect 5023 -21037 5093 -20951
rect 5481 -21037 5551 -20951
rect 5937 -21037 6007 -20951
rect 6393 -21037 6463 -20951
rect 6851 -21037 6921 -20951
rect 7307 -21037 7377 -20951
rect 7763 -21037 7833 -20951
rect 8237 -21037 8307 -20951
rect 8693 -21037 8763 -20951
rect 9151 -21037 9221 -20951
rect 66 -21047 400 -21037
rect 0 -21107 11 -21047
rect 71 -21107 331 -21047
rect 391 -21107 400 -21047
rect 0 -21397 14 -21107
rect 66 -21397 400 -21107
rect 0 -21457 11 -21397
rect 71 -21457 331 -21397
rect 391 -21457 400 -21397
rect 0 -21549 14 -21457
rect 66 -21467 400 -21457
rect 457 -21047 857 -21037
rect 457 -21107 467 -21047
rect 527 -21107 787 -21047
rect 847 -21107 857 -21047
rect 457 -21217 857 -21107
rect 913 -21047 1313 -21037
rect 913 -21107 923 -21047
rect 983 -21107 1243 -21047
rect 1303 -21107 1313 -21047
rect 913 -21217 1313 -21107
rect 1371 -21047 1771 -21037
rect 1371 -21107 1381 -21047
rect 1441 -21107 1701 -21047
rect 1761 -21107 1771 -21047
rect 1371 -21217 1771 -21107
rect 1827 -21047 2227 -21037
rect 1827 -21107 1837 -21047
rect 1897 -21107 2157 -21047
rect 2217 -21107 2227 -21047
rect 1827 -21217 2227 -21107
rect 2283 -21047 2683 -21037
rect 2283 -21107 2293 -21047
rect 2353 -21107 2613 -21047
rect 2673 -21107 2683 -21047
rect 2283 -21217 2683 -21107
rect 457 -21219 2683 -21217
rect 2741 -21047 3141 -21037
rect 2741 -21107 2751 -21047
rect 2811 -21107 3071 -21047
rect 3131 -21107 3141 -21047
rect 2741 -21217 3141 -21107
rect 3197 -21047 3597 -21037
rect 3197 -21107 3207 -21047
rect 3267 -21107 3527 -21047
rect 3587 -21107 3597 -21047
rect 3197 -21217 3597 -21107
rect 3653 -21047 4053 -21037
rect 3653 -21107 3663 -21047
rect 3723 -21107 3983 -21047
rect 4043 -21107 4053 -21047
rect 3653 -21217 4053 -21107
rect 2741 -21219 4053 -21217
rect 457 -21289 4053 -21219
rect 457 -21397 857 -21289
rect 457 -21457 467 -21397
rect 527 -21457 787 -21397
rect 847 -21457 857 -21397
rect 457 -21467 857 -21457
rect 913 -21397 1313 -21289
rect 913 -21457 923 -21397
rect 983 -21457 1243 -21397
rect 1303 -21457 1313 -21397
rect 913 -21467 1313 -21457
rect 1371 -21397 1771 -21289
rect 1371 -21457 1381 -21397
rect 1441 -21457 1701 -21397
rect 1761 -21457 1771 -21397
rect 1371 -21467 1771 -21457
rect 1827 -21397 2227 -21289
rect 1827 -21457 1837 -21397
rect 1897 -21457 2157 -21397
rect 2217 -21457 2227 -21397
rect 1827 -21467 2227 -21457
rect 2283 -21397 2683 -21289
rect 2283 -21457 2293 -21397
rect 2353 -21457 2613 -21397
rect 2673 -21457 2683 -21397
rect 2283 -21467 2683 -21457
rect 2741 -21397 3141 -21289
rect 2741 -21457 2751 -21397
rect 2811 -21457 3071 -21397
rect 3131 -21457 3141 -21397
rect 2741 -21467 3141 -21457
rect 3197 -21397 3597 -21289
rect 3197 -21457 3207 -21397
rect 3267 -21457 3527 -21397
rect 3587 -21457 3597 -21397
rect 3197 -21467 3597 -21457
rect 3653 -21397 4053 -21289
rect 3653 -21457 3663 -21397
rect 3723 -21457 3983 -21397
rect 4043 -21457 4053 -21397
rect 3653 -21467 4053 -21457
rect 4111 -21047 4511 -21037
rect 4111 -21107 4121 -21047
rect 4181 -21107 4441 -21047
rect 4501 -21107 4511 -21047
rect 4111 -21217 4511 -21107
rect 4567 -21047 4967 -21037
rect 4567 -21107 4577 -21047
rect 4637 -21107 4897 -21047
rect 4957 -21107 4967 -21047
rect 4567 -21217 4967 -21107
rect 5023 -21047 5423 -21037
rect 5023 -21107 5033 -21047
rect 5093 -21107 5353 -21047
rect 5413 -21107 5423 -21047
rect 5023 -21217 5423 -21107
rect 5481 -21047 5881 -21037
rect 5481 -21107 5491 -21047
rect 5551 -21107 5811 -21047
rect 5871 -21107 5881 -21047
rect 5481 -21217 5881 -21107
rect 5937 -21047 6337 -21037
rect 5937 -21107 5947 -21047
rect 6007 -21107 6267 -21047
rect 6327 -21107 6337 -21047
rect 5937 -21217 6337 -21107
rect 6393 -21047 6793 -21037
rect 6393 -21107 6403 -21047
rect 6463 -21107 6723 -21047
rect 6783 -21107 6793 -21047
rect 6393 -21217 6793 -21107
rect 6851 -21047 7251 -21037
rect 6851 -21107 6861 -21047
rect 6921 -21107 7181 -21047
rect 7241 -21107 7251 -21047
rect 6851 -21217 7251 -21107
rect 4111 -21289 7251 -21217
rect 4111 -21397 4511 -21289
rect 4111 -21457 4121 -21397
rect 4181 -21457 4441 -21397
rect 4501 -21457 4511 -21397
rect 4111 -21467 4511 -21457
rect 4567 -21397 4967 -21289
rect 4567 -21457 4577 -21397
rect 4637 -21457 4897 -21397
rect 4957 -21457 4967 -21397
rect 4567 -21467 4967 -21457
rect 5023 -21397 5423 -21289
rect 5023 -21457 5033 -21397
rect 5093 -21457 5353 -21397
rect 5413 -21457 5423 -21397
rect 5023 -21467 5423 -21457
rect 5481 -21397 5881 -21289
rect 5481 -21457 5491 -21397
rect 5551 -21457 5811 -21397
rect 5871 -21457 5881 -21397
rect 5481 -21467 5881 -21457
rect 5937 -21397 6337 -21289
rect 5937 -21457 5947 -21397
rect 6007 -21457 6267 -21397
rect 6327 -21457 6337 -21397
rect 5937 -21467 6337 -21457
rect 6393 -21397 6793 -21289
rect 6393 -21457 6403 -21397
rect 6463 -21457 6723 -21397
rect 6783 -21457 6793 -21397
rect 6393 -21467 6793 -21457
rect 6851 -21397 7251 -21289
rect 6851 -21457 6861 -21397
rect 6921 -21457 7181 -21397
rect 7241 -21457 7251 -21397
rect 6851 -21467 7251 -21457
rect 7307 -21047 7707 -21037
rect 7307 -21107 7317 -21047
rect 7377 -21107 7637 -21047
rect 7697 -21107 7707 -21047
rect 7307 -21217 7707 -21107
rect 7763 -21047 8163 -21037
rect 7763 -21107 7773 -21047
rect 7833 -21107 8093 -21047
rect 8153 -21107 8163 -21047
rect 7763 -21217 8163 -21107
rect 8237 -21047 8637 -21037
rect 8237 -21107 8247 -21047
rect 8307 -21107 8567 -21047
rect 8627 -21107 8637 -21047
rect 8237 -21217 8637 -21107
rect 8693 -21047 9093 -21037
rect 8693 -21107 8703 -21047
rect 8763 -21107 9023 -21047
rect 9083 -21107 9093 -21047
rect 8693 -21217 9093 -21107
rect 9151 -21047 9551 -21037
rect 9151 -21107 9161 -21047
rect 9221 -21107 9481 -21047
rect 9541 -21107 9551 -21047
rect 9151 -21217 9551 -21107
rect 9607 -21047 10007 -21037
rect 9607 -21107 9617 -21047
rect 9677 -21107 9937 -21047
rect 9997 -21107 10007 -21047
rect 9607 -21217 10007 -21107
rect 10063 -21047 10463 -21037
rect 10063 -21107 10073 -21047
rect 10133 -21107 10393 -21047
rect 10453 -21107 10463 -21047
rect 10063 -21217 10463 -21107
rect 7307 -21219 10463 -21217
rect 10521 -21047 10921 -21037
rect 10521 -21107 10531 -21047
rect 10591 -21107 10851 -21047
rect 10911 -21107 10921 -21047
rect 10521 -21217 10921 -21107
rect 10977 -21047 11377 -21037
rect 10977 -21107 10987 -21047
rect 11047 -21107 11307 -21047
rect 11367 -21107 11377 -21047
rect 10977 -21217 11377 -21107
rect 11433 -21047 11833 -21037
rect 11433 -21107 11443 -21047
rect 11503 -21107 11763 -21047
rect 11823 -21107 11833 -21047
rect 11433 -21217 11833 -21107
rect 11891 -21047 12291 -21037
rect 11891 -21107 11901 -21047
rect 11961 -21107 12221 -21047
rect 12281 -21107 12291 -21047
rect 11891 -21217 12291 -21107
rect 12347 -21047 12747 -21037
rect 12347 -21107 12357 -21047
rect 12417 -21107 12677 -21047
rect 12737 -21107 12747 -21047
rect 12347 -21217 12747 -21107
rect 12803 -21047 13203 -21037
rect 12803 -21107 12813 -21047
rect 12873 -21107 13133 -21047
rect 13193 -21107 13203 -21047
rect 12803 -21217 13203 -21107
rect 13261 -21047 13661 -21037
rect 13261 -21107 13271 -21047
rect 13331 -21107 13591 -21047
rect 13651 -21107 13661 -21047
rect 13261 -21217 13661 -21107
rect 13717 -21047 14117 -21037
rect 13717 -21107 13727 -21047
rect 13787 -21107 14047 -21047
rect 14107 -21107 14117 -21047
rect 13717 -21217 14117 -21107
rect 14173 -21047 14573 -21037
rect 14173 -21107 14183 -21047
rect 14243 -21107 14503 -21047
rect 14563 -21107 14573 -21047
rect 14173 -21217 14573 -21107
rect 14631 -21047 15031 -21037
rect 14631 -21107 14641 -21047
rect 14701 -21107 14961 -21047
rect 15021 -21107 15031 -21047
rect 14631 -21217 15031 -21107
rect 15087 -21047 15487 -21037
rect 15087 -21107 15097 -21047
rect 15157 -21107 15417 -21047
rect 15477 -21107 15487 -21047
rect 15087 -21217 15487 -21107
rect 10521 -21218 15487 -21217
rect 10521 -21219 15721 -21218
rect 7307 -21289 15721 -21219
rect 7307 -21397 7707 -21289
rect 7307 -21457 7317 -21397
rect 7377 -21457 7637 -21397
rect 7697 -21457 7707 -21397
rect 7307 -21467 7707 -21457
rect 7763 -21397 8163 -21289
rect 7763 -21457 7773 -21397
rect 7833 -21457 8093 -21397
rect 8153 -21457 8163 -21397
rect 7763 -21467 8163 -21457
rect 8237 -21397 8637 -21289
rect 8237 -21457 8247 -21397
rect 8307 -21457 8567 -21397
rect 8627 -21457 8637 -21397
rect 8237 -21467 8637 -21457
rect 8693 -21397 9093 -21289
rect 8693 -21457 8703 -21397
rect 8763 -21457 9023 -21397
rect 9083 -21457 9093 -21397
rect 8693 -21467 9093 -21457
rect 9151 -21397 9551 -21289
rect 9151 -21457 9161 -21397
rect 9221 -21457 9481 -21397
rect 9541 -21457 9551 -21397
rect 9151 -21467 9551 -21457
rect 9607 -21397 10007 -21289
rect 9607 -21457 9617 -21397
rect 9677 -21457 9937 -21397
rect 9997 -21457 10007 -21397
rect 9607 -21467 10007 -21457
rect 10063 -21397 10463 -21289
rect 10063 -21457 10073 -21397
rect 10133 -21457 10393 -21397
rect 10453 -21457 10463 -21397
rect 10063 -21467 10463 -21457
rect 10521 -21397 10921 -21289
rect 10521 -21457 10531 -21397
rect 10591 -21457 10851 -21397
rect 10911 -21457 10921 -21397
rect 10521 -21467 10921 -21457
rect 10977 -21397 11377 -21289
rect 10977 -21457 10987 -21397
rect 11047 -21457 11307 -21397
rect 11367 -21457 11377 -21397
rect 10977 -21467 11377 -21457
rect 11433 -21397 11833 -21289
rect 11433 -21457 11443 -21397
rect 11503 -21457 11763 -21397
rect 11823 -21457 11833 -21397
rect 11433 -21467 11833 -21457
rect 11891 -21397 12291 -21289
rect 11891 -21457 11901 -21397
rect 11961 -21457 12221 -21397
rect 12281 -21457 12291 -21397
rect 11891 -21467 12291 -21457
rect 12347 -21397 12747 -21289
rect 12347 -21457 12357 -21397
rect 12417 -21457 12677 -21397
rect 12737 -21457 12747 -21397
rect 12347 -21467 12747 -21457
rect 12803 -21397 13203 -21289
rect 12803 -21457 12813 -21397
rect 12873 -21457 13133 -21397
rect 13193 -21457 13203 -21397
rect 12803 -21467 13203 -21457
rect 13261 -21397 13661 -21289
rect 13261 -21457 13271 -21397
rect 13331 -21457 13591 -21397
rect 13651 -21457 13661 -21397
rect 13261 -21467 13661 -21457
rect 13717 -21397 14117 -21289
rect 13717 -21457 13727 -21397
rect 13787 -21457 14047 -21397
rect 14107 -21457 14117 -21397
rect 13717 -21467 14117 -21457
rect 14173 -21397 14573 -21289
rect 14173 -21457 14183 -21397
rect 14243 -21457 14503 -21397
rect 14563 -21457 14573 -21397
rect 14173 -21467 14573 -21457
rect 14631 -21397 15031 -21289
rect 14631 -21457 14641 -21397
rect 14701 -21457 14961 -21397
rect 15021 -21457 15031 -21397
rect 14631 -21467 15031 -21457
rect 15087 -21397 15487 -21289
rect 15087 -21457 15097 -21397
rect 15157 -21457 15417 -21397
rect 15477 -21457 15487 -21397
rect 15087 -21467 15487 -21457
rect 66 -21539 80 -21467
rect 457 -21539 527 -21467
rect 913 -21539 984 -21467
rect 1371 -21539 1442 -21467
rect 1827 -21539 1898 -21467
rect 2283 -21539 2354 -21467
rect 2741 -21539 2812 -21467
rect 3197 -21539 3268 -21467
rect 3653 -21539 3724 -21467
rect 4111 -21539 4182 -21467
rect 4567 -21539 4638 -21467
rect 5023 -21539 5094 -21467
rect 5481 -21539 5552 -21467
rect 5937 -21539 6008 -21467
rect 6393 -21539 6464 -21467
rect 6851 -21539 6922 -21467
rect 7307 -21539 7378 -21467
rect 7763 -21539 7834 -21467
rect 8237 -21539 8308 -21467
rect 8693 -21539 8764 -21467
rect 9151 -21539 9222 -21467
rect 9607 -21539 9678 -21467
rect 10063 -21539 10134 -21467
rect 10521 -21539 10592 -21467
rect 10977 -21539 11048 -21467
rect 11433 -21539 11504 -21467
rect 11891 -21539 11962 -21467
rect 12347 -21539 12418 -21467
rect 12803 -21539 12874 -21467
rect 13261 -21539 13332 -21467
rect 13717 -21539 13788 -21467
rect 14173 -21539 14244 -21467
rect 14631 -21539 14702 -21467
rect 66 -21549 400 -21539
rect 0 -21609 11 -21549
rect 71 -21609 331 -21549
rect 391 -21609 400 -21549
rect 0 -21899 14 -21609
rect 66 -21899 400 -21609
rect 0 -21959 11 -21899
rect 71 -21959 331 -21899
rect 391 -21959 400 -21899
rect 0 -22041 14 -21959
rect 66 -21969 400 -21959
rect 457 -21549 857 -21539
rect 457 -21609 467 -21549
rect 527 -21609 787 -21549
rect 847 -21609 857 -21549
rect 457 -21719 857 -21609
rect 913 -21549 1313 -21539
rect 913 -21609 923 -21549
rect 983 -21609 1243 -21549
rect 1303 -21609 1313 -21549
rect 913 -21719 1313 -21609
rect 1371 -21549 1771 -21539
rect 1371 -21609 1381 -21549
rect 1441 -21609 1701 -21549
rect 1761 -21609 1771 -21549
rect 1371 -21719 1771 -21609
rect 1827 -21549 2227 -21539
rect 1827 -21609 1837 -21549
rect 1897 -21609 2157 -21549
rect 2217 -21609 2227 -21549
rect 1827 -21719 2227 -21609
rect 2283 -21549 2683 -21539
rect 2283 -21609 2293 -21549
rect 2353 -21609 2613 -21549
rect 2673 -21609 2683 -21549
rect 2283 -21719 2683 -21609
rect 457 -21720 2683 -21719
rect 2741 -21549 3141 -21539
rect 2741 -21609 2751 -21549
rect 2811 -21609 3071 -21549
rect 3131 -21609 3141 -21549
rect 2741 -21719 3141 -21609
rect 3197 -21549 3597 -21539
rect 3197 -21609 3207 -21549
rect 3267 -21609 3527 -21549
rect 3587 -21609 3597 -21549
rect 3197 -21719 3597 -21609
rect 3653 -21549 4053 -21539
rect 3653 -21609 3663 -21549
rect 3723 -21609 3983 -21549
rect 4043 -21609 4053 -21549
rect 3653 -21719 4053 -21609
rect 2741 -21720 4053 -21719
rect 457 -21790 4053 -21720
rect 457 -21899 857 -21790
rect 457 -21959 467 -21899
rect 527 -21959 787 -21899
rect 847 -21959 857 -21899
rect 457 -21969 857 -21959
rect 913 -21899 1313 -21790
rect 913 -21959 923 -21899
rect 983 -21959 1243 -21899
rect 1303 -21959 1313 -21899
rect 913 -21969 1313 -21959
rect 1371 -21899 1771 -21790
rect 1371 -21959 1381 -21899
rect 1441 -21959 1701 -21899
rect 1761 -21959 1771 -21899
rect 1371 -21969 1771 -21959
rect 1827 -21899 2227 -21790
rect 1827 -21959 1837 -21899
rect 1897 -21959 2157 -21899
rect 2217 -21959 2227 -21899
rect 1827 -21969 2227 -21959
rect 2283 -21899 2683 -21790
rect 2283 -21959 2293 -21899
rect 2353 -21959 2613 -21899
rect 2673 -21959 2683 -21899
rect 2283 -21969 2683 -21959
rect 2741 -21899 3141 -21790
rect 2741 -21959 2751 -21899
rect 2811 -21959 3071 -21899
rect 3131 -21959 3141 -21899
rect 2741 -21969 3141 -21959
rect 3197 -21899 3597 -21790
rect 3197 -21959 3207 -21899
rect 3267 -21959 3527 -21899
rect 3587 -21959 3597 -21899
rect 3197 -21969 3597 -21959
rect 3653 -21899 4053 -21790
rect 3653 -21959 3663 -21899
rect 3723 -21959 3983 -21899
rect 4043 -21959 4053 -21899
rect 3653 -21969 4053 -21959
rect 4111 -21549 4511 -21539
rect 4111 -21609 4121 -21549
rect 4181 -21609 4441 -21549
rect 4501 -21609 4511 -21549
rect 4111 -21719 4511 -21609
rect 4567 -21549 4967 -21539
rect 4567 -21609 4577 -21549
rect 4637 -21609 4897 -21549
rect 4957 -21609 4967 -21549
rect 4567 -21719 4967 -21609
rect 5023 -21549 5423 -21539
rect 5023 -21609 5033 -21549
rect 5093 -21609 5353 -21549
rect 5413 -21609 5423 -21549
rect 5023 -21719 5423 -21609
rect 5481 -21549 5881 -21539
rect 5481 -21609 5491 -21549
rect 5551 -21609 5811 -21549
rect 5871 -21609 5881 -21549
rect 5481 -21719 5881 -21609
rect 5937 -21549 6337 -21539
rect 5937 -21609 5947 -21549
rect 6007 -21609 6267 -21549
rect 6327 -21609 6337 -21549
rect 5937 -21719 6337 -21609
rect 6393 -21549 6793 -21539
rect 6393 -21609 6403 -21549
rect 6463 -21609 6723 -21549
rect 6783 -21609 6793 -21549
rect 6393 -21719 6793 -21609
rect 6851 -21549 7251 -21539
rect 6851 -21609 6861 -21549
rect 6921 -21609 7181 -21549
rect 7241 -21609 7251 -21549
rect 6851 -21719 7251 -21609
rect 4111 -21790 7251 -21719
rect 4111 -21899 4511 -21790
rect 4111 -21959 4121 -21899
rect 4181 -21959 4441 -21899
rect 4501 -21959 4511 -21899
rect 4111 -21969 4511 -21959
rect 4567 -21899 4967 -21790
rect 4567 -21959 4577 -21899
rect 4637 -21959 4897 -21899
rect 4957 -21959 4967 -21899
rect 4567 -21969 4967 -21959
rect 5023 -21899 5423 -21790
rect 5023 -21959 5033 -21899
rect 5093 -21959 5353 -21899
rect 5413 -21959 5423 -21899
rect 5023 -21969 5423 -21959
rect 5481 -21899 5881 -21790
rect 5481 -21959 5491 -21899
rect 5551 -21959 5811 -21899
rect 5871 -21959 5881 -21899
rect 5481 -21969 5881 -21959
rect 5937 -21899 6337 -21790
rect 5937 -21959 5947 -21899
rect 6007 -21959 6267 -21899
rect 6327 -21959 6337 -21899
rect 5937 -21969 6337 -21959
rect 6393 -21899 6793 -21790
rect 6393 -21959 6403 -21899
rect 6463 -21959 6723 -21899
rect 6783 -21959 6793 -21899
rect 6393 -21969 6793 -21959
rect 6851 -21899 7251 -21790
rect 6851 -21959 6861 -21899
rect 6921 -21959 7181 -21899
rect 7241 -21959 7251 -21899
rect 6851 -21969 7251 -21959
rect 7307 -21549 7707 -21539
rect 7307 -21609 7317 -21549
rect 7377 -21609 7637 -21549
rect 7697 -21609 7707 -21549
rect 7307 -21719 7707 -21609
rect 7763 -21549 8163 -21539
rect 7763 -21609 7773 -21549
rect 7833 -21609 8093 -21549
rect 8153 -21609 8163 -21549
rect 7763 -21719 8163 -21609
rect 8237 -21549 8637 -21539
rect 8237 -21609 8247 -21549
rect 8307 -21609 8567 -21549
rect 8627 -21609 8637 -21549
rect 8237 -21719 8637 -21609
rect 8693 -21549 9093 -21539
rect 8693 -21609 8703 -21549
rect 8763 -21609 9023 -21549
rect 9083 -21609 9093 -21549
rect 8693 -21719 9093 -21609
rect 9151 -21549 9551 -21539
rect 9151 -21609 9161 -21549
rect 9221 -21609 9481 -21549
rect 9541 -21609 9551 -21549
rect 9151 -21719 9551 -21609
rect 9607 -21549 10007 -21539
rect 9607 -21609 9617 -21549
rect 9677 -21609 9937 -21549
rect 9997 -21609 10007 -21549
rect 9607 -21719 10007 -21609
rect 10063 -21549 10463 -21539
rect 10063 -21609 10073 -21549
rect 10133 -21609 10393 -21549
rect 10453 -21609 10463 -21549
rect 10063 -21719 10463 -21609
rect 7307 -21720 10463 -21719
rect 10521 -21549 10921 -21539
rect 10521 -21609 10531 -21549
rect 10591 -21609 10851 -21549
rect 10911 -21609 10921 -21549
rect 10521 -21719 10921 -21609
rect 10977 -21549 11377 -21539
rect 10977 -21609 10987 -21549
rect 11047 -21609 11307 -21549
rect 11367 -21609 11377 -21549
rect 10977 -21719 11377 -21609
rect 11433 -21549 11833 -21539
rect 11433 -21609 11443 -21549
rect 11503 -21609 11763 -21549
rect 11823 -21609 11833 -21549
rect 11433 -21719 11833 -21609
rect 11891 -21549 12291 -21539
rect 11891 -21609 11901 -21549
rect 11961 -21609 12221 -21549
rect 12281 -21609 12291 -21549
rect 11891 -21719 12291 -21609
rect 12347 -21549 12747 -21539
rect 12347 -21609 12357 -21549
rect 12417 -21609 12677 -21549
rect 12737 -21609 12747 -21549
rect 12347 -21719 12747 -21609
rect 12803 -21549 13203 -21539
rect 12803 -21609 12813 -21549
rect 12873 -21609 13133 -21549
rect 13193 -21609 13203 -21549
rect 12803 -21719 13203 -21609
rect 13261 -21549 13661 -21539
rect 13261 -21609 13271 -21549
rect 13331 -21609 13591 -21549
rect 13651 -21609 13661 -21549
rect 13261 -21719 13661 -21609
rect 13717 -21549 14117 -21539
rect 13717 -21609 13727 -21549
rect 13787 -21609 14047 -21549
rect 14107 -21609 14117 -21549
rect 13717 -21719 14117 -21609
rect 14173 -21549 14573 -21539
rect 14173 -21609 14183 -21549
rect 14243 -21609 14503 -21549
rect 14563 -21609 14573 -21549
rect 14173 -21719 14573 -21609
rect 14631 -21549 15031 -21539
rect 14631 -21609 14641 -21549
rect 14701 -21609 14961 -21549
rect 15021 -21609 15031 -21549
rect 14631 -21719 15031 -21609
rect 15087 -21549 15487 -21539
rect 15087 -21609 15097 -21549
rect 15157 -21609 15417 -21549
rect 15477 -21609 15487 -21549
rect 15087 -21719 15487 -21609
rect 10521 -21720 15487 -21719
rect 7307 -21790 15487 -21720
rect 7307 -21899 7707 -21790
rect 7307 -21959 7317 -21899
rect 7377 -21959 7637 -21899
rect 7697 -21959 7707 -21899
rect 7307 -21969 7707 -21959
rect 7763 -21899 8163 -21790
rect 7763 -21959 7773 -21899
rect 7833 -21959 8093 -21899
rect 8153 -21959 8163 -21899
rect 7763 -21969 8163 -21959
rect 8237 -21899 8637 -21790
rect 8237 -21959 8247 -21899
rect 8307 -21959 8567 -21899
rect 8627 -21959 8637 -21899
rect 8237 -21969 8637 -21959
rect 8693 -21899 9093 -21790
rect 8693 -21959 8703 -21899
rect 8763 -21959 9023 -21899
rect 9083 -21959 9093 -21899
rect 8693 -21969 9093 -21959
rect 9151 -21899 9551 -21790
rect 9151 -21959 9161 -21899
rect 9221 -21959 9481 -21899
rect 9541 -21959 9551 -21899
rect 9151 -21969 9551 -21959
rect 9607 -21899 10007 -21790
rect 9607 -21959 9617 -21899
rect 9677 -21959 9937 -21899
rect 9997 -21959 10007 -21899
rect 9607 -21969 10007 -21959
rect 10063 -21899 10463 -21790
rect 10063 -21959 10073 -21899
rect 10133 -21959 10393 -21899
rect 10453 -21959 10463 -21899
rect 10063 -21969 10463 -21959
rect 10521 -21899 10921 -21790
rect 10521 -21959 10531 -21899
rect 10591 -21959 10851 -21899
rect 10911 -21959 10921 -21899
rect 10521 -21969 10921 -21959
rect 10977 -21899 11377 -21790
rect 10977 -21959 10987 -21899
rect 11047 -21959 11307 -21899
rect 11367 -21959 11377 -21899
rect 10977 -21969 11377 -21959
rect 11433 -21899 11833 -21790
rect 11433 -21959 11443 -21899
rect 11503 -21959 11763 -21899
rect 11823 -21959 11833 -21899
rect 11433 -21969 11833 -21959
rect 11891 -21899 12291 -21790
rect 11891 -21959 11901 -21899
rect 11961 -21959 12221 -21899
rect 12281 -21959 12291 -21899
rect 11891 -21969 12291 -21959
rect 12347 -21899 12747 -21790
rect 12347 -21959 12357 -21899
rect 12417 -21959 12677 -21899
rect 12737 -21959 12747 -21899
rect 12347 -21969 12747 -21959
rect 12803 -21899 13203 -21790
rect 12803 -21959 12813 -21899
rect 12873 -21959 13133 -21899
rect 13193 -21959 13203 -21899
rect 12803 -21969 13203 -21959
rect 13261 -21899 13661 -21790
rect 13261 -21959 13271 -21899
rect 13331 -21959 13591 -21899
rect 13651 -21959 13661 -21899
rect 13261 -21969 13661 -21959
rect 13717 -21899 14117 -21790
rect 13717 -21959 13727 -21899
rect 13787 -21959 14047 -21899
rect 14107 -21959 14117 -21899
rect 13717 -21969 14117 -21959
rect 14173 -21899 14573 -21790
rect 14173 -21959 14183 -21899
rect 14243 -21959 14503 -21899
rect 14563 -21959 14573 -21899
rect 14173 -21969 14573 -21959
rect 14631 -21899 15031 -21790
rect 14631 -21959 14641 -21899
rect 14701 -21959 14961 -21899
rect 15021 -21959 15031 -21899
rect 14631 -21969 15031 -21959
rect 15087 -21899 15487 -21790
rect 15087 -21959 15097 -21899
rect 15157 -21959 15417 -21899
rect 15477 -21959 15487 -21899
rect 15087 -21969 15487 -21959
rect 66 -22031 80 -21969
rect 457 -22031 528 -21969
rect 913 -22031 984 -21969
rect 1371 -22031 1442 -21969
rect 1827 -22031 1898 -21969
rect 2283 -22031 2354 -21969
rect 2741 -22031 2811 -21969
rect 3197 -22031 3267 -21969
rect 3653 -22031 3723 -21969
rect 4111 -22031 4181 -21969
rect 4567 -22031 4637 -21969
rect 5023 -22031 5093 -21969
rect 5481 -22031 5551 -21969
rect 5937 -22031 6007 -21969
rect 6393 -22031 6463 -21969
rect 6851 -22031 6921 -21969
rect 7307 -22031 7377 -21969
rect 7763 -22031 7833 -21969
rect 8237 -22031 8307 -21969
rect 8693 -22031 8763 -21969
rect 9151 -22031 9221 -21969
rect 9607 -22031 9677 -21969
rect 10063 -22031 10133 -21969
rect 10521 -22031 10591 -21969
rect 10977 -22031 11047 -21969
rect 11433 -22031 11503 -21969
rect 11891 -22031 11961 -21969
rect 12347 -22031 12417 -21969
rect 12803 -22031 12873 -21969
rect 13261 -22031 13331 -21969
rect 13717 -22031 13787 -21969
rect 14173 -22031 14243 -21969
rect 14631 -22031 14701 -21969
rect 66 -22041 400 -22031
rect 0 -22101 11 -22041
rect 71 -22101 331 -22041
rect 391 -22101 400 -22041
rect 0 -22391 14 -22101
rect 66 -22391 400 -22101
rect 0 -22451 11 -22391
rect 71 -22451 331 -22391
rect 391 -22451 400 -22391
rect 0 -22528 14 -22451
rect 66 -22461 400 -22451
rect 457 -22041 857 -22031
rect 457 -22101 467 -22041
rect 527 -22101 787 -22041
rect 847 -22101 857 -22041
rect 457 -22211 857 -22101
rect 913 -22041 1313 -22031
rect 913 -22101 923 -22041
rect 983 -22101 1243 -22041
rect 1303 -22101 1313 -22041
rect 913 -22211 1313 -22101
rect 1371 -22041 1771 -22031
rect 1371 -22101 1381 -22041
rect 1441 -22101 1701 -22041
rect 1761 -22101 1771 -22041
rect 1371 -22211 1771 -22101
rect 1827 -22041 2227 -22031
rect 1827 -22101 1837 -22041
rect 1897 -22101 2157 -22041
rect 2217 -22101 2227 -22041
rect 1827 -22211 2227 -22101
rect 2283 -22041 2683 -22031
rect 2283 -22101 2293 -22041
rect 2353 -22101 2613 -22041
rect 2673 -22101 2683 -22041
rect 2283 -22211 2683 -22101
rect 2741 -22041 3141 -22031
rect 2741 -22101 2751 -22041
rect 2811 -22101 3071 -22041
rect 3131 -22101 3141 -22041
rect 2741 -22211 3141 -22101
rect 3197 -22041 3597 -22031
rect 3197 -22101 3207 -22041
rect 3267 -22101 3527 -22041
rect 3587 -22101 3597 -22041
rect 3197 -22211 3597 -22101
rect 3653 -22041 4053 -22031
rect 3653 -22101 3663 -22041
rect 3723 -22101 3983 -22041
rect 4043 -22101 4053 -22041
rect 3653 -22211 4053 -22101
rect 457 -22281 4053 -22211
rect 457 -22391 857 -22281
rect 457 -22451 467 -22391
rect 527 -22451 787 -22391
rect 847 -22451 857 -22391
rect 457 -22461 857 -22451
rect 913 -22391 1313 -22281
rect 913 -22451 923 -22391
rect 983 -22451 1243 -22391
rect 1303 -22451 1313 -22391
rect 913 -22461 1313 -22451
rect 1371 -22391 1771 -22281
rect 1371 -22451 1381 -22391
rect 1441 -22451 1701 -22391
rect 1761 -22451 1771 -22391
rect 1371 -22461 1771 -22451
rect 1827 -22391 2227 -22281
rect 1827 -22451 1837 -22391
rect 1897 -22451 2157 -22391
rect 2217 -22451 2227 -22391
rect 1827 -22461 2227 -22451
rect 2283 -22391 2683 -22281
rect 2283 -22451 2293 -22391
rect 2353 -22451 2613 -22391
rect 2673 -22451 2683 -22391
rect 2283 -22461 2683 -22451
rect 2741 -22391 3141 -22281
rect 2741 -22451 2751 -22391
rect 2811 -22451 3071 -22391
rect 3131 -22451 3141 -22391
rect 2741 -22461 3141 -22451
rect 3197 -22391 3597 -22281
rect 3197 -22451 3207 -22391
rect 3267 -22451 3527 -22391
rect 3587 -22451 3597 -22391
rect 3197 -22461 3597 -22451
rect 3653 -22391 4053 -22281
rect 3653 -22451 3663 -22391
rect 3723 -22451 3983 -22391
rect 4043 -22451 4053 -22391
rect 3653 -22461 4053 -22451
rect 4111 -22041 4511 -22031
rect 4111 -22101 4121 -22041
rect 4181 -22101 4441 -22041
rect 4501 -22101 4511 -22041
rect 4111 -22211 4511 -22101
rect 4567 -22041 4967 -22031
rect 4567 -22101 4577 -22041
rect 4637 -22101 4897 -22041
rect 4957 -22101 4967 -22041
rect 4567 -22211 4967 -22101
rect 5023 -22041 5423 -22031
rect 5023 -22101 5033 -22041
rect 5093 -22101 5353 -22041
rect 5413 -22101 5423 -22041
rect 5023 -22211 5423 -22101
rect 5481 -22041 5881 -22031
rect 5481 -22101 5491 -22041
rect 5551 -22101 5811 -22041
rect 5871 -22101 5881 -22041
rect 5481 -22211 5881 -22101
rect 5937 -22041 6337 -22031
rect 5937 -22101 5947 -22041
rect 6007 -22101 6267 -22041
rect 6327 -22101 6337 -22041
rect 5937 -22211 6337 -22101
rect 6393 -22041 6793 -22031
rect 6393 -22101 6403 -22041
rect 6463 -22101 6723 -22041
rect 6783 -22101 6793 -22041
rect 6393 -22211 6793 -22101
rect 6851 -22041 7251 -22031
rect 6851 -22101 6861 -22041
rect 6921 -22101 7181 -22041
rect 7241 -22101 7251 -22041
rect 6851 -22211 7251 -22101
rect 4111 -22281 7251 -22211
rect 4111 -22391 4511 -22281
rect 4111 -22451 4121 -22391
rect 4181 -22451 4441 -22391
rect 4501 -22451 4511 -22391
rect 4111 -22461 4511 -22451
rect 4567 -22391 4967 -22281
rect 4567 -22451 4577 -22391
rect 4637 -22451 4897 -22391
rect 4957 -22451 4967 -22391
rect 4567 -22461 4967 -22451
rect 5023 -22391 5423 -22281
rect 5023 -22451 5033 -22391
rect 5093 -22451 5353 -22391
rect 5413 -22451 5423 -22391
rect 5023 -22461 5423 -22451
rect 5481 -22391 5881 -22281
rect 5481 -22451 5491 -22391
rect 5551 -22451 5811 -22391
rect 5871 -22451 5881 -22391
rect 5481 -22461 5881 -22451
rect 5937 -22391 6337 -22281
rect 5937 -22451 5947 -22391
rect 6007 -22451 6267 -22391
rect 6327 -22451 6337 -22391
rect 5937 -22461 6337 -22451
rect 6393 -22391 6793 -22281
rect 6393 -22451 6403 -22391
rect 6463 -22451 6723 -22391
rect 6783 -22451 6793 -22391
rect 6393 -22461 6793 -22451
rect 6851 -22391 7251 -22281
rect 6851 -22451 6861 -22391
rect 6921 -22451 7181 -22391
rect 7241 -22451 7251 -22391
rect 6851 -22461 7251 -22451
rect 7307 -22041 7707 -22031
rect 7307 -22101 7317 -22041
rect 7377 -22101 7637 -22041
rect 7697 -22101 7707 -22041
rect 7307 -22211 7707 -22101
rect 7763 -22041 8163 -22031
rect 7763 -22101 7773 -22041
rect 7833 -22101 8093 -22041
rect 8153 -22101 8163 -22041
rect 7763 -22211 8163 -22101
rect 8237 -22041 8637 -22031
rect 8237 -22101 8247 -22041
rect 8307 -22101 8567 -22041
rect 8627 -22101 8637 -22041
rect 8237 -22211 8637 -22101
rect 8693 -22041 9093 -22031
rect 8693 -22101 8703 -22041
rect 8763 -22101 9023 -22041
rect 9083 -22101 9093 -22041
rect 8693 -22211 9093 -22101
rect 9151 -22041 9551 -22031
rect 9151 -22101 9161 -22041
rect 9221 -22101 9481 -22041
rect 9541 -22101 9551 -22041
rect 9151 -22211 9551 -22101
rect 9607 -22041 10007 -22031
rect 9607 -22101 9617 -22041
rect 9677 -22101 9937 -22041
rect 9997 -22101 10007 -22041
rect 9607 -22211 10007 -22101
rect 10063 -22041 10463 -22031
rect 10063 -22101 10073 -22041
rect 10133 -22101 10393 -22041
rect 10453 -22101 10463 -22041
rect 10063 -22211 10463 -22101
rect 10521 -22041 10921 -22031
rect 10521 -22101 10531 -22041
rect 10591 -22101 10851 -22041
rect 10911 -22101 10921 -22041
rect 10521 -22211 10921 -22101
rect 10977 -22041 11377 -22031
rect 10977 -22101 10987 -22041
rect 11047 -22101 11307 -22041
rect 11367 -22101 11377 -22041
rect 10977 -22211 11377 -22101
rect 11433 -22041 11833 -22031
rect 11433 -22101 11443 -22041
rect 11503 -22101 11763 -22041
rect 11823 -22101 11833 -22041
rect 11433 -22211 11833 -22101
rect 11891 -22041 12291 -22031
rect 11891 -22101 11901 -22041
rect 11961 -22101 12221 -22041
rect 12281 -22101 12291 -22041
rect 11891 -22211 12291 -22101
rect 12347 -22041 12747 -22031
rect 12347 -22101 12357 -22041
rect 12417 -22101 12677 -22041
rect 12737 -22101 12747 -22041
rect 12347 -22211 12747 -22101
rect 12803 -22041 13203 -22031
rect 12803 -22101 12813 -22041
rect 12873 -22101 13133 -22041
rect 13193 -22101 13203 -22041
rect 12803 -22211 13203 -22101
rect 13261 -22041 13661 -22031
rect 13261 -22101 13271 -22041
rect 13331 -22101 13591 -22041
rect 13651 -22101 13661 -22041
rect 13261 -22211 13661 -22101
rect 13717 -22041 14117 -22031
rect 13717 -22101 13727 -22041
rect 13787 -22101 14047 -22041
rect 14107 -22101 14117 -22041
rect 13717 -22211 14117 -22101
rect 14173 -22041 14573 -22031
rect 14173 -22101 14183 -22041
rect 14243 -22101 14503 -22041
rect 14563 -22101 14573 -22041
rect 14173 -22211 14573 -22101
rect 14631 -22041 15031 -22031
rect 14631 -22101 14641 -22041
rect 14701 -22101 14961 -22041
rect 15021 -22101 15031 -22041
rect 14631 -22211 15031 -22101
rect 15087 -22041 15487 -22031
rect 15087 -22101 15097 -22041
rect 15157 -22101 15417 -22041
rect 15477 -22101 15487 -22041
rect 15087 -22211 15487 -22101
rect 7307 -22281 15487 -22211
rect 7307 -22391 7707 -22281
rect 7307 -22451 7317 -22391
rect 7377 -22451 7637 -22391
rect 7697 -22451 7707 -22391
rect 7307 -22461 7707 -22451
rect 7763 -22391 8163 -22281
rect 7763 -22451 7773 -22391
rect 7833 -22451 8093 -22391
rect 8153 -22451 8163 -22391
rect 7763 -22461 8163 -22451
rect 8237 -22391 8637 -22281
rect 8237 -22451 8247 -22391
rect 8307 -22451 8567 -22391
rect 8627 -22451 8637 -22391
rect 8237 -22461 8637 -22451
rect 8693 -22391 9093 -22281
rect 8693 -22451 8703 -22391
rect 8763 -22451 9023 -22391
rect 9083 -22451 9093 -22391
rect 8693 -22461 9093 -22451
rect 9151 -22391 9551 -22281
rect 9151 -22451 9161 -22391
rect 9221 -22451 9481 -22391
rect 9541 -22451 9551 -22391
rect 9151 -22461 9551 -22451
rect 9607 -22391 10007 -22281
rect 9607 -22451 9617 -22391
rect 9677 -22451 9937 -22391
rect 9997 -22451 10007 -22391
rect 9607 -22461 10007 -22451
rect 10063 -22391 10463 -22281
rect 10063 -22451 10073 -22391
rect 10133 -22451 10393 -22391
rect 10453 -22451 10463 -22391
rect 10063 -22461 10463 -22451
rect 10521 -22391 10921 -22281
rect 10521 -22451 10531 -22391
rect 10591 -22451 10851 -22391
rect 10911 -22451 10921 -22391
rect 10521 -22461 10921 -22451
rect 10977 -22391 11377 -22281
rect 10977 -22451 10987 -22391
rect 11047 -22451 11307 -22391
rect 11367 -22451 11377 -22391
rect 10977 -22461 11377 -22451
rect 11433 -22391 11833 -22281
rect 11433 -22451 11443 -22391
rect 11503 -22451 11763 -22391
rect 11823 -22451 11833 -22391
rect 11433 -22461 11833 -22451
rect 11891 -22391 12291 -22281
rect 11891 -22451 11901 -22391
rect 11961 -22451 12221 -22391
rect 12281 -22451 12291 -22391
rect 11891 -22461 12291 -22451
rect 12347 -22391 12747 -22281
rect 12347 -22451 12357 -22391
rect 12417 -22451 12677 -22391
rect 12737 -22451 12747 -22391
rect 12347 -22461 12747 -22451
rect 12803 -22391 13203 -22281
rect 12803 -22451 12813 -22391
rect 12873 -22451 13133 -22391
rect 13193 -22451 13203 -22391
rect 12803 -22461 13203 -22451
rect 13261 -22391 13661 -22281
rect 13261 -22451 13271 -22391
rect 13331 -22451 13591 -22391
rect 13651 -22451 13661 -22391
rect 13261 -22461 13661 -22451
rect 13717 -22391 14117 -22281
rect 13717 -22451 13727 -22391
rect 13787 -22451 14047 -22391
rect 14107 -22451 14117 -22391
rect 13717 -22461 14117 -22451
rect 14173 -22391 14573 -22281
rect 14173 -22451 14183 -22391
rect 14243 -22451 14503 -22391
rect 14563 -22451 14573 -22391
rect 14173 -22461 14573 -22451
rect 14631 -22391 15031 -22281
rect 14631 -22451 14641 -22391
rect 14701 -22451 14961 -22391
rect 15021 -22451 15031 -22391
rect 14631 -22461 15031 -22451
rect 15087 -22391 15487 -22281
rect 15087 -22451 15097 -22391
rect 15157 -22451 15417 -22391
rect 15477 -22451 15487 -22391
rect 15087 -22461 15487 -22451
rect 66 -22518 80 -22461
rect 457 -22518 529 -22461
rect 913 -22518 985 -22461
rect 1371 -22518 1443 -22461
rect 1827 -22518 1899 -22461
rect 2283 -22518 2355 -22461
rect 2741 -22518 2813 -22461
rect 3197 -22518 3269 -22461
rect 3653 -22518 3725 -22461
rect 4111 -22518 4183 -22461
rect 4567 -22518 4639 -22461
rect 5023 -22518 5095 -22461
rect 5481 -22518 5553 -22461
rect 5937 -22518 6007 -22461
rect 6393 -22518 6463 -22461
rect 6851 -22518 6921 -22461
rect 7307 -22518 7380 -22461
rect 7763 -22518 7836 -22461
rect 8237 -22518 8310 -22461
rect 8693 -22518 8766 -22461
rect 9151 -22518 9224 -22461
rect 9607 -22518 9680 -22461
rect 10063 -22518 10136 -22461
rect 10521 -22518 10594 -22461
rect 10977 -22518 11050 -22461
rect 11433 -22518 11506 -22461
rect 11891 -22518 11964 -22461
rect 12347 -22518 12420 -22461
rect 12803 -22518 12876 -22461
rect 13261 -22518 13334 -22461
rect 13717 -22518 13790 -22461
rect 14173 -22518 14246 -22461
rect 14631 -22518 14704 -22461
rect 66 -22528 400 -22518
rect 0 -22588 11 -22528
rect 71 -22588 331 -22528
rect 391 -22588 400 -22528
rect 0 -22878 14 -22588
rect 66 -22878 400 -22588
rect 0 -22938 11 -22878
rect 71 -22938 331 -22878
rect 391 -22938 400 -22878
rect 0 -23030 14 -22938
rect 66 -22948 400 -22938
rect 457 -22528 857 -22518
rect 457 -22588 467 -22528
rect 527 -22588 787 -22528
rect 847 -22588 857 -22528
rect 457 -22698 857 -22588
rect 913 -22528 1313 -22518
rect 913 -22588 923 -22528
rect 983 -22588 1243 -22528
rect 1303 -22588 1313 -22528
rect 913 -22698 1313 -22588
rect 1371 -22528 1771 -22518
rect 1371 -22588 1381 -22528
rect 1441 -22588 1701 -22528
rect 1761 -22588 1771 -22528
rect 1371 -22698 1771 -22588
rect 1827 -22528 2227 -22518
rect 1827 -22588 1837 -22528
rect 1897 -22588 2157 -22528
rect 2217 -22588 2227 -22528
rect 1827 -22698 2227 -22588
rect 2283 -22528 2683 -22518
rect 2283 -22588 2293 -22528
rect 2353 -22588 2613 -22528
rect 2673 -22588 2683 -22528
rect 2283 -22698 2683 -22588
rect 457 -22699 2683 -22698
rect 2741 -22528 3141 -22518
rect 2741 -22588 2751 -22528
rect 2811 -22588 3071 -22528
rect 3131 -22588 3141 -22528
rect 2741 -22698 3141 -22588
rect 3197 -22528 3597 -22518
rect 3197 -22588 3207 -22528
rect 3267 -22588 3527 -22528
rect 3587 -22588 3597 -22528
rect 3197 -22698 3597 -22588
rect 3653 -22528 4053 -22518
rect 3653 -22588 3663 -22528
rect 3723 -22588 3983 -22528
rect 4043 -22588 4053 -22528
rect 3653 -22698 4053 -22588
rect 2741 -22699 4053 -22698
rect 457 -22769 4053 -22699
rect 457 -22878 857 -22769
rect 457 -22938 467 -22878
rect 527 -22938 787 -22878
rect 847 -22938 857 -22878
rect 457 -22948 857 -22938
rect 913 -22878 1313 -22769
rect 913 -22938 923 -22878
rect 983 -22938 1243 -22878
rect 1303 -22938 1313 -22878
rect 913 -22948 1313 -22938
rect 1371 -22878 1771 -22769
rect 1371 -22938 1381 -22878
rect 1441 -22938 1701 -22878
rect 1761 -22938 1771 -22878
rect 1371 -22948 1771 -22938
rect 1827 -22878 2227 -22769
rect 1827 -22938 1837 -22878
rect 1897 -22938 2157 -22878
rect 2217 -22938 2227 -22878
rect 1827 -22948 2227 -22938
rect 2283 -22878 2683 -22769
rect 2283 -22938 2293 -22878
rect 2353 -22938 2613 -22878
rect 2673 -22938 2683 -22878
rect 2283 -22948 2683 -22938
rect 2741 -22878 3141 -22769
rect 2741 -22938 2751 -22878
rect 2811 -22938 3071 -22878
rect 3131 -22938 3141 -22878
rect 2741 -22948 3141 -22938
rect 3197 -22878 3597 -22769
rect 3197 -22938 3207 -22878
rect 3267 -22938 3527 -22878
rect 3587 -22938 3597 -22878
rect 3197 -22948 3597 -22938
rect 3653 -22878 4053 -22769
rect 3653 -22938 3663 -22878
rect 3723 -22938 3983 -22878
rect 4043 -22938 4053 -22878
rect 3653 -22948 4053 -22938
rect 4111 -22528 4511 -22518
rect 4111 -22588 4121 -22528
rect 4181 -22588 4441 -22528
rect 4501 -22588 4511 -22528
rect 4111 -22698 4511 -22588
rect 4567 -22528 4967 -22518
rect 4567 -22588 4577 -22528
rect 4637 -22588 4897 -22528
rect 4957 -22588 4967 -22528
rect 4567 -22698 4967 -22588
rect 5023 -22528 5423 -22518
rect 5023 -22588 5033 -22528
rect 5093 -22588 5353 -22528
rect 5413 -22588 5423 -22528
rect 5023 -22698 5423 -22588
rect 5481 -22528 5881 -22518
rect 5481 -22588 5491 -22528
rect 5551 -22588 5811 -22528
rect 5871 -22588 5881 -22528
rect 5481 -22698 5881 -22588
rect 5937 -22528 6337 -22518
rect 5937 -22588 5947 -22528
rect 6007 -22588 6267 -22528
rect 6327 -22588 6337 -22528
rect 5937 -22698 6337 -22588
rect 6393 -22528 6793 -22518
rect 6393 -22588 6403 -22528
rect 6463 -22588 6723 -22528
rect 6783 -22588 6793 -22528
rect 6393 -22698 6793 -22588
rect 6851 -22528 7251 -22518
rect 6851 -22588 6861 -22528
rect 6921 -22588 7181 -22528
rect 7241 -22588 7251 -22528
rect 6851 -22698 7251 -22588
rect 4111 -22769 7251 -22698
rect 4111 -22878 4511 -22769
rect 4111 -22938 4121 -22878
rect 4181 -22938 4441 -22878
rect 4501 -22938 4511 -22878
rect 4111 -22948 4511 -22938
rect 4567 -22878 4967 -22769
rect 4567 -22938 4577 -22878
rect 4637 -22938 4897 -22878
rect 4957 -22938 4967 -22878
rect 4567 -22948 4967 -22938
rect 5023 -22878 5423 -22769
rect 5023 -22938 5033 -22878
rect 5093 -22938 5353 -22878
rect 5413 -22938 5423 -22878
rect 5023 -22948 5423 -22938
rect 5481 -22878 5881 -22769
rect 5481 -22938 5491 -22878
rect 5551 -22938 5811 -22878
rect 5871 -22938 5881 -22878
rect 5481 -22948 5881 -22938
rect 5937 -22878 6337 -22769
rect 5937 -22938 5947 -22878
rect 6007 -22938 6267 -22878
rect 6327 -22938 6337 -22878
rect 5937 -22948 6337 -22938
rect 6393 -22878 6793 -22769
rect 6393 -22938 6403 -22878
rect 6463 -22938 6723 -22878
rect 6783 -22938 6793 -22878
rect 6393 -22948 6793 -22938
rect 6851 -22878 7251 -22769
rect 6851 -22938 6861 -22878
rect 6921 -22938 7181 -22878
rect 7241 -22938 7251 -22878
rect 6851 -22948 7251 -22938
rect 7307 -22528 7707 -22518
rect 7307 -22588 7317 -22528
rect 7377 -22588 7637 -22528
rect 7697 -22588 7707 -22528
rect 7307 -22698 7707 -22588
rect 7763 -22528 8163 -22518
rect 7763 -22588 7773 -22528
rect 7833 -22588 8093 -22528
rect 8153 -22588 8163 -22528
rect 7763 -22698 8163 -22588
rect 8237 -22528 8637 -22518
rect 8237 -22588 8247 -22528
rect 8307 -22588 8567 -22528
rect 8627 -22588 8637 -22528
rect 8237 -22698 8637 -22588
rect 8693 -22528 9093 -22518
rect 8693 -22588 8703 -22528
rect 8763 -22588 9023 -22528
rect 9083 -22588 9093 -22528
rect 8693 -22698 9093 -22588
rect 9151 -22528 9551 -22518
rect 9151 -22588 9161 -22528
rect 9221 -22588 9481 -22528
rect 9541 -22588 9551 -22528
rect 9151 -22698 9551 -22588
rect 9607 -22528 10007 -22518
rect 9607 -22588 9617 -22528
rect 9677 -22588 9937 -22528
rect 9997 -22588 10007 -22528
rect 9607 -22698 10007 -22588
rect 10063 -22528 10463 -22518
rect 10063 -22588 10073 -22528
rect 10133 -22588 10393 -22528
rect 10453 -22588 10463 -22528
rect 10063 -22698 10463 -22588
rect 7307 -22699 10463 -22698
rect 10521 -22528 10921 -22518
rect 10521 -22588 10531 -22528
rect 10591 -22588 10851 -22528
rect 10911 -22588 10921 -22528
rect 10521 -22698 10921 -22588
rect 10977 -22528 11377 -22518
rect 10977 -22588 10987 -22528
rect 11047 -22588 11307 -22528
rect 11367 -22588 11377 -22528
rect 10977 -22698 11377 -22588
rect 11433 -22528 11833 -22518
rect 11433 -22588 11443 -22528
rect 11503 -22588 11763 -22528
rect 11823 -22588 11833 -22528
rect 11433 -22698 11833 -22588
rect 11891 -22528 12291 -22518
rect 11891 -22588 11901 -22528
rect 11961 -22588 12221 -22528
rect 12281 -22588 12291 -22528
rect 11891 -22698 12291 -22588
rect 12347 -22528 12747 -22518
rect 12347 -22588 12357 -22528
rect 12417 -22588 12677 -22528
rect 12737 -22588 12747 -22528
rect 12347 -22698 12747 -22588
rect 12803 -22528 13203 -22518
rect 12803 -22588 12813 -22528
rect 12873 -22588 13133 -22528
rect 13193 -22588 13203 -22528
rect 12803 -22698 13203 -22588
rect 13261 -22528 13661 -22518
rect 13261 -22588 13271 -22528
rect 13331 -22588 13591 -22528
rect 13651 -22588 13661 -22528
rect 13261 -22698 13661 -22588
rect 13717 -22528 14117 -22518
rect 13717 -22588 13727 -22528
rect 13787 -22588 14047 -22528
rect 14107 -22588 14117 -22528
rect 13717 -22698 14117 -22588
rect 14173 -22528 14573 -22518
rect 14173 -22588 14183 -22528
rect 14243 -22588 14503 -22528
rect 14563 -22588 14573 -22528
rect 14173 -22698 14573 -22588
rect 14631 -22528 15031 -22518
rect 14631 -22588 14641 -22528
rect 14701 -22588 14961 -22528
rect 15021 -22588 15031 -22528
rect 14631 -22698 15031 -22588
rect 15087 -22528 15487 -22518
rect 15087 -22588 15097 -22528
rect 15157 -22588 15417 -22528
rect 15477 -22588 15487 -22528
rect 15087 -22698 15487 -22588
rect 10521 -22699 15487 -22698
rect 7307 -22769 15487 -22699
rect 7307 -22878 7707 -22769
rect 7307 -22938 7317 -22878
rect 7377 -22938 7637 -22878
rect 7697 -22938 7707 -22878
rect 7307 -22948 7707 -22938
rect 7763 -22878 8163 -22769
rect 7763 -22938 7773 -22878
rect 7833 -22938 8093 -22878
rect 8153 -22938 8163 -22878
rect 7763 -22948 8163 -22938
rect 8237 -22878 8637 -22769
rect 8237 -22938 8247 -22878
rect 8307 -22938 8567 -22878
rect 8627 -22938 8637 -22878
rect 8237 -22948 8637 -22938
rect 8693 -22878 9093 -22769
rect 8693 -22938 8703 -22878
rect 8763 -22938 9023 -22878
rect 9083 -22938 9093 -22878
rect 8693 -22948 9093 -22938
rect 9151 -22878 9551 -22769
rect 9151 -22938 9161 -22878
rect 9221 -22938 9481 -22878
rect 9541 -22938 9551 -22878
rect 9151 -22948 9551 -22938
rect 9607 -22878 10007 -22769
rect 9607 -22938 9617 -22878
rect 9677 -22938 9937 -22878
rect 9997 -22938 10007 -22878
rect 9607 -22948 10007 -22938
rect 10063 -22878 10463 -22769
rect 10063 -22938 10073 -22878
rect 10133 -22938 10393 -22878
rect 10453 -22938 10463 -22878
rect 10063 -22948 10463 -22938
rect 10521 -22878 10921 -22769
rect 10521 -22938 10531 -22878
rect 10591 -22938 10851 -22878
rect 10911 -22938 10921 -22878
rect 10521 -22948 10921 -22938
rect 10977 -22878 11377 -22769
rect 10977 -22938 10987 -22878
rect 11047 -22938 11307 -22878
rect 11367 -22938 11377 -22878
rect 10977 -22948 11377 -22938
rect 11433 -22878 11833 -22769
rect 11433 -22938 11443 -22878
rect 11503 -22938 11763 -22878
rect 11823 -22938 11833 -22878
rect 11433 -22948 11833 -22938
rect 11891 -22878 12291 -22769
rect 11891 -22938 11901 -22878
rect 11961 -22938 12221 -22878
rect 12281 -22938 12291 -22878
rect 11891 -22948 12291 -22938
rect 12347 -22878 12747 -22769
rect 12347 -22938 12357 -22878
rect 12417 -22938 12677 -22878
rect 12737 -22938 12747 -22878
rect 12347 -22948 12747 -22938
rect 12803 -22878 13203 -22769
rect 12803 -22938 12813 -22878
rect 12873 -22938 13133 -22878
rect 13193 -22938 13203 -22878
rect 12803 -22948 13203 -22938
rect 13261 -22878 13661 -22769
rect 13261 -22938 13271 -22878
rect 13331 -22938 13591 -22878
rect 13651 -22938 13661 -22878
rect 13261 -22948 13661 -22938
rect 13717 -22878 14117 -22769
rect 13717 -22938 13727 -22878
rect 13787 -22938 14047 -22878
rect 14107 -22938 14117 -22878
rect 13717 -22948 14117 -22938
rect 14173 -22878 14573 -22769
rect 14173 -22938 14183 -22878
rect 14243 -22938 14503 -22878
rect 14563 -22938 14573 -22878
rect 14173 -22948 14573 -22938
rect 14631 -22878 15031 -22769
rect 14631 -22938 14641 -22878
rect 14701 -22938 14961 -22878
rect 15021 -22938 15031 -22878
rect 14631 -22948 15031 -22938
rect 15087 -22878 15487 -22769
rect 15087 -22938 15097 -22878
rect 15157 -22938 15417 -22878
rect 15477 -22938 15487 -22878
rect 15087 -22948 15487 -22938
rect 66 -23020 80 -22948
rect 457 -23020 527 -22948
rect 913 -23020 984 -22948
rect 1371 -23020 1442 -22948
rect 1827 -23020 1898 -22948
rect 2283 -23020 2354 -22948
rect 2741 -23020 2812 -22948
rect 3197 -23020 3268 -22948
rect 3653 -23020 3724 -22948
rect 4111 -23020 4182 -22948
rect 4567 -23020 4638 -22948
rect 5023 -23020 5094 -22948
rect 5481 -23020 5552 -22948
rect 5937 -23020 6008 -22948
rect 6393 -23020 6464 -22948
rect 6851 -23020 6922 -22948
rect 7307 -23020 7378 -22948
rect 7763 -23020 7834 -22948
rect 8237 -23020 8308 -22948
rect 8693 -23020 8764 -22948
rect 9151 -23020 9222 -22948
rect 9607 -23020 9678 -22948
rect 10063 -23020 10134 -22948
rect 10521 -23020 10592 -22948
rect 10977 -23020 11048 -22948
rect 11433 -23020 11504 -22948
rect 11891 -23020 11962 -22948
rect 12347 -23020 12418 -22948
rect 12803 -23020 12874 -22948
rect 13261 -23020 13332 -22948
rect 13717 -23020 13788 -22948
rect 14173 -23020 14244 -22948
rect 14631 -23020 14702 -22948
rect 66 -23030 400 -23020
rect 0 -23090 11 -23030
rect 71 -23090 331 -23030
rect 391 -23090 400 -23030
rect 0 -23380 14 -23090
rect 66 -23380 400 -23090
rect 0 -23440 11 -23380
rect 71 -23440 331 -23380
rect 391 -23440 400 -23380
rect 0 -23524 14 -23440
rect 66 -23450 400 -23440
rect 457 -23030 857 -23020
rect 457 -23090 467 -23030
rect 527 -23090 787 -23030
rect 847 -23090 857 -23030
rect 457 -23200 857 -23090
rect 913 -23030 1313 -23020
rect 913 -23090 923 -23030
rect 983 -23090 1243 -23030
rect 1303 -23090 1313 -23030
rect 913 -23200 1313 -23090
rect 1371 -23030 1771 -23020
rect 1371 -23090 1381 -23030
rect 1441 -23090 1701 -23030
rect 1761 -23090 1771 -23030
rect 1371 -23200 1771 -23090
rect 1827 -23030 2227 -23020
rect 1827 -23090 1837 -23030
rect 1897 -23090 2157 -23030
rect 2217 -23090 2227 -23030
rect 1827 -23200 2227 -23090
rect 2283 -23030 2683 -23020
rect 2283 -23090 2293 -23030
rect 2353 -23090 2613 -23030
rect 2673 -23090 2683 -23030
rect 2283 -23200 2683 -23090
rect 2741 -23030 3141 -23020
rect 2741 -23090 2751 -23030
rect 2811 -23090 3071 -23030
rect 3131 -23090 3141 -23030
rect 2741 -23200 3141 -23090
rect 3197 -23030 3597 -23020
rect 3197 -23090 3207 -23030
rect 3267 -23090 3527 -23030
rect 3587 -23090 3597 -23030
rect 3197 -23200 3597 -23090
rect 3653 -23030 4053 -23020
rect 3653 -23090 3663 -23030
rect 3723 -23090 3983 -23030
rect 4043 -23090 4053 -23030
rect 3653 -23200 4053 -23090
rect 457 -23271 4053 -23200
rect 457 -23380 857 -23271
rect 457 -23440 467 -23380
rect 527 -23440 787 -23380
rect 847 -23440 857 -23380
rect 457 -23450 857 -23440
rect 913 -23380 1313 -23271
rect 913 -23440 923 -23380
rect 983 -23440 1243 -23380
rect 1303 -23440 1313 -23380
rect 913 -23450 1313 -23440
rect 1371 -23380 1771 -23271
rect 1371 -23440 1381 -23380
rect 1441 -23440 1701 -23380
rect 1761 -23440 1771 -23380
rect 1371 -23450 1771 -23440
rect 1827 -23380 2227 -23271
rect 1827 -23440 1837 -23380
rect 1897 -23440 2157 -23380
rect 2217 -23440 2227 -23380
rect 1827 -23450 2227 -23440
rect 2283 -23380 2683 -23271
rect 2283 -23440 2293 -23380
rect 2353 -23440 2613 -23380
rect 2673 -23440 2683 -23380
rect 2283 -23450 2683 -23440
rect 2741 -23380 3141 -23271
rect 2741 -23440 2751 -23380
rect 2811 -23440 3071 -23380
rect 3131 -23440 3141 -23380
rect 2741 -23450 3141 -23440
rect 3197 -23380 3597 -23271
rect 3197 -23440 3207 -23380
rect 3267 -23440 3527 -23380
rect 3587 -23440 3597 -23380
rect 3197 -23450 3597 -23440
rect 3653 -23380 4053 -23271
rect 3653 -23440 3663 -23380
rect 3723 -23440 3983 -23380
rect 4043 -23440 4053 -23380
rect 3653 -23450 4053 -23440
rect 4111 -23030 4511 -23020
rect 4111 -23090 4121 -23030
rect 4181 -23090 4441 -23030
rect 4501 -23090 4511 -23030
rect 4111 -23200 4511 -23090
rect 4567 -23030 4967 -23020
rect 4567 -23090 4577 -23030
rect 4637 -23090 4897 -23030
rect 4957 -23090 4967 -23030
rect 4567 -23200 4967 -23090
rect 5023 -23030 5423 -23020
rect 5023 -23090 5033 -23030
rect 5093 -23090 5353 -23030
rect 5413 -23090 5423 -23030
rect 5023 -23200 5423 -23090
rect 5481 -23030 5881 -23020
rect 5481 -23090 5491 -23030
rect 5551 -23090 5811 -23030
rect 5871 -23090 5881 -23030
rect 5481 -23200 5881 -23090
rect 5937 -23030 6337 -23020
rect 5937 -23090 5947 -23030
rect 6007 -23090 6267 -23030
rect 6327 -23090 6337 -23030
rect 5937 -23200 6337 -23090
rect 6393 -23030 6793 -23020
rect 6393 -23090 6403 -23030
rect 6463 -23090 6723 -23030
rect 6783 -23090 6793 -23030
rect 6393 -23200 6793 -23090
rect 6851 -23030 7251 -23020
rect 6851 -23090 6861 -23030
rect 6921 -23090 7181 -23030
rect 7241 -23090 7251 -23030
rect 6851 -23200 7251 -23090
rect 4111 -23271 7251 -23200
rect 4111 -23380 4511 -23271
rect 4111 -23440 4121 -23380
rect 4181 -23440 4441 -23380
rect 4501 -23440 4511 -23380
rect 4111 -23450 4511 -23440
rect 4567 -23380 4967 -23271
rect 4567 -23440 4577 -23380
rect 4637 -23440 4897 -23380
rect 4957 -23440 4967 -23380
rect 4567 -23450 4967 -23440
rect 5023 -23380 5423 -23271
rect 5023 -23440 5033 -23380
rect 5093 -23440 5353 -23380
rect 5413 -23440 5423 -23380
rect 5023 -23450 5423 -23440
rect 5481 -23380 5881 -23271
rect 5481 -23440 5491 -23380
rect 5551 -23440 5811 -23380
rect 5871 -23440 5881 -23380
rect 5481 -23450 5881 -23440
rect 5937 -23380 6337 -23271
rect 5937 -23440 5947 -23380
rect 6007 -23440 6267 -23380
rect 6327 -23440 6337 -23380
rect 5937 -23450 6337 -23440
rect 6393 -23380 6793 -23271
rect 6393 -23440 6403 -23380
rect 6463 -23440 6723 -23380
rect 6783 -23440 6793 -23380
rect 6393 -23450 6793 -23440
rect 6851 -23380 7251 -23271
rect 6851 -23440 6861 -23380
rect 6921 -23440 7181 -23380
rect 7241 -23440 7251 -23380
rect 6851 -23450 7251 -23440
rect 7307 -23030 7707 -23020
rect 7307 -23090 7317 -23030
rect 7377 -23090 7637 -23030
rect 7697 -23090 7707 -23030
rect 7307 -23200 7707 -23090
rect 7763 -23030 8163 -23020
rect 7763 -23090 7773 -23030
rect 7833 -23090 8093 -23030
rect 8153 -23090 8163 -23030
rect 7763 -23200 8163 -23090
rect 8237 -23030 8637 -23020
rect 8237 -23090 8247 -23030
rect 8307 -23090 8567 -23030
rect 8627 -23090 8637 -23030
rect 8237 -23200 8637 -23090
rect 8693 -23030 9093 -23020
rect 8693 -23090 8703 -23030
rect 8763 -23090 9023 -23030
rect 9083 -23090 9093 -23030
rect 8693 -23200 9093 -23090
rect 9151 -23030 9551 -23020
rect 9151 -23090 9161 -23030
rect 9221 -23090 9481 -23030
rect 9541 -23090 9551 -23030
rect 9151 -23200 9551 -23090
rect 9607 -23030 10007 -23020
rect 9607 -23090 9617 -23030
rect 9677 -23090 9937 -23030
rect 9997 -23090 10007 -23030
rect 9607 -23200 10007 -23090
rect 10063 -23030 10463 -23020
rect 10063 -23090 10073 -23030
rect 10133 -23090 10393 -23030
rect 10453 -23090 10463 -23030
rect 10063 -23200 10463 -23090
rect 10521 -23030 10921 -23020
rect 10521 -23090 10531 -23030
rect 10591 -23090 10851 -23030
rect 10911 -23090 10921 -23030
rect 10521 -23200 10921 -23090
rect 10977 -23030 11377 -23020
rect 10977 -23090 10987 -23030
rect 11047 -23090 11307 -23030
rect 11367 -23090 11377 -23030
rect 10977 -23200 11377 -23090
rect 11433 -23030 11833 -23020
rect 11433 -23090 11443 -23030
rect 11503 -23090 11763 -23030
rect 11823 -23090 11833 -23030
rect 11433 -23200 11833 -23090
rect 11891 -23030 12291 -23020
rect 11891 -23090 11901 -23030
rect 11961 -23090 12221 -23030
rect 12281 -23090 12291 -23030
rect 11891 -23200 12291 -23090
rect 12347 -23030 12747 -23020
rect 12347 -23090 12357 -23030
rect 12417 -23090 12677 -23030
rect 12737 -23090 12747 -23030
rect 12347 -23200 12747 -23090
rect 12803 -23030 13203 -23020
rect 12803 -23090 12813 -23030
rect 12873 -23090 13133 -23030
rect 13193 -23090 13203 -23030
rect 12803 -23200 13203 -23090
rect 13261 -23030 13661 -23020
rect 13261 -23090 13271 -23030
rect 13331 -23090 13591 -23030
rect 13651 -23090 13661 -23030
rect 13261 -23200 13661 -23090
rect 13717 -23030 14117 -23020
rect 13717 -23090 13727 -23030
rect 13787 -23090 14047 -23030
rect 14107 -23090 14117 -23030
rect 13717 -23200 14117 -23090
rect 14173 -23030 14573 -23020
rect 14173 -23090 14183 -23030
rect 14243 -23090 14503 -23030
rect 14563 -23090 14573 -23030
rect 14173 -23200 14573 -23090
rect 14631 -23030 15031 -23020
rect 14631 -23090 14641 -23030
rect 14701 -23090 14961 -23030
rect 15021 -23090 15031 -23030
rect 14631 -23200 15031 -23090
rect 15087 -23030 15487 -23020
rect 15087 -23090 15097 -23030
rect 15157 -23090 15417 -23030
rect 15477 -23090 15487 -23030
rect 15087 -23200 15487 -23090
rect 7307 -23271 15487 -23200
rect 7307 -23380 7707 -23271
rect 7307 -23440 7317 -23380
rect 7377 -23440 7637 -23380
rect 7697 -23440 7707 -23380
rect 7307 -23450 7707 -23440
rect 7763 -23380 8163 -23271
rect 7763 -23440 7773 -23380
rect 7833 -23440 8093 -23380
rect 8153 -23440 8163 -23380
rect 7763 -23450 8163 -23440
rect 8237 -23380 8637 -23271
rect 8237 -23440 8247 -23380
rect 8307 -23440 8567 -23380
rect 8627 -23440 8637 -23380
rect 8237 -23450 8637 -23440
rect 8693 -23380 9093 -23271
rect 8693 -23440 8703 -23380
rect 8763 -23440 9023 -23380
rect 9083 -23440 9093 -23380
rect 8693 -23450 9093 -23440
rect 9151 -23380 9551 -23271
rect 9151 -23440 9161 -23380
rect 9221 -23440 9481 -23380
rect 9541 -23440 9551 -23380
rect 9151 -23450 9551 -23440
rect 9607 -23380 10007 -23271
rect 9607 -23440 9617 -23380
rect 9677 -23440 9937 -23380
rect 9997 -23440 10007 -23380
rect 9607 -23450 10007 -23440
rect 10063 -23380 10463 -23271
rect 10063 -23440 10073 -23380
rect 10133 -23440 10393 -23380
rect 10453 -23440 10463 -23380
rect 10063 -23450 10463 -23440
rect 10521 -23380 10921 -23271
rect 10521 -23440 10531 -23380
rect 10591 -23440 10851 -23380
rect 10911 -23440 10921 -23380
rect 10521 -23450 10921 -23440
rect 10977 -23380 11377 -23271
rect 10977 -23440 10987 -23380
rect 11047 -23440 11307 -23380
rect 11367 -23440 11377 -23380
rect 10977 -23450 11377 -23440
rect 11433 -23380 11833 -23271
rect 11433 -23440 11443 -23380
rect 11503 -23440 11763 -23380
rect 11823 -23440 11833 -23380
rect 11433 -23450 11833 -23440
rect 11891 -23380 12291 -23271
rect 11891 -23440 11901 -23380
rect 11961 -23440 12221 -23380
rect 12281 -23440 12291 -23380
rect 11891 -23450 12291 -23440
rect 12347 -23380 12747 -23271
rect 12347 -23440 12357 -23380
rect 12417 -23440 12677 -23380
rect 12737 -23440 12747 -23380
rect 12347 -23450 12747 -23440
rect 12803 -23380 13203 -23271
rect 12803 -23440 12813 -23380
rect 12873 -23440 13133 -23380
rect 13193 -23440 13203 -23380
rect 12803 -23450 13203 -23440
rect 13261 -23380 13661 -23271
rect 13261 -23440 13271 -23380
rect 13331 -23440 13591 -23380
rect 13651 -23440 13661 -23380
rect 13261 -23450 13661 -23440
rect 13717 -23380 14117 -23271
rect 13717 -23440 13727 -23380
rect 13787 -23440 14047 -23380
rect 14107 -23440 14117 -23380
rect 13717 -23450 14117 -23440
rect 14173 -23380 14573 -23271
rect 14173 -23440 14183 -23380
rect 14243 -23440 14503 -23380
rect 14563 -23440 14573 -23380
rect 14173 -23450 14573 -23440
rect 14631 -23380 15031 -23271
rect 14631 -23440 14641 -23380
rect 14701 -23440 14961 -23380
rect 15021 -23440 15031 -23380
rect 14631 -23450 15031 -23440
rect 15087 -23380 15487 -23271
rect 15087 -23440 15097 -23380
rect 15157 -23440 15417 -23380
rect 15477 -23440 15487 -23380
rect 15087 -23450 15487 -23440
rect 66 -23514 80 -23450
rect 457 -23514 527 -23450
rect 913 -23514 983 -23450
rect 1371 -23514 1441 -23450
rect 1827 -23514 1897 -23450
rect 2283 -23514 2353 -23450
rect 2741 -23514 2811 -23450
rect 3197 -23514 3267 -23450
rect 3653 -23514 3723 -23450
rect 4111 -23514 4181 -23450
rect 4567 -23514 4637 -23450
rect 5023 -23514 5093 -23450
rect 5481 -23514 5551 -23450
rect 5937 -23514 6007 -23450
rect 6393 -23514 6463 -23450
rect 6851 -23514 6921 -23450
rect 66 -23524 400 -23514
rect 0 -23584 11 -23524
rect 71 -23584 331 -23524
rect 391 -23584 400 -23524
rect 0 -23874 14 -23584
rect 66 -23874 400 -23584
rect 0 -23934 11 -23874
rect 71 -23934 331 -23874
rect 391 -23934 400 -23874
rect 0 -24016 14 -23934
rect 66 -23944 400 -23934
rect 457 -23524 857 -23514
rect 457 -23584 467 -23524
rect 527 -23584 787 -23524
rect 847 -23584 857 -23524
rect 457 -23694 857 -23584
rect 913 -23524 1313 -23514
rect 913 -23584 923 -23524
rect 983 -23584 1243 -23524
rect 1303 -23584 1313 -23524
rect 913 -23694 1313 -23584
rect 1371 -23524 1771 -23514
rect 1371 -23584 1381 -23524
rect 1441 -23584 1701 -23524
rect 1761 -23584 1771 -23524
rect 1371 -23694 1771 -23584
rect 1827 -23524 2227 -23514
rect 1827 -23584 1837 -23524
rect 1897 -23584 2157 -23524
rect 2217 -23584 2227 -23524
rect 1827 -23694 2227 -23584
rect 2283 -23524 2683 -23514
rect 2283 -23584 2293 -23524
rect 2353 -23584 2613 -23524
rect 2673 -23584 2683 -23524
rect 2283 -23694 2683 -23584
rect 457 -23697 2683 -23694
rect 2741 -23524 3141 -23514
rect 2741 -23584 2751 -23524
rect 2811 -23584 3071 -23524
rect 3131 -23584 3141 -23524
rect 2741 -23694 3141 -23584
rect 3197 -23524 3597 -23514
rect 3197 -23584 3207 -23524
rect 3267 -23584 3527 -23524
rect 3587 -23584 3597 -23524
rect 3197 -23694 3597 -23584
rect 3653 -23524 4053 -23514
rect 3653 -23584 3663 -23524
rect 3723 -23584 3983 -23524
rect 4043 -23584 4053 -23524
rect 3653 -23694 4053 -23584
rect 2741 -23697 4053 -23694
rect 457 -23767 4053 -23697
rect 457 -23874 857 -23767
rect 457 -23934 467 -23874
rect 527 -23934 787 -23874
rect 847 -23934 857 -23874
rect 457 -23944 857 -23934
rect 913 -23874 1313 -23767
rect 913 -23934 923 -23874
rect 983 -23934 1243 -23874
rect 1303 -23934 1313 -23874
rect 913 -23944 1313 -23934
rect 1371 -23874 1771 -23767
rect 1371 -23934 1381 -23874
rect 1441 -23934 1701 -23874
rect 1761 -23934 1771 -23874
rect 1371 -23944 1771 -23934
rect 1827 -23874 2227 -23767
rect 1827 -23934 1837 -23874
rect 1897 -23934 2157 -23874
rect 2217 -23934 2227 -23874
rect 1827 -23944 2227 -23934
rect 2283 -23874 2683 -23767
rect 2283 -23934 2293 -23874
rect 2353 -23934 2613 -23874
rect 2673 -23934 2683 -23874
rect 2283 -23944 2683 -23934
rect 2741 -23874 3141 -23767
rect 2741 -23934 2751 -23874
rect 2811 -23934 3071 -23874
rect 3131 -23934 3141 -23874
rect 2741 -23944 3141 -23934
rect 3197 -23874 3597 -23767
rect 3197 -23934 3207 -23874
rect 3267 -23934 3527 -23874
rect 3587 -23934 3597 -23874
rect 3197 -23944 3597 -23934
rect 3653 -23874 4053 -23767
rect 3653 -23934 3663 -23874
rect 3723 -23934 3983 -23874
rect 4043 -23934 4053 -23874
rect 3653 -23944 4053 -23934
rect 4111 -23524 4511 -23514
rect 4111 -23584 4121 -23524
rect 4181 -23584 4441 -23524
rect 4501 -23584 4511 -23524
rect 4111 -23694 4511 -23584
rect 4567 -23524 4967 -23514
rect 4567 -23584 4577 -23524
rect 4637 -23584 4897 -23524
rect 4957 -23584 4967 -23524
rect 4567 -23694 4967 -23584
rect 5023 -23524 5423 -23514
rect 5023 -23584 5033 -23524
rect 5093 -23584 5353 -23524
rect 5413 -23584 5423 -23524
rect 5023 -23694 5423 -23584
rect 5481 -23524 5881 -23514
rect 5481 -23584 5491 -23524
rect 5551 -23584 5811 -23524
rect 5871 -23584 5881 -23524
rect 5481 -23694 5881 -23584
rect 5937 -23524 6337 -23514
rect 5937 -23584 5947 -23524
rect 6007 -23584 6267 -23524
rect 6327 -23584 6337 -23524
rect 5937 -23694 6337 -23584
rect 6393 -23524 6793 -23514
rect 6393 -23584 6403 -23524
rect 6463 -23584 6723 -23524
rect 6783 -23584 6793 -23524
rect 6393 -23694 6793 -23584
rect 6851 -23524 7251 -23514
rect 6851 -23584 6861 -23524
rect 6921 -23584 7181 -23524
rect 7241 -23584 7251 -23524
rect 6851 -23694 7251 -23584
rect 7307 -23524 7707 -23514
rect 7307 -23584 7317 -23524
rect 7377 -23584 7637 -23524
rect 7697 -23584 7707 -23524
rect 7307 -23694 7707 -23584
rect 7763 -23524 8163 -23514
rect 7763 -23584 7773 -23524
rect 7833 -23584 8093 -23524
rect 8153 -23584 8163 -23524
rect 7763 -23694 8163 -23584
rect 8237 -23524 8637 -23514
rect 8237 -23584 8247 -23524
rect 8307 -23584 8567 -23524
rect 8627 -23584 8637 -23524
rect 8237 -23694 8637 -23584
rect 8693 -23524 9093 -23514
rect 8693 -23584 8703 -23524
rect 8763 -23584 9023 -23524
rect 9083 -23584 9093 -23524
rect 8693 -23694 9093 -23584
rect 9151 -23524 9551 -23514
rect 9151 -23584 9161 -23524
rect 9221 -23584 9481 -23524
rect 9541 -23584 9551 -23524
rect 9151 -23694 9551 -23584
rect 9607 -23524 10007 -23514
rect 9607 -23584 9617 -23524
rect 9677 -23584 9937 -23524
rect 9997 -23584 10007 -23524
rect 9607 -23694 10007 -23584
rect 10063 -23524 10463 -23514
rect 10063 -23584 10073 -23524
rect 10133 -23584 10393 -23524
rect 10453 -23584 10463 -23524
rect 10063 -23694 10463 -23584
rect 4111 -23697 10463 -23694
rect 10521 -23524 10921 -23514
rect 10521 -23584 10531 -23524
rect 10591 -23584 10851 -23524
rect 10911 -23584 10921 -23524
rect 10521 -23694 10921 -23584
rect 10977 -23524 11377 -23514
rect 10977 -23584 10987 -23524
rect 11047 -23584 11307 -23524
rect 11367 -23584 11377 -23524
rect 10977 -23694 11377 -23584
rect 11433 -23524 11833 -23514
rect 11433 -23584 11443 -23524
rect 11503 -23584 11763 -23524
rect 11823 -23584 11833 -23524
rect 11433 -23694 11833 -23584
rect 11891 -23524 12291 -23514
rect 11891 -23584 11901 -23524
rect 11961 -23584 12221 -23524
rect 12281 -23584 12291 -23524
rect 11891 -23694 12291 -23584
rect 12347 -23524 12747 -23514
rect 12347 -23584 12357 -23524
rect 12417 -23584 12677 -23524
rect 12737 -23584 12747 -23524
rect 12347 -23694 12747 -23584
rect 12803 -23524 13203 -23514
rect 12803 -23584 12813 -23524
rect 12873 -23584 13133 -23524
rect 13193 -23584 13203 -23524
rect 12803 -23694 13203 -23584
rect 13261 -23524 13661 -23514
rect 13261 -23584 13271 -23524
rect 13331 -23584 13591 -23524
rect 13651 -23584 13661 -23524
rect 13261 -23694 13661 -23584
rect 13717 -23524 14117 -23514
rect 13717 -23584 13727 -23524
rect 13787 -23584 14047 -23524
rect 14107 -23584 14117 -23524
rect 13717 -23694 14117 -23584
rect 14173 -23524 14573 -23514
rect 14173 -23584 14183 -23524
rect 14243 -23584 14503 -23524
rect 14563 -23584 14573 -23524
rect 14173 -23694 14573 -23584
rect 14631 -23524 15031 -23514
rect 14631 -23584 14641 -23524
rect 14701 -23584 14961 -23524
rect 15021 -23584 15031 -23524
rect 14631 -23694 15031 -23584
rect 15087 -23524 15487 -23514
rect 15087 -23584 15097 -23524
rect 15157 -23584 15417 -23524
rect 15477 -23584 15487 -23524
rect 15087 -23694 15487 -23584
rect 10521 -23695 15487 -23694
rect 10521 -23697 15721 -23695
rect 4111 -23766 15721 -23697
rect 4111 -23767 15487 -23766
rect 4111 -23874 4511 -23767
rect 4111 -23934 4121 -23874
rect 4181 -23934 4441 -23874
rect 4501 -23934 4511 -23874
rect 4111 -23944 4511 -23934
rect 4567 -23874 4967 -23767
rect 4567 -23934 4577 -23874
rect 4637 -23934 4897 -23874
rect 4957 -23934 4967 -23874
rect 4567 -23944 4967 -23934
rect 5023 -23874 5423 -23767
rect 5023 -23934 5033 -23874
rect 5093 -23934 5353 -23874
rect 5413 -23934 5423 -23874
rect 5023 -23944 5423 -23934
rect 5481 -23874 5881 -23767
rect 5481 -23934 5491 -23874
rect 5551 -23934 5811 -23874
rect 5871 -23934 5881 -23874
rect 5481 -23944 5881 -23934
rect 5937 -23874 6337 -23767
rect 5937 -23934 5947 -23874
rect 6007 -23934 6267 -23874
rect 6327 -23934 6337 -23874
rect 5937 -23944 6337 -23934
rect 6393 -23874 6793 -23767
rect 6393 -23934 6403 -23874
rect 6463 -23934 6723 -23874
rect 6783 -23934 6793 -23874
rect 6393 -23944 6793 -23934
rect 6851 -23874 7251 -23767
rect 6851 -23934 6861 -23874
rect 6921 -23934 7181 -23874
rect 7241 -23934 7251 -23874
rect 6851 -23944 7251 -23934
rect 7307 -23874 7707 -23767
rect 7307 -23934 7317 -23874
rect 7377 -23934 7637 -23874
rect 7697 -23934 7707 -23874
rect 7307 -23944 7707 -23934
rect 7763 -23874 8163 -23767
rect 7763 -23934 7773 -23874
rect 7833 -23934 8093 -23874
rect 8153 -23934 8163 -23874
rect 7763 -23944 8163 -23934
rect 8237 -23874 8637 -23767
rect 8237 -23934 8247 -23874
rect 8307 -23934 8567 -23874
rect 8627 -23934 8637 -23874
rect 8237 -23944 8637 -23934
rect 8693 -23874 9093 -23767
rect 8693 -23934 8703 -23874
rect 8763 -23934 9023 -23874
rect 9083 -23934 9093 -23874
rect 8693 -23944 9093 -23934
rect 9151 -23874 9551 -23767
rect 9151 -23934 9161 -23874
rect 9221 -23934 9481 -23874
rect 9541 -23934 9551 -23874
rect 9151 -23944 9551 -23934
rect 9607 -23874 10007 -23767
rect 9607 -23934 9617 -23874
rect 9677 -23934 9937 -23874
rect 9997 -23934 10007 -23874
rect 9607 -23944 10007 -23934
rect 10063 -23874 10463 -23767
rect 10063 -23934 10073 -23874
rect 10133 -23934 10393 -23874
rect 10453 -23934 10463 -23874
rect 10063 -23944 10463 -23934
rect 10521 -23874 10921 -23767
rect 10521 -23934 10531 -23874
rect 10591 -23934 10851 -23874
rect 10911 -23934 10921 -23874
rect 10521 -23944 10921 -23934
rect 10977 -23874 11377 -23767
rect 10977 -23934 10987 -23874
rect 11047 -23934 11307 -23874
rect 11367 -23934 11377 -23874
rect 10977 -23944 11377 -23934
rect 11433 -23874 11833 -23767
rect 11433 -23934 11443 -23874
rect 11503 -23934 11763 -23874
rect 11823 -23934 11833 -23874
rect 11433 -23944 11833 -23934
rect 11891 -23874 12291 -23767
rect 11891 -23934 11901 -23874
rect 11961 -23934 12221 -23874
rect 12281 -23934 12291 -23874
rect 11891 -23944 12291 -23934
rect 12347 -23874 12747 -23767
rect 12347 -23934 12357 -23874
rect 12417 -23934 12677 -23874
rect 12737 -23934 12747 -23874
rect 12347 -23944 12747 -23934
rect 12803 -23874 13203 -23767
rect 12803 -23934 12813 -23874
rect 12873 -23934 13133 -23874
rect 13193 -23934 13203 -23874
rect 12803 -23944 13203 -23934
rect 13261 -23874 13661 -23767
rect 13261 -23934 13271 -23874
rect 13331 -23934 13591 -23874
rect 13651 -23934 13661 -23874
rect 13261 -23944 13661 -23934
rect 13717 -23874 14117 -23767
rect 13717 -23934 13727 -23874
rect 13787 -23934 14047 -23874
rect 14107 -23934 14117 -23874
rect 13717 -23944 14117 -23934
rect 14173 -23874 14573 -23767
rect 14173 -23934 14183 -23874
rect 14243 -23934 14503 -23874
rect 14563 -23934 14573 -23874
rect 14173 -23944 14573 -23934
rect 14631 -23874 15031 -23767
rect 14631 -23934 14641 -23874
rect 14701 -23934 14961 -23874
rect 15021 -23934 15031 -23874
rect 14631 -23944 15031 -23934
rect 15087 -23874 15487 -23767
rect 15087 -23934 15097 -23874
rect 15157 -23934 15417 -23874
rect 15477 -23934 15487 -23874
rect 15087 -23944 15487 -23934
rect 66 -24006 80 -23944
rect 457 -24006 528 -23944
rect 913 -24006 984 -23944
rect 1371 -24006 1442 -23944
rect 1827 -24006 1898 -23944
rect 2283 -24006 2354 -23944
rect 2741 -24006 2811 -23944
rect 3197 -24006 3267 -23944
rect 3653 -24006 3723 -23944
rect 4111 -24006 4181 -23944
rect 4567 -24006 4637 -23944
rect 5023 -24006 5093 -23944
rect 5481 -24006 5551 -23944
rect 5937 -24006 6007 -23944
rect 6393 -24006 6463 -23944
rect 6851 -24006 6921 -23944
rect 7307 -24006 7377 -23944
rect 7763 -24006 7833 -23944
rect 8237 -24006 8307 -23944
rect 8693 -24006 8763 -23944
rect 9151 -24006 9221 -23944
rect 9607 -24006 9677 -23944
rect 10063 -24006 10133 -23944
rect 10521 -24006 10591 -23944
rect 10977 -24006 11047 -23944
rect 11433 -24006 11503 -23944
rect 11891 -24006 11961 -23944
rect 12347 -24006 12417 -23944
rect 12803 -24006 12873 -23944
rect 13261 -24006 13331 -23944
rect 13717 -24006 13787 -23944
rect 14173 -24006 14243 -23944
rect 14631 -24006 14701 -23944
rect 66 -24016 400 -24006
rect 0 -24076 11 -24016
rect 71 -24076 331 -24016
rect 391 -24076 400 -24016
rect 0 -24366 14 -24076
rect 66 -24366 400 -24076
rect 0 -24426 11 -24366
rect 71 -24426 331 -24366
rect 391 -24426 400 -24366
rect 0 -24518 14 -24426
rect 66 -24436 400 -24426
rect 457 -24016 857 -24006
rect 457 -24076 467 -24016
rect 527 -24076 787 -24016
rect 847 -24076 857 -24016
rect 457 -24186 857 -24076
rect 913 -24016 1313 -24006
rect 913 -24076 923 -24016
rect 983 -24076 1243 -24016
rect 1303 -24076 1313 -24016
rect 913 -24186 1313 -24076
rect 1371 -24016 1771 -24006
rect 1371 -24076 1381 -24016
rect 1441 -24076 1701 -24016
rect 1761 -24076 1771 -24016
rect 1371 -24186 1771 -24076
rect 1827 -24016 2227 -24006
rect 1827 -24076 1837 -24016
rect 1897 -24076 2157 -24016
rect 2217 -24076 2227 -24016
rect 1827 -24186 2227 -24076
rect 2283 -24016 2683 -24006
rect 2283 -24076 2293 -24016
rect 2353 -24076 2613 -24016
rect 2673 -24076 2683 -24016
rect 2283 -24186 2683 -24076
rect 457 -24187 2683 -24186
rect 2741 -24016 3141 -24006
rect 2741 -24076 2751 -24016
rect 2811 -24076 3071 -24016
rect 3131 -24076 3141 -24016
rect 2741 -24186 3141 -24076
rect 3197 -24016 3597 -24006
rect 3197 -24076 3207 -24016
rect 3267 -24076 3527 -24016
rect 3587 -24076 3597 -24016
rect 3197 -24186 3597 -24076
rect 3653 -24016 4053 -24006
rect 3653 -24076 3663 -24016
rect 3723 -24076 3983 -24016
rect 4043 -24076 4053 -24016
rect 3653 -24186 4053 -24076
rect 2741 -24187 4053 -24186
rect 457 -24257 4053 -24187
rect 457 -24366 857 -24257
rect 457 -24426 467 -24366
rect 527 -24426 787 -24366
rect 847 -24426 857 -24366
rect 457 -24436 857 -24426
rect 913 -24366 1313 -24257
rect 913 -24426 923 -24366
rect 983 -24426 1243 -24366
rect 1303 -24426 1313 -24366
rect 913 -24436 1313 -24426
rect 1371 -24366 1771 -24257
rect 1371 -24426 1381 -24366
rect 1441 -24426 1701 -24366
rect 1761 -24426 1771 -24366
rect 1371 -24436 1771 -24426
rect 1827 -24366 2227 -24257
rect 1827 -24426 1837 -24366
rect 1897 -24426 2157 -24366
rect 2217 -24426 2227 -24366
rect 1827 -24436 2227 -24426
rect 2283 -24366 2683 -24257
rect 2283 -24426 2293 -24366
rect 2353 -24426 2613 -24366
rect 2673 -24426 2683 -24366
rect 2283 -24436 2683 -24426
rect 2741 -24366 3141 -24257
rect 2741 -24426 2751 -24366
rect 2811 -24426 3071 -24366
rect 3131 -24426 3141 -24366
rect 2741 -24436 3141 -24426
rect 3197 -24366 3597 -24257
rect 3197 -24426 3207 -24366
rect 3267 -24426 3527 -24366
rect 3587 -24426 3597 -24366
rect 3197 -24436 3597 -24426
rect 3653 -24366 4053 -24257
rect 3653 -24426 3663 -24366
rect 3723 -24426 3983 -24366
rect 4043 -24426 4053 -24366
rect 3653 -24436 4053 -24426
rect 4111 -24016 4511 -24006
rect 4111 -24076 4121 -24016
rect 4181 -24076 4441 -24016
rect 4501 -24076 4511 -24016
rect 4111 -24186 4511 -24076
rect 4567 -24016 4967 -24006
rect 4567 -24076 4577 -24016
rect 4637 -24076 4897 -24016
rect 4957 -24076 4967 -24016
rect 4567 -24186 4967 -24076
rect 5023 -24016 5423 -24006
rect 5023 -24076 5033 -24016
rect 5093 -24076 5353 -24016
rect 5413 -24076 5423 -24016
rect 5023 -24186 5423 -24076
rect 5481 -24016 5881 -24006
rect 5481 -24076 5491 -24016
rect 5551 -24076 5811 -24016
rect 5871 -24076 5881 -24016
rect 5481 -24186 5881 -24076
rect 5937 -24016 6337 -24006
rect 5937 -24076 5947 -24016
rect 6007 -24076 6267 -24016
rect 6327 -24076 6337 -24016
rect 5937 -24186 6337 -24076
rect 6393 -24016 6793 -24006
rect 6393 -24076 6403 -24016
rect 6463 -24076 6723 -24016
rect 6783 -24076 6793 -24016
rect 6393 -24186 6793 -24076
rect 6851 -24016 7251 -24006
rect 6851 -24076 6861 -24016
rect 6921 -24076 7181 -24016
rect 7241 -24076 7251 -24016
rect 6851 -24186 7251 -24076
rect 7307 -24016 7707 -24006
rect 7307 -24076 7317 -24016
rect 7377 -24076 7637 -24016
rect 7697 -24076 7707 -24016
rect 7307 -24186 7707 -24076
rect 7763 -24016 8163 -24006
rect 7763 -24076 7773 -24016
rect 7833 -24076 8093 -24016
rect 8153 -24076 8163 -24016
rect 7763 -24186 8163 -24076
rect 8237 -24016 8637 -24006
rect 8237 -24076 8247 -24016
rect 8307 -24076 8567 -24016
rect 8627 -24076 8637 -24016
rect 8237 -24186 8637 -24076
rect 8693 -24016 9093 -24006
rect 8693 -24076 8703 -24016
rect 8763 -24076 9023 -24016
rect 9083 -24076 9093 -24016
rect 8693 -24186 9093 -24076
rect 9151 -24016 9551 -24006
rect 9151 -24076 9161 -24016
rect 9221 -24076 9481 -24016
rect 9541 -24076 9551 -24016
rect 9151 -24186 9551 -24076
rect 9607 -24016 10007 -24006
rect 9607 -24076 9617 -24016
rect 9677 -24076 9937 -24016
rect 9997 -24076 10007 -24016
rect 9607 -24186 10007 -24076
rect 10063 -24016 10463 -24006
rect 10063 -24076 10073 -24016
rect 10133 -24076 10393 -24016
rect 10453 -24076 10463 -24016
rect 10063 -24186 10463 -24076
rect 4111 -24187 10463 -24186
rect 10521 -24016 10921 -24006
rect 10521 -24076 10531 -24016
rect 10591 -24076 10851 -24016
rect 10911 -24076 10921 -24016
rect 10521 -24186 10921 -24076
rect 10977 -24016 11377 -24006
rect 10977 -24076 10987 -24016
rect 11047 -24076 11307 -24016
rect 11367 -24076 11377 -24016
rect 10977 -24186 11377 -24076
rect 11433 -24016 11833 -24006
rect 11433 -24076 11443 -24016
rect 11503 -24076 11763 -24016
rect 11823 -24076 11833 -24016
rect 11433 -24186 11833 -24076
rect 11891 -24016 12291 -24006
rect 11891 -24076 11901 -24016
rect 11961 -24076 12221 -24016
rect 12281 -24076 12291 -24016
rect 11891 -24186 12291 -24076
rect 12347 -24016 12747 -24006
rect 12347 -24076 12357 -24016
rect 12417 -24076 12677 -24016
rect 12737 -24076 12747 -24016
rect 12347 -24186 12747 -24076
rect 12803 -24016 13203 -24006
rect 12803 -24076 12813 -24016
rect 12873 -24076 13133 -24016
rect 13193 -24076 13203 -24016
rect 12803 -24186 13203 -24076
rect 13261 -24016 13661 -24006
rect 13261 -24076 13271 -24016
rect 13331 -24076 13591 -24016
rect 13651 -24076 13661 -24016
rect 13261 -24186 13661 -24076
rect 13717 -24016 14117 -24006
rect 13717 -24076 13727 -24016
rect 13787 -24076 14047 -24016
rect 14107 -24076 14117 -24016
rect 13717 -24186 14117 -24076
rect 14173 -24016 14573 -24006
rect 14173 -24076 14183 -24016
rect 14243 -24076 14503 -24016
rect 14563 -24076 14573 -24016
rect 14173 -24186 14573 -24076
rect 14631 -24016 15031 -24006
rect 14631 -24076 14641 -24016
rect 14701 -24076 14961 -24016
rect 15021 -24076 15031 -24016
rect 14631 -24186 15031 -24076
rect 15087 -24016 15487 -24006
rect 15087 -24076 15097 -24016
rect 15157 -24076 15417 -24016
rect 15477 -24076 15487 -24016
rect 15087 -24186 15487 -24076
rect 10521 -24187 15487 -24186
rect 4111 -24257 15487 -24187
rect 4111 -24366 4511 -24257
rect 4111 -24426 4121 -24366
rect 4181 -24426 4441 -24366
rect 4501 -24426 4511 -24366
rect 4111 -24436 4511 -24426
rect 4567 -24366 4967 -24257
rect 4567 -24426 4577 -24366
rect 4637 -24426 4897 -24366
rect 4957 -24426 4967 -24366
rect 4567 -24436 4967 -24426
rect 5023 -24366 5423 -24257
rect 5023 -24426 5033 -24366
rect 5093 -24426 5353 -24366
rect 5413 -24426 5423 -24366
rect 5023 -24436 5423 -24426
rect 5481 -24366 5881 -24257
rect 5481 -24426 5491 -24366
rect 5551 -24426 5811 -24366
rect 5871 -24426 5881 -24366
rect 5481 -24436 5881 -24426
rect 5937 -24366 6337 -24257
rect 5937 -24426 5947 -24366
rect 6007 -24426 6267 -24366
rect 6327 -24426 6337 -24366
rect 5937 -24436 6337 -24426
rect 6393 -24366 6793 -24257
rect 6393 -24426 6403 -24366
rect 6463 -24426 6723 -24366
rect 6783 -24426 6793 -24366
rect 6393 -24436 6793 -24426
rect 6851 -24366 7251 -24257
rect 6851 -24426 6861 -24366
rect 6921 -24426 7181 -24366
rect 7241 -24426 7251 -24366
rect 6851 -24436 7251 -24426
rect 7307 -24366 7707 -24257
rect 7307 -24426 7317 -24366
rect 7377 -24426 7637 -24366
rect 7697 -24426 7707 -24366
rect 7307 -24436 7707 -24426
rect 7763 -24366 8163 -24257
rect 7763 -24426 7773 -24366
rect 7833 -24426 8093 -24366
rect 8153 -24426 8163 -24366
rect 7763 -24436 8163 -24426
rect 8237 -24366 8637 -24257
rect 8237 -24426 8247 -24366
rect 8307 -24426 8567 -24366
rect 8627 -24426 8637 -24366
rect 8237 -24436 8637 -24426
rect 8693 -24366 9093 -24257
rect 8693 -24426 8703 -24366
rect 8763 -24426 9023 -24366
rect 9083 -24426 9093 -24366
rect 8693 -24436 9093 -24426
rect 9151 -24366 9551 -24257
rect 9151 -24426 9161 -24366
rect 9221 -24426 9481 -24366
rect 9541 -24426 9551 -24366
rect 9151 -24436 9551 -24426
rect 9607 -24366 10007 -24257
rect 9607 -24426 9617 -24366
rect 9677 -24426 9937 -24366
rect 9997 -24426 10007 -24366
rect 9607 -24436 10007 -24426
rect 10063 -24366 10463 -24257
rect 10063 -24426 10073 -24366
rect 10133 -24426 10393 -24366
rect 10453 -24426 10463 -24366
rect 10063 -24436 10463 -24426
rect 10521 -24366 10921 -24257
rect 10521 -24426 10531 -24366
rect 10591 -24426 10851 -24366
rect 10911 -24426 10921 -24366
rect 10521 -24436 10921 -24426
rect 10977 -24366 11377 -24257
rect 10977 -24426 10987 -24366
rect 11047 -24426 11307 -24366
rect 11367 -24426 11377 -24366
rect 10977 -24436 11377 -24426
rect 11433 -24366 11833 -24257
rect 11433 -24426 11443 -24366
rect 11503 -24426 11763 -24366
rect 11823 -24426 11833 -24366
rect 11433 -24436 11833 -24426
rect 11891 -24366 12291 -24257
rect 11891 -24426 11901 -24366
rect 11961 -24426 12221 -24366
rect 12281 -24426 12291 -24366
rect 11891 -24436 12291 -24426
rect 12347 -24366 12747 -24257
rect 12347 -24426 12357 -24366
rect 12417 -24426 12677 -24366
rect 12737 -24426 12747 -24366
rect 12347 -24436 12747 -24426
rect 12803 -24366 13203 -24257
rect 12803 -24426 12813 -24366
rect 12873 -24426 13133 -24366
rect 13193 -24426 13203 -24366
rect 12803 -24436 13203 -24426
rect 13261 -24366 13661 -24257
rect 13261 -24426 13271 -24366
rect 13331 -24426 13591 -24366
rect 13651 -24426 13661 -24366
rect 13261 -24436 13661 -24426
rect 13717 -24366 14117 -24257
rect 13717 -24426 13727 -24366
rect 13787 -24426 14047 -24366
rect 14107 -24426 14117 -24366
rect 13717 -24436 14117 -24426
rect 14173 -24366 14573 -24257
rect 14173 -24426 14183 -24366
rect 14243 -24426 14503 -24366
rect 14563 -24426 14573 -24366
rect 14173 -24436 14573 -24426
rect 14631 -24366 15031 -24257
rect 14631 -24426 14641 -24366
rect 14701 -24426 14961 -24366
rect 15021 -24426 15031 -24366
rect 14631 -24436 15031 -24426
rect 15087 -24366 15487 -24257
rect 15087 -24426 15097 -24366
rect 15157 -24426 15417 -24366
rect 15477 -24426 15487 -24366
rect 15087 -24436 15487 -24426
rect 66 -24508 80 -24436
rect 457 -24508 527 -24436
rect 913 -24508 984 -24436
rect 1371 -24508 1442 -24436
rect 1827 -24508 1898 -24436
rect 2283 -24508 2354 -24436
rect 2741 -24508 2812 -24436
rect 3197 -24508 3268 -24436
rect 3653 -24508 3724 -24436
rect 4111 -24508 4182 -24436
rect 4567 -24508 4638 -24436
rect 5023 -24508 5094 -24436
rect 5481 -24508 5552 -24436
rect 5937 -24508 6008 -24436
rect 6393 -24508 6464 -24436
rect 6851 -24508 6922 -24436
rect 7307 -24508 7378 -24436
rect 7763 -24508 7834 -24436
rect 8237 -24508 8308 -24436
rect 8693 -24508 8764 -24436
rect 9151 -24508 9222 -24436
rect 9607 -24508 9678 -24436
rect 10063 -24508 10134 -24436
rect 10521 -24508 10592 -24436
rect 10977 -24508 11048 -24436
rect 11433 -24508 11504 -24436
rect 11891 -24508 11962 -24436
rect 12347 -24508 12418 -24436
rect 12803 -24508 12874 -24436
rect 13261 -24508 13332 -24436
rect 13717 -24508 13788 -24436
rect 14173 -24508 14244 -24436
rect 14631 -24508 14702 -24436
rect 66 -24518 400 -24508
rect 0 -24578 11 -24518
rect 71 -24578 331 -24518
rect 391 -24578 400 -24518
rect 0 -24868 14 -24578
rect 66 -24868 400 -24578
rect 0 -24928 11 -24868
rect 71 -24928 331 -24868
rect 391 -24928 400 -24868
rect 0 -25034 14 -24928
rect 66 -24938 400 -24928
rect 457 -24518 857 -24508
rect 457 -24578 467 -24518
rect 527 -24578 787 -24518
rect 847 -24578 857 -24518
rect 457 -24688 857 -24578
rect 913 -24518 1313 -24508
rect 913 -24578 923 -24518
rect 983 -24578 1243 -24518
rect 1303 -24578 1313 -24518
rect 913 -24688 1313 -24578
rect 1371 -24518 1771 -24508
rect 1371 -24578 1381 -24518
rect 1441 -24578 1701 -24518
rect 1761 -24578 1771 -24518
rect 1371 -24688 1771 -24578
rect 1827 -24518 2227 -24508
rect 1827 -24578 1837 -24518
rect 1897 -24578 2157 -24518
rect 2217 -24578 2227 -24518
rect 1827 -24688 2227 -24578
rect 2283 -24518 2683 -24508
rect 2283 -24578 2293 -24518
rect 2353 -24578 2613 -24518
rect 2673 -24578 2683 -24518
rect 2283 -24688 2683 -24578
rect 457 -24689 2683 -24688
rect 2741 -24518 3141 -24508
rect 2741 -24578 2751 -24518
rect 2811 -24578 3071 -24518
rect 3131 -24578 3141 -24518
rect 2741 -24688 3141 -24578
rect 3197 -24518 3597 -24508
rect 3197 -24578 3207 -24518
rect 3267 -24578 3527 -24518
rect 3587 -24578 3597 -24518
rect 3197 -24688 3597 -24578
rect 3653 -24518 4053 -24508
rect 3653 -24578 3663 -24518
rect 3723 -24578 3983 -24518
rect 4043 -24578 4053 -24518
rect 3653 -24688 4053 -24578
rect 2741 -24689 4053 -24688
rect 457 -24759 4053 -24689
rect 457 -24868 857 -24759
rect 457 -24928 467 -24868
rect 527 -24928 787 -24868
rect 847 -24928 857 -24868
rect 457 -24938 857 -24928
rect 913 -24868 1313 -24759
rect 913 -24928 923 -24868
rect 983 -24928 1243 -24868
rect 1303 -24928 1313 -24868
rect 913 -24938 1313 -24928
rect 1371 -24868 1771 -24759
rect 1371 -24928 1381 -24868
rect 1441 -24928 1701 -24868
rect 1761 -24928 1771 -24868
rect 1371 -24938 1771 -24928
rect 1827 -24868 2227 -24759
rect 1827 -24928 1837 -24868
rect 1897 -24928 2157 -24868
rect 2217 -24928 2227 -24868
rect 1827 -24938 2227 -24928
rect 2283 -24868 2683 -24759
rect 2283 -24928 2293 -24868
rect 2353 -24928 2613 -24868
rect 2673 -24928 2683 -24868
rect 2283 -24938 2683 -24928
rect 2741 -24868 3141 -24759
rect 2741 -24928 2751 -24868
rect 2811 -24928 3071 -24868
rect 3131 -24928 3141 -24868
rect 2741 -24938 3141 -24928
rect 3197 -24868 3597 -24759
rect 3197 -24928 3207 -24868
rect 3267 -24928 3527 -24868
rect 3587 -24928 3597 -24868
rect 3197 -24938 3597 -24928
rect 3653 -24868 4053 -24759
rect 3653 -24928 3663 -24868
rect 3723 -24928 3983 -24868
rect 4043 -24928 4053 -24868
rect 3653 -24938 4053 -24928
rect 4111 -24518 4511 -24508
rect 4111 -24578 4121 -24518
rect 4181 -24578 4441 -24518
rect 4501 -24578 4511 -24518
rect 4111 -24688 4511 -24578
rect 4567 -24518 4967 -24508
rect 4567 -24578 4577 -24518
rect 4637 -24578 4897 -24518
rect 4957 -24578 4967 -24518
rect 4567 -24688 4967 -24578
rect 5023 -24518 5423 -24508
rect 5023 -24578 5033 -24518
rect 5093 -24578 5353 -24518
rect 5413 -24578 5423 -24518
rect 5023 -24688 5423 -24578
rect 5481 -24518 5881 -24508
rect 5481 -24578 5491 -24518
rect 5551 -24578 5811 -24518
rect 5871 -24578 5881 -24518
rect 5481 -24688 5881 -24578
rect 5937 -24518 6337 -24508
rect 5937 -24578 5947 -24518
rect 6007 -24578 6267 -24518
rect 6327 -24578 6337 -24518
rect 5937 -24688 6337 -24578
rect 6393 -24518 6793 -24508
rect 6393 -24578 6403 -24518
rect 6463 -24578 6723 -24518
rect 6783 -24578 6793 -24518
rect 6393 -24688 6793 -24578
rect 6851 -24518 7251 -24508
rect 6851 -24578 6861 -24518
rect 6921 -24578 7181 -24518
rect 7241 -24578 7251 -24518
rect 6851 -24688 7251 -24578
rect 7307 -24518 7707 -24508
rect 7307 -24578 7317 -24518
rect 7377 -24578 7637 -24518
rect 7697 -24578 7707 -24518
rect 7307 -24688 7707 -24578
rect 7763 -24518 8163 -24508
rect 7763 -24578 7773 -24518
rect 7833 -24578 8093 -24518
rect 8153 -24578 8163 -24518
rect 7763 -24688 8163 -24578
rect 8237 -24518 8637 -24508
rect 8237 -24578 8247 -24518
rect 8307 -24578 8567 -24518
rect 8627 -24578 8637 -24518
rect 8237 -24688 8637 -24578
rect 8693 -24518 9093 -24508
rect 8693 -24578 8703 -24518
rect 8763 -24578 9023 -24518
rect 9083 -24578 9093 -24518
rect 8693 -24688 9093 -24578
rect 9151 -24518 9551 -24508
rect 9151 -24578 9161 -24518
rect 9221 -24578 9481 -24518
rect 9541 -24578 9551 -24518
rect 9151 -24688 9551 -24578
rect 9607 -24518 10007 -24508
rect 9607 -24578 9617 -24518
rect 9677 -24578 9937 -24518
rect 9997 -24578 10007 -24518
rect 9607 -24688 10007 -24578
rect 10063 -24518 10463 -24508
rect 10063 -24578 10073 -24518
rect 10133 -24578 10393 -24518
rect 10453 -24578 10463 -24518
rect 10063 -24688 10463 -24578
rect 4111 -24689 10463 -24688
rect 10521 -24518 10921 -24508
rect 10521 -24578 10531 -24518
rect 10591 -24578 10851 -24518
rect 10911 -24578 10921 -24518
rect 10521 -24688 10921 -24578
rect 10977 -24518 11377 -24508
rect 10977 -24578 10987 -24518
rect 11047 -24578 11307 -24518
rect 11367 -24578 11377 -24518
rect 10977 -24688 11377 -24578
rect 11433 -24518 11833 -24508
rect 11433 -24578 11443 -24518
rect 11503 -24578 11763 -24518
rect 11823 -24578 11833 -24518
rect 11433 -24688 11833 -24578
rect 11891 -24518 12291 -24508
rect 11891 -24578 11901 -24518
rect 11961 -24578 12221 -24518
rect 12281 -24578 12291 -24518
rect 11891 -24688 12291 -24578
rect 12347 -24518 12747 -24508
rect 12347 -24578 12357 -24518
rect 12417 -24578 12677 -24518
rect 12737 -24578 12747 -24518
rect 12347 -24688 12747 -24578
rect 12803 -24518 13203 -24508
rect 12803 -24578 12813 -24518
rect 12873 -24578 13133 -24518
rect 13193 -24578 13203 -24518
rect 12803 -24688 13203 -24578
rect 13261 -24518 13661 -24508
rect 13261 -24578 13271 -24518
rect 13331 -24578 13591 -24518
rect 13651 -24578 13661 -24518
rect 13261 -24688 13661 -24578
rect 13717 -24518 14117 -24508
rect 13717 -24578 13727 -24518
rect 13787 -24578 14047 -24518
rect 14107 -24578 14117 -24518
rect 13717 -24688 14117 -24578
rect 14173 -24518 14573 -24508
rect 14173 -24578 14183 -24518
rect 14243 -24578 14503 -24518
rect 14563 -24578 14573 -24518
rect 14173 -24688 14573 -24578
rect 14631 -24518 15031 -24508
rect 14631 -24578 14641 -24518
rect 14701 -24578 14961 -24518
rect 15021 -24578 15031 -24518
rect 14631 -24688 15031 -24578
rect 15087 -24518 15487 -24508
rect 15087 -24578 15097 -24518
rect 15157 -24578 15417 -24518
rect 15477 -24578 15487 -24518
rect 15087 -24688 15487 -24578
rect 10521 -24689 15487 -24688
rect 4111 -24759 15487 -24689
rect 4111 -24868 4511 -24759
rect 4111 -24928 4121 -24868
rect 4181 -24928 4441 -24868
rect 4501 -24928 4511 -24868
rect 4111 -24938 4511 -24928
rect 4567 -24868 4967 -24759
rect 4567 -24928 4577 -24868
rect 4637 -24928 4897 -24868
rect 4957 -24928 4967 -24868
rect 4567 -24938 4967 -24928
rect 5023 -24868 5423 -24759
rect 5023 -24928 5033 -24868
rect 5093 -24928 5353 -24868
rect 5413 -24928 5423 -24868
rect 5023 -24938 5423 -24928
rect 5481 -24868 5881 -24759
rect 5481 -24928 5491 -24868
rect 5551 -24928 5811 -24868
rect 5871 -24928 5881 -24868
rect 5481 -24938 5881 -24928
rect 5937 -24868 6337 -24759
rect 5937 -24928 5947 -24868
rect 6007 -24928 6267 -24868
rect 6327 -24928 6337 -24868
rect 5937 -24938 6337 -24928
rect 6393 -24868 6793 -24759
rect 6393 -24928 6403 -24868
rect 6463 -24928 6723 -24868
rect 6783 -24928 6793 -24868
rect 6393 -24938 6793 -24928
rect 6851 -24868 7251 -24759
rect 6851 -24928 6861 -24868
rect 6921 -24928 7181 -24868
rect 7241 -24928 7251 -24868
rect 6851 -24938 7251 -24928
rect 7307 -24868 7707 -24759
rect 7307 -24928 7317 -24868
rect 7377 -24928 7637 -24868
rect 7697 -24928 7707 -24868
rect 7307 -24938 7707 -24928
rect 7763 -24868 8163 -24759
rect 7763 -24928 7773 -24868
rect 7833 -24928 8093 -24868
rect 8153 -24928 8163 -24868
rect 7763 -24938 8163 -24928
rect 8237 -24868 8637 -24759
rect 8237 -24928 8247 -24868
rect 8307 -24928 8567 -24868
rect 8627 -24928 8637 -24868
rect 8237 -24938 8637 -24928
rect 8693 -24868 9093 -24759
rect 8693 -24928 8703 -24868
rect 8763 -24928 9023 -24868
rect 9083 -24928 9093 -24868
rect 8693 -24938 9093 -24928
rect 9151 -24868 9551 -24759
rect 9151 -24928 9161 -24868
rect 9221 -24928 9481 -24868
rect 9541 -24928 9551 -24868
rect 9151 -24938 9551 -24928
rect 9607 -24868 10007 -24759
rect 9607 -24928 9617 -24868
rect 9677 -24928 9937 -24868
rect 9997 -24928 10007 -24868
rect 9607 -24938 10007 -24928
rect 10063 -24868 10463 -24759
rect 10063 -24928 10073 -24868
rect 10133 -24928 10393 -24868
rect 10453 -24928 10463 -24868
rect 10063 -24938 10463 -24928
rect 10521 -24868 10921 -24759
rect 10521 -24928 10531 -24868
rect 10591 -24928 10851 -24868
rect 10911 -24928 10921 -24868
rect 10521 -24938 10921 -24928
rect 10977 -24868 11377 -24759
rect 10977 -24928 10987 -24868
rect 11047 -24928 11307 -24868
rect 11367 -24928 11377 -24868
rect 10977 -24938 11377 -24928
rect 11433 -24868 11833 -24759
rect 11433 -24928 11443 -24868
rect 11503 -24928 11763 -24868
rect 11823 -24928 11833 -24868
rect 11433 -24938 11833 -24928
rect 11891 -24868 12291 -24759
rect 11891 -24928 11901 -24868
rect 11961 -24928 12221 -24868
rect 12281 -24928 12291 -24868
rect 11891 -24938 12291 -24928
rect 12347 -24868 12747 -24759
rect 12347 -24928 12357 -24868
rect 12417 -24928 12677 -24868
rect 12737 -24928 12747 -24868
rect 12347 -24938 12747 -24928
rect 12803 -24868 13203 -24759
rect 12803 -24928 12813 -24868
rect 12873 -24928 13133 -24868
rect 13193 -24928 13203 -24868
rect 12803 -24938 13203 -24928
rect 13261 -24868 13661 -24759
rect 13261 -24928 13271 -24868
rect 13331 -24928 13591 -24868
rect 13651 -24928 13661 -24868
rect 13261 -24938 13661 -24928
rect 13717 -24868 14117 -24759
rect 13717 -24928 13727 -24868
rect 13787 -24928 14047 -24868
rect 14107 -24928 14117 -24868
rect 13717 -24938 14117 -24928
rect 14173 -24868 14573 -24759
rect 14173 -24928 14183 -24868
rect 14243 -24928 14503 -24868
rect 14563 -24928 14573 -24868
rect 14173 -24938 14573 -24928
rect 14631 -24868 15031 -24759
rect 14631 -24928 14641 -24868
rect 14701 -24928 14961 -24868
rect 15021 -24928 15031 -24868
rect 14631 -24938 15031 -24928
rect 15087 -24868 15487 -24759
rect 15087 -24928 15097 -24868
rect 15157 -24928 15417 -24868
rect 15477 -24928 15487 -24868
rect 15087 -24938 15487 -24928
rect 66 -25024 80 -24938
rect 457 -25024 527 -24938
rect 913 -25024 983 -24938
rect 1371 -25024 1441 -24938
rect 1827 -25024 1897 -24938
rect 2283 -25024 2353 -24938
rect 2741 -25024 2811 -24938
rect 3197 -25024 3267 -24938
rect 3653 -25024 3723 -24938
rect 4111 -25024 4181 -24938
rect 4567 -25024 4637 -24938
rect 5023 -25024 5093 -24938
rect 5481 -25024 5551 -24938
rect 5937 -25024 6007 -24938
rect 6393 -25024 6463 -24938
rect 6851 -25024 6921 -24938
rect 7307 -25024 7377 -24938
rect 7763 -25024 7833 -24938
rect 8237 -25024 8307 -24938
rect 8693 -25024 8763 -24938
rect 9151 -25024 9221 -24938
rect 9607 -25024 9677 -24938
rect 10063 -25024 10133 -24938
rect 10521 -25024 10591 -24938
rect 10977 -25024 11047 -24938
rect 11433 -25024 11503 -24938
rect 11891 -25024 11961 -24938
rect 12347 -25024 12417 -24938
rect 12803 -25024 12873 -24938
rect 13261 -25024 13331 -24938
rect 13717 -25024 13787 -24938
rect 14173 -25024 14243 -24938
rect 14631 -25024 14701 -24938
rect 66 -25034 400 -25024
rect 0 -25094 11 -25034
rect 71 -25094 331 -25034
rect 391 -25094 400 -25034
rect 0 -25384 14 -25094
rect 66 -25384 400 -25094
rect 0 -25444 11 -25384
rect 71 -25444 331 -25384
rect 391 -25444 400 -25384
rect 0 -25526 14 -25444
rect 66 -25454 400 -25444
rect 457 -25034 857 -25024
rect 457 -25094 467 -25034
rect 527 -25094 787 -25034
rect 847 -25094 857 -25034
rect 457 -25203 857 -25094
rect 913 -25034 1313 -25024
rect 913 -25094 923 -25034
rect 983 -25094 1243 -25034
rect 1303 -25094 1313 -25034
rect 913 -25203 1313 -25094
rect 1371 -25034 1771 -25024
rect 1371 -25094 1381 -25034
rect 1441 -25094 1701 -25034
rect 1761 -25094 1771 -25034
rect 1371 -25203 1771 -25094
rect 1827 -25034 2227 -25024
rect 1827 -25094 1837 -25034
rect 1897 -25094 2157 -25034
rect 2217 -25094 2227 -25034
rect 1827 -25203 2227 -25094
rect 2283 -25034 2683 -25024
rect 2283 -25094 2293 -25034
rect 2353 -25094 2613 -25034
rect 2673 -25094 2683 -25034
rect 2283 -25203 2683 -25094
rect 2741 -25034 3141 -25024
rect 2741 -25094 2751 -25034
rect 2811 -25094 3071 -25034
rect 3131 -25094 3141 -25034
rect 2741 -25203 3141 -25094
rect 3197 -25034 3597 -25024
rect 3197 -25094 3207 -25034
rect 3267 -25094 3527 -25034
rect 3587 -25094 3597 -25034
rect 3197 -25203 3597 -25094
rect 3653 -25034 4053 -25024
rect 3653 -25094 3663 -25034
rect 3723 -25094 3983 -25034
rect 4043 -25094 4053 -25034
rect 3653 -25203 4053 -25094
rect 457 -25273 4053 -25203
rect 457 -25274 2683 -25273
rect 457 -25384 857 -25274
rect 457 -25444 467 -25384
rect 527 -25444 787 -25384
rect 847 -25444 857 -25384
rect 457 -25454 857 -25444
rect 913 -25384 1313 -25274
rect 913 -25444 923 -25384
rect 983 -25444 1243 -25384
rect 1303 -25444 1313 -25384
rect 913 -25454 1313 -25444
rect 1371 -25384 1771 -25274
rect 1371 -25444 1381 -25384
rect 1441 -25444 1701 -25384
rect 1761 -25444 1771 -25384
rect 1371 -25454 1771 -25444
rect 1827 -25384 2227 -25274
rect 1827 -25444 1837 -25384
rect 1897 -25444 2157 -25384
rect 2217 -25444 2227 -25384
rect 1827 -25454 2227 -25444
rect 2283 -25384 2683 -25274
rect 2283 -25444 2293 -25384
rect 2353 -25444 2613 -25384
rect 2673 -25444 2683 -25384
rect 2283 -25454 2683 -25444
rect 2741 -25274 4053 -25273
rect 2741 -25384 3141 -25274
rect 2741 -25444 2751 -25384
rect 2811 -25444 3071 -25384
rect 3131 -25444 3141 -25384
rect 2741 -25454 3141 -25444
rect 3197 -25384 3597 -25274
rect 3197 -25444 3207 -25384
rect 3267 -25444 3527 -25384
rect 3587 -25444 3597 -25384
rect 3197 -25454 3597 -25444
rect 3653 -25384 4053 -25274
rect 3653 -25444 3663 -25384
rect 3723 -25444 3983 -25384
rect 4043 -25444 4053 -25384
rect 3653 -25454 4053 -25444
rect 4111 -25034 4511 -25024
rect 4111 -25094 4121 -25034
rect 4181 -25094 4441 -25034
rect 4501 -25094 4511 -25034
rect 4111 -25203 4511 -25094
rect 4567 -25034 4967 -25024
rect 4567 -25094 4577 -25034
rect 4637 -25094 4897 -25034
rect 4957 -25094 4967 -25034
rect 4567 -25203 4967 -25094
rect 5023 -25034 5423 -25024
rect 5023 -25094 5033 -25034
rect 5093 -25094 5353 -25034
rect 5413 -25094 5423 -25034
rect 5023 -25203 5423 -25094
rect 5481 -25034 5881 -25024
rect 5481 -25094 5491 -25034
rect 5551 -25094 5811 -25034
rect 5871 -25094 5881 -25034
rect 5481 -25203 5881 -25094
rect 5937 -25034 6337 -25024
rect 5937 -25094 5947 -25034
rect 6007 -25094 6267 -25034
rect 6327 -25094 6337 -25034
rect 5937 -25203 6337 -25094
rect 6393 -25034 6793 -25024
rect 6393 -25094 6403 -25034
rect 6463 -25094 6723 -25034
rect 6783 -25094 6793 -25034
rect 6393 -25203 6793 -25094
rect 6851 -25034 7251 -25024
rect 6851 -25094 6861 -25034
rect 6921 -25094 7181 -25034
rect 7241 -25094 7251 -25034
rect 6851 -25203 7251 -25094
rect 7307 -25034 7707 -25024
rect 7307 -25094 7317 -25034
rect 7377 -25094 7637 -25034
rect 7697 -25094 7707 -25034
rect 7307 -25203 7707 -25094
rect 7763 -25034 8163 -25024
rect 7763 -25094 7773 -25034
rect 7833 -25094 8093 -25034
rect 8153 -25094 8163 -25034
rect 7763 -25203 8163 -25094
rect 8237 -25034 8637 -25024
rect 8237 -25094 8247 -25034
rect 8307 -25094 8567 -25034
rect 8627 -25094 8637 -25034
rect 8237 -25203 8637 -25094
rect 8693 -25034 9093 -25024
rect 8693 -25094 8703 -25034
rect 8763 -25094 9023 -25034
rect 9083 -25094 9093 -25034
rect 8693 -25203 9093 -25094
rect 9151 -25034 9551 -25024
rect 9151 -25094 9161 -25034
rect 9221 -25094 9481 -25034
rect 9541 -25094 9551 -25034
rect 9151 -25203 9551 -25094
rect 9607 -25034 10007 -25024
rect 9607 -25094 9617 -25034
rect 9677 -25094 9937 -25034
rect 9997 -25094 10007 -25034
rect 9607 -25203 10007 -25094
rect 10063 -25034 10463 -25024
rect 10063 -25094 10073 -25034
rect 10133 -25094 10393 -25034
rect 10453 -25094 10463 -25034
rect 10063 -25203 10463 -25094
rect 10521 -25034 10921 -25024
rect 10521 -25094 10531 -25034
rect 10591 -25094 10851 -25034
rect 10911 -25094 10921 -25034
rect 10521 -25203 10921 -25094
rect 10977 -25034 11377 -25024
rect 10977 -25094 10987 -25034
rect 11047 -25094 11307 -25034
rect 11367 -25094 11377 -25034
rect 10977 -25203 11377 -25094
rect 11433 -25034 11833 -25024
rect 11433 -25094 11443 -25034
rect 11503 -25094 11763 -25034
rect 11823 -25094 11833 -25034
rect 11433 -25203 11833 -25094
rect 11891 -25034 12291 -25024
rect 11891 -25094 11901 -25034
rect 11961 -25094 12221 -25034
rect 12281 -25094 12291 -25034
rect 11891 -25203 12291 -25094
rect 12347 -25034 12747 -25024
rect 12347 -25094 12357 -25034
rect 12417 -25094 12677 -25034
rect 12737 -25094 12747 -25034
rect 12347 -25203 12747 -25094
rect 12803 -25034 13203 -25024
rect 12803 -25094 12813 -25034
rect 12873 -25094 13133 -25034
rect 13193 -25094 13203 -25034
rect 12803 -25203 13203 -25094
rect 13261 -25034 13661 -25024
rect 13261 -25094 13271 -25034
rect 13331 -25094 13591 -25034
rect 13651 -25094 13661 -25034
rect 13261 -25203 13661 -25094
rect 13717 -25034 14117 -25024
rect 13717 -25094 13727 -25034
rect 13787 -25094 14047 -25034
rect 14107 -25094 14117 -25034
rect 13717 -25203 14117 -25094
rect 14173 -25034 14573 -25024
rect 14173 -25094 14183 -25034
rect 14243 -25094 14503 -25034
rect 14563 -25094 14573 -25034
rect 14173 -25203 14573 -25094
rect 14631 -25034 15031 -25024
rect 14631 -25094 14641 -25034
rect 14701 -25094 14961 -25034
rect 15021 -25094 15031 -25034
rect 14631 -25203 15031 -25094
rect 15087 -25034 15487 -25024
rect 15087 -25094 15097 -25034
rect 15157 -25094 15417 -25034
rect 15477 -25094 15487 -25034
rect 15087 -25203 15487 -25094
rect 4111 -25273 15487 -25203
rect 4111 -25274 10463 -25273
rect 4111 -25384 4511 -25274
rect 4111 -25444 4121 -25384
rect 4181 -25444 4441 -25384
rect 4501 -25444 4511 -25384
rect 4111 -25454 4511 -25444
rect 4567 -25384 4967 -25274
rect 4567 -25444 4577 -25384
rect 4637 -25444 4897 -25384
rect 4957 -25444 4967 -25384
rect 4567 -25454 4967 -25444
rect 5023 -25384 5423 -25274
rect 5023 -25444 5033 -25384
rect 5093 -25444 5353 -25384
rect 5413 -25444 5423 -25384
rect 5023 -25454 5423 -25444
rect 5481 -25384 5881 -25274
rect 5481 -25444 5491 -25384
rect 5551 -25444 5811 -25384
rect 5871 -25444 5881 -25384
rect 5481 -25454 5881 -25444
rect 5937 -25384 6337 -25274
rect 5937 -25444 5947 -25384
rect 6007 -25444 6267 -25384
rect 6327 -25444 6337 -25384
rect 5937 -25454 6337 -25444
rect 6393 -25384 6793 -25274
rect 6393 -25444 6403 -25384
rect 6463 -25444 6723 -25384
rect 6783 -25444 6793 -25384
rect 6393 -25454 6793 -25444
rect 6851 -25384 7251 -25274
rect 6851 -25444 6861 -25384
rect 6921 -25444 7181 -25384
rect 7241 -25444 7251 -25384
rect 6851 -25454 7251 -25444
rect 7307 -25384 7707 -25274
rect 7307 -25444 7317 -25384
rect 7377 -25444 7637 -25384
rect 7697 -25444 7707 -25384
rect 7307 -25454 7707 -25444
rect 7763 -25384 8163 -25274
rect 7763 -25444 7773 -25384
rect 7833 -25444 8093 -25384
rect 8153 -25444 8163 -25384
rect 7763 -25454 8163 -25444
rect 8237 -25384 8637 -25274
rect 8237 -25444 8247 -25384
rect 8307 -25444 8567 -25384
rect 8627 -25444 8637 -25384
rect 8237 -25454 8637 -25444
rect 8693 -25384 9093 -25274
rect 8693 -25444 8703 -25384
rect 8763 -25444 9023 -25384
rect 9083 -25444 9093 -25384
rect 8693 -25454 9093 -25444
rect 9151 -25384 9551 -25274
rect 9151 -25444 9161 -25384
rect 9221 -25444 9481 -25384
rect 9541 -25444 9551 -25384
rect 9151 -25454 9551 -25444
rect 9607 -25384 10007 -25274
rect 9607 -25444 9617 -25384
rect 9677 -25444 9937 -25384
rect 9997 -25444 10007 -25384
rect 9607 -25454 10007 -25444
rect 10063 -25384 10463 -25274
rect 10063 -25444 10073 -25384
rect 10133 -25444 10393 -25384
rect 10453 -25444 10463 -25384
rect 10063 -25454 10463 -25444
rect 10521 -25274 15487 -25273
rect 10521 -25384 10921 -25274
rect 10521 -25444 10531 -25384
rect 10591 -25444 10851 -25384
rect 10911 -25444 10921 -25384
rect 10521 -25454 10921 -25444
rect 10977 -25384 11377 -25274
rect 10977 -25444 10987 -25384
rect 11047 -25444 11307 -25384
rect 11367 -25444 11377 -25384
rect 10977 -25454 11377 -25444
rect 11433 -25384 11833 -25274
rect 11433 -25444 11443 -25384
rect 11503 -25444 11763 -25384
rect 11823 -25444 11833 -25384
rect 11433 -25454 11833 -25444
rect 11891 -25384 12291 -25274
rect 11891 -25444 11901 -25384
rect 11961 -25444 12221 -25384
rect 12281 -25444 12291 -25384
rect 11891 -25454 12291 -25444
rect 12347 -25384 12747 -25274
rect 12347 -25444 12357 -25384
rect 12417 -25444 12677 -25384
rect 12737 -25444 12747 -25384
rect 12347 -25454 12747 -25444
rect 12803 -25384 13203 -25274
rect 12803 -25444 12813 -25384
rect 12873 -25444 13133 -25384
rect 13193 -25444 13203 -25384
rect 12803 -25454 13203 -25444
rect 13261 -25384 13661 -25274
rect 13261 -25444 13271 -25384
rect 13331 -25444 13591 -25384
rect 13651 -25444 13661 -25384
rect 13261 -25454 13661 -25444
rect 13717 -25384 14117 -25274
rect 13717 -25444 13727 -25384
rect 13787 -25444 14047 -25384
rect 14107 -25444 14117 -25384
rect 13717 -25454 14117 -25444
rect 14173 -25384 14573 -25274
rect 14173 -25444 14183 -25384
rect 14243 -25444 14503 -25384
rect 14563 -25444 14573 -25384
rect 14173 -25454 14573 -25444
rect 14631 -25384 15031 -25274
rect 14631 -25444 14641 -25384
rect 14701 -25444 14961 -25384
rect 15021 -25444 15031 -25384
rect 14631 -25454 15031 -25444
rect 15087 -25384 15487 -25274
rect 15087 -25444 15097 -25384
rect 15157 -25444 15417 -25384
rect 15477 -25444 15487 -25384
rect 15087 -25454 15487 -25444
rect 66 -25516 80 -25454
rect 457 -25516 528 -25454
rect 913 -25516 984 -25454
rect 1371 -25516 1442 -25454
rect 1827 -25516 1898 -25454
rect 2283 -25516 2354 -25454
rect 2741 -25516 2811 -25454
rect 3197 -25516 3267 -25454
rect 3653 -25516 3723 -25454
rect 4111 -25516 4181 -25454
rect 4567 -25516 4637 -25454
rect 5023 -25516 5093 -25454
rect 5481 -25516 5551 -25454
rect 5937 -25516 6007 -25454
rect 6393 -25516 6463 -25454
rect 6851 -25516 6921 -25454
rect 7307 -25516 7377 -25454
rect 7763 -25516 7833 -25454
rect 8237 -25516 8307 -25454
rect 8693 -25516 8763 -25454
rect 9151 -25516 9221 -25454
rect 9607 -25516 9677 -25454
rect 10063 -25516 10133 -25454
rect 10521 -25516 10591 -25454
rect 10977 -25516 11047 -25454
rect 11433 -25516 11503 -25454
rect 11891 -25516 11961 -25454
rect 12347 -25516 12417 -25454
rect 12803 -25516 12873 -25454
rect 13261 -25516 13331 -25454
rect 13717 -25516 13787 -25454
rect 14173 -25516 14243 -25454
rect 14631 -25516 14701 -25454
rect 66 -25526 400 -25516
rect 0 -25586 11 -25526
rect 71 -25586 331 -25526
rect 391 -25586 400 -25526
rect 0 -25876 14 -25586
rect 66 -25876 400 -25586
rect 0 -25936 11 -25876
rect 71 -25936 331 -25876
rect 391 -25936 400 -25876
rect 0 -26023 14 -25936
rect 66 -25946 400 -25936
rect 457 -25526 857 -25516
rect 457 -25586 467 -25526
rect 527 -25586 787 -25526
rect 847 -25586 857 -25526
rect 457 -25696 857 -25586
rect 913 -25526 1313 -25516
rect 913 -25586 923 -25526
rect 983 -25586 1243 -25526
rect 1303 -25586 1313 -25526
rect 913 -25696 1313 -25586
rect 1371 -25526 1771 -25516
rect 1371 -25586 1381 -25526
rect 1441 -25586 1701 -25526
rect 1761 -25586 1771 -25526
rect 1371 -25696 1771 -25586
rect 1827 -25526 2227 -25516
rect 1827 -25586 1837 -25526
rect 1897 -25586 2157 -25526
rect 2217 -25586 2227 -25526
rect 1827 -25696 2227 -25586
rect 2283 -25526 2683 -25516
rect 2283 -25586 2293 -25526
rect 2353 -25586 2613 -25526
rect 2673 -25586 2683 -25526
rect 2283 -25696 2683 -25586
rect 2741 -25526 3141 -25516
rect 2741 -25586 2751 -25526
rect 2811 -25586 3071 -25526
rect 3131 -25586 3141 -25526
rect 2741 -25696 3141 -25586
rect 3197 -25526 3597 -25516
rect 3197 -25586 3207 -25526
rect 3267 -25586 3527 -25526
rect 3587 -25586 3597 -25526
rect 3197 -25696 3597 -25586
rect 3653 -25526 4053 -25516
rect 3653 -25586 3663 -25526
rect 3723 -25586 3983 -25526
rect 4043 -25586 4053 -25526
rect 3653 -25696 4053 -25586
rect 457 -25766 4053 -25696
rect 457 -25876 857 -25766
rect 457 -25936 467 -25876
rect 527 -25936 787 -25876
rect 847 -25936 857 -25876
rect 457 -25946 857 -25936
rect 913 -25876 1313 -25766
rect 913 -25936 923 -25876
rect 983 -25936 1243 -25876
rect 1303 -25936 1313 -25876
rect 913 -25946 1313 -25936
rect 1371 -25876 1771 -25766
rect 1371 -25936 1381 -25876
rect 1441 -25936 1701 -25876
rect 1761 -25936 1771 -25876
rect 1371 -25946 1771 -25936
rect 1827 -25876 2227 -25766
rect 1827 -25936 1837 -25876
rect 1897 -25936 2157 -25876
rect 2217 -25936 2227 -25876
rect 1827 -25946 2227 -25936
rect 2283 -25876 2683 -25766
rect 2283 -25936 2293 -25876
rect 2353 -25936 2613 -25876
rect 2673 -25936 2683 -25876
rect 2283 -25946 2683 -25936
rect 2741 -25876 3141 -25766
rect 2741 -25936 2751 -25876
rect 2811 -25936 3071 -25876
rect 3131 -25936 3141 -25876
rect 2741 -25946 3141 -25936
rect 3197 -25876 3597 -25766
rect 3197 -25936 3207 -25876
rect 3267 -25936 3527 -25876
rect 3587 -25936 3597 -25876
rect 3197 -25946 3597 -25936
rect 3653 -25876 4053 -25766
rect 3653 -25936 3663 -25876
rect 3723 -25936 3983 -25876
rect 4043 -25936 4053 -25876
rect 3653 -25946 4053 -25936
rect 4111 -25526 4511 -25516
rect 4111 -25586 4121 -25526
rect 4181 -25586 4441 -25526
rect 4501 -25586 4511 -25526
rect 4111 -25696 4511 -25586
rect 4567 -25526 4967 -25516
rect 4567 -25586 4577 -25526
rect 4637 -25586 4897 -25526
rect 4957 -25586 4967 -25526
rect 4567 -25696 4967 -25586
rect 5023 -25526 5423 -25516
rect 5023 -25586 5033 -25526
rect 5093 -25586 5353 -25526
rect 5413 -25586 5423 -25526
rect 5023 -25696 5423 -25586
rect 5481 -25526 5881 -25516
rect 5481 -25586 5491 -25526
rect 5551 -25586 5811 -25526
rect 5871 -25586 5881 -25526
rect 5481 -25696 5881 -25586
rect 5937 -25526 6337 -25516
rect 5937 -25586 5947 -25526
rect 6007 -25586 6267 -25526
rect 6327 -25586 6337 -25526
rect 5937 -25696 6337 -25586
rect 6393 -25526 6793 -25516
rect 6393 -25586 6403 -25526
rect 6463 -25586 6723 -25526
rect 6783 -25586 6793 -25526
rect 6393 -25696 6793 -25586
rect 6851 -25526 7251 -25516
rect 6851 -25586 6861 -25526
rect 6921 -25586 7181 -25526
rect 7241 -25586 7251 -25526
rect 6851 -25696 7251 -25586
rect 7307 -25526 7707 -25516
rect 7307 -25586 7317 -25526
rect 7377 -25586 7637 -25526
rect 7697 -25586 7707 -25526
rect 7307 -25696 7707 -25586
rect 7763 -25526 8163 -25516
rect 7763 -25586 7773 -25526
rect 7833 -25586 8093 -25526
rect 8153 -25586 8163 -25526
rect 7763 -25696 8163 -25586
rect 8237 -25526 8637 -25516
rect 8237 -25586 8247 -25526
rect 8307 -25586 8567 -25526
rect 8627 -25586 8637 -25526
rect 8237 -25696 8637 -25586
rect 8693 -25526 9093 -25516
rect 8693 -25586 8703 -25526
rect 8763 -25586 9023 -25526
rect 9083 -25586 9093 -25526
rect 8693 -25696 9093 -25586
rect 9151 -25526 9551 -25516
rect 9151 -25586 9161 -25526
rect 9221 -25586 9481 -25526
rect 9541 -25586 9551 -25526
rect 9151 -25696 9551 -25586
rect 9607 -25526 10007 -25516
rect 9607 -25586 9617 -25526
rect 9677 -25586 9937 -25526
rect 9997 -25586 10007 -25526
rect 9607 -25696 10007 -25586
rect 10063 -25526 10463 -25516
rect 10063 -25586 10073 -25526
rect 10133 -25586 10393 -25526
rect 10453 -25586 10463 -25526
rect 10063 -25696 10463 -25586
rect 10521 -25526 10921 -25516
rect 10521 -25586 10531 -25526
rect 10591 -25586 10851 -25526
rect 10911 -25586 10921 -25526
rect 10521 -25696 10921 -25586
rect 10977 -25526 11377 -25516
rect 10977 -25586 10987 -25526
rect 11047 -25586 11307 -25526
rect 11367 -25586 11377 -25526
rect 10977 -25696 11377 -25586
rect 11433 -25526 11833 -25516
rect 11433 -25586 11443 -25526
rect 11503 -25586 11763 -25526
rect 11823 -25586 11833 -25526
rect 11433 -25696 11833 -25586
rect 11891 -25526 12291 -25516
rect 11891 -25586 11901 -25526
rect 11961 -25586 12221 -25526
rect 12281 -25586 12291 -25526
rect 11891 -25696 12291 -25586
rect 12347 -25526 12747 -25516
rect 12347 -25586 12357 -25526
rect 12417 -25586 12677 -25526
rect 12737 -25586 12747 -25526
rect 12347 -25696 12747 -25586
rect 12803 -25526 13203 -25516
rect 12803 -25586 12813 -25526
rect 12873 -25586 13133 -25526
rect 13193 -25586 13203 -25526
rect 12803 -25696 13203 -25586
rect 13261 -25526 13661 -25516
rect 13261 -25586 13271 -25526
rect 13331 -25586 13591 -25526
rect 13651 -25586 13661 -25526
rect 13261 -25696 13661 -25586
rect 13717 -25526 14117 -25516
rect 13717 -25586 13727 -25526
rect 13787 -25586 14047 -25526
rect 14107 -25586 14117 -25526
rect 13717 -25696 14117 -25586
rect 14173 -25526 14573 -25516
rect 14173 -25586 14183 -25526
rect 14243 -25586 14503 -25526
rect 14563 -25586 14573 -25526
rect 14173 -25696 14573 -25586
rect 14631 -25526 15031 -25516
rect 14631 -25586 14641 -25526
rect 14701 -25586 14961 -25526
rect 15021 -25586 15031 -25526
rect 14631 -25696 15031 -25586
rect 15087 -25526 15487 -25516
rect 15087 -25586 15097 -25526
rect 15157 -25586 15417 -25526
rect 15477 -25586 15487 -25526
rect 15087 -25696 15487 -25586
rect 4111 -25766 15487 -25696
rect 4111 -25876 4511 -25766
rect 4111 -25936 4121 -25876
rect 4181 -25936 4441 -25876
rect 4501 -25936 4511 -25876
rect 4111 -25946 4511 -25936
rect 4567 -25876 4967 -25766
rect 4567 -25936 4577 -25876
rect 4637 -25936 4897 -25876
rect 4957 -25936 4967 -25876
rect 4567 -25946 4967 -25936
rect 5023 -25876 5423 -25766
rect 5023 -25936 5033 -25876
rect 5093 -25936 5353 -25876
rect 5413 -25936 5423 -25876
rect 5023 -25946 5423 -25936
rect 5481 -25876 5881 -25766
rect 5481 -25936 5491 -25876
rect 5551 -25936 5811 -25876
rect 5871 -25936 5881 -25876
rect 5481 -25946 5881 -25936
rect 5937 -25876 6337 -25766
rect 5937 -25936 5947 -25876
rect 6007 -25936 6267 -25876
rect 6327 -25936 6337 -25876
rect 5937 -25946 6337 -25936
rect 6393 -25876 6793 -25766
rect 6393 -25936 6403 -25876
rect 6463 -25936 6723 -25876
rect 6783 -25936 6793 -25876
rect 6393 -25946 6793 -25936
rect 6851 -25876 7251 -25766
rect 6851 -25936 6861 -25876
rect 6921 -25936 7181 -25876
rect 7241 -25936 7251 -25876
rect 6851 -25946 7251 -25936
rect 7307 -25876 7707 -25766
rect 7307 -25936 7317 -25876
rect 7377 -25936 7637 -25876
rect 7697 -25936 7707 -25876
rect 7307 -25946 7707 -25936
rect 7763 -25876 8163 -25766
rect 7763 -25936 7773 -25876
rect 7833 -25936 8093 -25876
rect 8153 -25936 8163 -25876
rect 7763 -25946 8163 -25936
rect 8237 -25876 8637 -25766
rect 8237 -25936 8247 -25876
rect 8307 -25936 8567 -25876
rect 8627 -25936 8637 -25876
rect 8237 -25946 8637 -25936
rect 8693 -25876 9093 -25766
rect 8693 -25936 8703 -25876
rect 8763 -25936 9023 -25876
rect 9083 -25936 9093 -25876
rect 8693 -25946 9093 -25936
rect 9151 -25876 9551 -25766
rect 9151 -25936 9161 -25876
rect 9221 -25936 9481 -25876
rect 9541 -25936 9551 -25876
rect 9151 -25946 9551 -25936
rect 9607 -25876 10007 -25766
rect 9607 -25936 9617 -25876
rect 9677 -25936 9937 -25876
rect 9997 -25936 10007 -25876
rect 9607 -25946 10007 -25936
rect 10063 -25876 10463 -25766
rect 10063 -25936 10073 -25876
rect 10133 -25936 10393 -25876
rect 10453 -25936 10463 -25876
rect 10063 -25946 10463 -25936
rect 10521 -25876 10921 -25766
rect 10521 -25936 10531 -25876
rect 10591 -25936 10851 -25876
rect 10911 -25936 10921 -25876
rect 10521 -25946 10921 -25936
rect 10977 -25876 11377 -25766
rect 10977 -25936 10987 -25876
rect 11047 -25936 11307 -25876
rect 11367 -25936 11377 -25876
rect 10977 -25946 11377 -25936
rect 11433 -25876 11833 -25766
rect 11433 -25936 11443 -25876
rect 11503 -25936 11763 -25876
rect 11823 -25936 11833 -25876
rect 11433 -25946 11833 -25936
rect 11891 -25876 12291 -25766
rect 11891 -25936 11901 -25876
rect 11961 -25936 12221 -25876
rect 12281 -25936 12291 -25876
rect 11891 -25946 12291 -25936
rect 12347 -25876 12747 -25766
rect 12347 -25936 12357 -25876
rect 12417 -25936 12677 -25876
rect 12737 -25936 12747 -25876
rect 12347 -25946 12747 -25936
rect 12803 -25876 13203 -25766
rect 12803 -25936 12813 -25876
rect 12873 -25936 13133 -25876
rect 13193 -25936 13203 -25876
rect 12803 -25946 13203 -25936
rect 13261 -25876 13661 -25766
rect 13261 -25936 13271 -25876
rect 13331 -25936 13591 -25876
rect 13651 -25936 13661 -25876
rect 13261 -25946 13661 -25936
rect 13717 -25876 14117 -25766
rect 13717 -25936 13727 -25876
rect 13787 -25936 14047 -25876
rect 14107 -25936 14117 -25876
rect 13717 -25946 14117 -25936
rect 14173 -25876 14573 -25766
rect 14173 -25936 14183 -25876
rect 14243 -25936 14503 -25876
rect 14563 -25936 14573 -25876
rect 14173 -25946 14573 -25936
rect 14631 -25876 15031 -25766
rect 14631 -25936 14641 -25876
rect 14701 -25936 14961 -25876
rect 15021 -25936 15031 -25876
rect 14631 -25946 15031 -25936
rect 15087 -25876 15487 -25766
rect 15087 -25936 15097 -25876
rect 15157 -25936 15417 -25876
rect 15477 -25936 15487 -25876
rect 15087 -25946 15487 -25936
rect 66 -26013 80 -25946
rect 457 -26012 527 -25946
rect 456 -26013 527 -26012
rect 913 -26013 984 -25946
rect 1371 -26013 1442 -25946
rect 1827 -26013 1898 -25946
rect 2283 -26013 2354 -25946
rect 2741 -26013 2812 -25946
rect 3197 -26013 3268 -25946
rect 3653 -26013 3724 -25946
rect 4111 -26013 4182 -25946
rect 4567 -26013 4638 -25946
rect 5023 -26013 5094 -25946
rect 5481 -26013 5552 -25946
rect 5937 -26013 6008 -25946
rect 6393 -26013 6464 -25946
rect 6851 -26013 6922 -25946
rect 7307 -26013 7378 -25946
rect 7763 -26013 7834 -25946
rect 8237 -26013 8308 -25946
rect 8693 -26013 8764 -25946
rect 9151 -26013 9222 -25946
rect 9607 -26013 9678 -25946
rect 10063 -26013 10134 -25946
rect 10521 -26013 10592 -25946
rect 10977 -26013 11048 -25946
rect 11433 -26013 11504 -25946
rect 11891 -26013 11962 -25946
rect 12347 -26013 12418 -25946
rect 12803 -26013 12874 -25946
rect 13261 -26013 13332 -25946
rect 13717 -26013 13788 -25946
rect 14173 -26013 14244 -25946
rect 14631 -26013 14702 -25946
rect 66 -26023 400 -26013
rect 0 -26083 10 -26023
rect 70 -26083 330 -26023
rect 390 -26083 400 -26023
rect 0 -26373 14 -26083
rect 66 -26373 400 -26083
rect 0 -26433 10 -26373
rect 70 -26433 330 -26373
rect 390 -26433 400 -26373
rect 0 -26515 14 -26433
rect 66 -26443 400 -26433
rect 456 -26023 856 -26013
rect 456 -26083 466 -26023
rect 526 -26083 786 -26023
rect 846 -26083 856 -26023
rect 456 -26193 856 -26083
rect 912 -26023 1312 -26013
rect 912 -26083 922 -26023
rect 982 -26083 1242 -26023
rect 1302 -26083 1312 -26023
rect 912 -26193 1312 -26083
rect 1370 -26023 1770 -26013
rect 1370 -26083 1380 -26023
rect 1440 -26083 1700 -26023
rect 1760 -26083 1770 -26023
rect 1370 -26193 1770 -26083
rect 1826 -26023 2226 -26013
rect 1826 -26083 1836 -26023
rect 1896 -26083 2156 -26023
rect 2216 -26083 2226 -26023
rect 1826 -26193 2226 -26083
rect 2282 -26023 2682 -26013
rect 2282 -26083 2292 -26023
rect 2352 -26083 2612 -26023
rect 2672 -26083 2682 -26023
rect 2282 -26193 2682 -26083
rect 2740 -26023 3140 -26013
rect 2740 -26083 2750 -26023
rect 2810 -26083 3070 -26023
rect 3130 -26083 3140 -26023
rect 2740 -26193 3140 -26083
rect 3196 -26023 3596 -26013
rect 3196 -26083 3206 -26023
rect 3266 -26083 3526 -26023
rect 3586 -26083 3596 -26023
rect 3196 -26193 3596 -26083
rect 3652 -26023 4052 -26013
rect 3652 -26083 3662 -26023
rect 3722 -26083 3982 -26023
rect 4042 -26083 4052 -26023
rect 3652 -26193 4052 -26083
rect 456 -26263 4052 -26193
rect 456 -26373 856 -26263
rect 456 -26433 466 -26373
rect 526 -26433 786 -26373
rect 846 -26433 856 -26373
rect 456 -26443 856 -26433
rect 912 -26373 1312 -26263
rect 912 -26433 922 -26373
rect 982 -26433 1242 -26373
rect 1302 -26433 1312 -26373
rect 912 -26443 1312 -26433
rect 1370 -26373 1770 -26263
rect 1370 -26433 1380 -26373
rect 1440 -26433 1700 -26373
rect 1760 -26433 1770 -26373
rect 1370 -26443 1770 -26433
rect 1826 -26373 2226 -26263
rect 1826 -26433 1836 -26373
rect 1896 -26433 2156 -26373
rect 2216 -26433 2226 -26373
rect 1826 -26443 2226 -26433
rect 2282 -26373 2682 -26263
rect 2282 -26433 2292 -26373
rect 2352 -26433 2612 -26373
rect 2672 -26433 2682 -26373
rect 2282 -26443 2682 -26433
rect 2740 -26373 3140 -26263
rect 2740 -26433 2750 -26373
rect 2810 -26433 3070 -26373
rect 3130 -26433 3140 -26373
rect 2740 -26443 3140 -26433
rect 3196 -26373 3596 -26263
rect 3196 -26433 3206 -26373
rect 3266 -26433 3526 -26373
rect 3586 -26433 3596 -26373
rect 3196 -26443 3596 -26433
rect 3652 -26373 4052 -26263
rect 3652 -26433 3662 -26373
rect 3722 -26433 3982 -26373
rect 4042 -26433 4052 -26373
rect 3652 -26443 4052 -26433
rect 4110 -26023 4510 -26013
rect 4110 -26083 4120 -26023
rect 4180 -26083 4440 -26023
rect 4500 -26083 4510 -26023
rect 4110 -26193 4510 -26083
rect 4566 -26023 4966 -26013
rect 4566 -26083 4576 -26023
rect 4636 -26083 4896 -26023
rect 4956 -26083 4966 -26023
rect 4566 -26193 4966 -26083
rect 5022 -26023 5422 -26013
rect 5022 -26083 5032 -26023
rect 5092 -26083 5352 -26023
rect 5412 -26083 5422 -26023
rect 5022 -26193 5422 -26083
rect 5480 -26023 5880 -26013
rect 5480 -26083 5490 -26023
rect 5550 -26083 5810 -26023
rect 5870 -26083 5880 -26023
rect 5480 -26193 5880 -26083
rect 5936 -26023 6336 -26013
rect 5936 -26083 5946 -26023
rect 6006 -26083 6266 -26023
rect 6326 -26083 6336 -26023
rect 5936 -26193 6336 -26083
rect 6392 -26023 6792 -26013
rect 6392 -26083 6402 -26023
rect 6462 -26083 6722 -26023
rect 6782 -26083 6792 -26023
rect 6392 -26193 6792 -26083
rect 6850 -26023 7250 -26013
rect 6850 -26083 6860 -26023
rect 6920 -26083 7180 -26023
rect 7240 -26083 7250 -26023
rect 6850 -26193 7250 -26083
rect 7306 -26023 7706 -26013
rect 7306 -26083 7316 -26023
rect 7376 -26083 7636 -26023
rect 7696 -26083 7706 -26023
rect 7306 -26193 7706 -26083
rect 7762 -26023 8162 -26013
rect 7762 -26083 7772 -26023
rect 7832 -26083 8092 -26023
rect 8152 -26083 8162 -26023
rect 7762 -26193 8162 -26083
rect 8236 -26023 8636 -26013
rect 8236 -26083 8246 -26023
rect 8306 -26083 8566 -26023
rect 8626 -26083 8636 -26023
rect 8236 -26193 8636 -26083
rect 8692 -26023 9092 -26013
rect 8692 -26083 8702 -26023
rect 8762 -26083 9022 -26023
rect 9082 -26083 9092 -26023
rect 8692 -26193 9092 -26083
rect 9150 -26023 9550 -26013
rect 9150 -26083 9160 -26023
rect 9220 -26083 9480 -26023
rect 9540 -26083 9550 -26023
rect 9150 -26193 9550 -26083
rect 9606 -26023 10006 -26013
rect 9606 -26083 9616 -26023
rect 9676 -26083 9936 -26023
rect 9996 -26083 10006 -26023
rect 9606 -26193 10006 -26083
rect 10062 -26023 10462 -26013
rect 10062 -26083 10072 -26023
rect 10132 -26083 10392 -26023
rect 10452 -26083 10462 -26023
rect 10062 -26193 10462 -26083
rect 10520 -26023 10920 -26013
rect 10520 -26083 10530 -26023
rect 10590 -26083 10850 -26023
rect 10910 -26083 10920 -26023
rect 10520 -26193 10920 -26083
rect 10976 -26023 11376 -26013
rect 10976 -26083 10986 -26023
rect 11046 -26083 11306 -26023
rect 11366 -26083 11376 -26023
rect 10976 -26193 11376 -26083
rect 11432 -26023 11832 -26013
rect 11432 -26083 11442 -26023
rect 11502 -26083 11762 -26023
rect 11822 -26083 11832 -26023
rect 11432 -26193 11832 -26083
rect 11890 -26023 12290 -26013
rect 11890 -26083 11900 -26023
rect 11960 -26083 12220 -26023
rect 12280 -26083 12290 -26023
rect 11890 -26193 12290 -26083
rect 12346 -26023 12746 -26013
rect 12346 -26083 12356 -26023
rect 12416 -26083 12676 -26023
rect 12736 -26083 12746 -26023
rect 12346 -26193 12746 -26083
rect 12802 -26023 13202 -26013
rect 12802 -26083 12812 -26023
rect 12872 -26083 13132 -26023
rect 13192 -26083 13202 -26023
rect 12802 -26193 13202 -26083
rect 13260 -26023 13660 -26013
rect 13260 -26083 13270 -26023
rect 13330 -26083 13590 -26023
rect 13650 -26083 13660 -26023
rect 13260 -26193 13660 -26083
rect 13716 -26023 14116 -26013
rect 13716 -26083 13726 -26023
rect 13786 -26083 14046 -26023
rect 14106 -26083 14116 -26023
rect 13716 -26193 14116 -26083
rect 14172 -26023 14572 -26013
rect 14172 -26083 14182 -26023
rect 14242 -26083 14502 -26023
rect 14562 -26083 14572 -26023
rect 14172 -26193 14572 -26083
rect 14630 -26023 15030 -26013
rect 14630 -26083 14640 -26023
rect 14700 -26083 14960 -26023
rect 15020 -26083 15030 -26023
rect 14630 -26193 15030 -26083
rect 15086 -26023 15486 -26013
rect 15086 -26083 15096 -26023
rect 15156 -26083 15416 -26023
rect 15476 -26083 15486 -26023
rect 15086 -26193 15486 -26083
rect 4110 -26263 15486 -26193
rect 4110 -26373 4510 -26263
rect 4110 -26433 4120 -26373
rect 4180 -26433 4440 -26373
rect 4500 -26433 4510 -26373
rect 4110 -26443 4510 -26433
rect 4566 -26373 4966 -26263
rect 4566 -26433 4576 -26373
rect 4636 -26433 4896 -26373
rect 4956 -26433 4966 -26373
rect 4566 -26443 4966 -26433
rect 5022 -26373 5422 -26263
rect 5022 -26433 5032 -26373
rect 5092 -26433 5352 -26373
rect 5412 -26433 5422 -26373
rect 5022 -26443 5422 -26433
rect 5480 -26373 5880 -26263
rect 5480 -26433 5490 -26373
rect 5550 -26433 5810 -26373
rect 5870 -26433 5880 -26373
rect 5480 -26443 5880 -26433
rect 5936 -26373 6336 -26263
rect 5936 -26433 5946 -26373
rect 6006 -26433 6266 -26373
rect 6326 -26433 6336 -26373
rect 5936 -26443 6336 -26433
rect 6392 -26373 6792 -26263
rect 6392 -26433 6402 -26373
rect 6462 -26433 6722 -26373
rect 6782 -26433 6792 -26373
rect 6392 -26443 6792 -26433
rect 6850 -26373 7250 -26263
rect 6850 -26433 6860 -26373
rect 6920 -26433 7180 -26373
rect 7240 -26433 7250 -26373
rect 6850 -26443 7250 -26433
rect 7306 -26373 7706 -26263
rect 7306 -26433 7316 -26373
rect 7376 -26433 7636 -26373
rect 7696 -26433 7706 -26373
rect 7306 -26443 7706 -26433
rect 7762 -26373 8162 -26263
rect 7762 -26433 7772 -26373
rect 7832 -26433 8092 -26373
rect 8152 -26433 8162 -26373
rect 7762 -26443 8162 -26433
rect 8236 -26373 8636 -26263
rect 8236 -26433 8246 -26373
rect 8306 -26433 8566 -26373
rect 8626 -26433 8636 -26373
rect 8236 -26443 8636 -26433
rect 8692 -26373 9092 -26263
rect 8692 -26433 8702 -26373
rect 8762 -26433 9022 -26373
rect 9082 -26433 9092 -26373
rect 8692 -26443 9092 -26433
rect 9150 -26373 9550 -26263
rect 9150 -26433 9160 -26373
rect 9220 -26433 9480 -26373
rect 9540 -26433 9550 -26373
rect 9150 -26443 9550 -26433
rect 9606 -26373 10006 -26263
rect 9606 -26433 9616 -26373
rect 9676 -26433 9936 -26373
rect 9996 -26433 10006 -26373
rect 9606 -26443 10006 -26433
rect 10062 -26373 10462 -26263
rect 10062 -26433 10072 -26373
rect 10132 -26433 10392 -26373
rect 10452 -26433 10462 -26373
rect 10062 -26443 10462 -26433
rect 10520 -26373 10920 -26263
rect 10520 -26433 10530 -26373
rect 10590 -26433 10850 -26373
rect 10910 -26433 10920 -26373
rect 10520 -26443 10920 -26433
rect 10976 -26373 11376 -26263
rect 10976 -26433 10986 -26373
rect 11046 -26433 11306 -26373
rect 11366 -26433 11376 -26373
rect 10976 -26443 11376 -26433
rect 11432 -26373 11832 -26263
rect 11432 -26433 11442 -26373
rect 11502 -26433 11762 -26373
rect 11822 -26433 11832 -26373
rect 11432 -26443 11832 -26433
rect 11890 -26373 12290 -26263
rect 11890 -26433 11900 -26373
rect 11960 -26433 12220 -26373
rect 12280 -26433 12290 -26373
rect 11890 -26443 12290 -26433
rect 12346 -26373 12746 -26263
rect 12346 -26433 12356 -26373
rect 12416 -26433 12676 -26373
rect 12736 -26433 12746 -26373
rect 12346 -26443 12746 -26433
rect 12802 -26373 13202 -26263
rect 12802 -26433 12812 -26373
rect 12872 -26433 13132 -26373
rect 13192 -26433 13202 -26373
rect 12802 -26443 13202 -26433
rect 13260 -26373 13660 -26263
rect 13260 -26433 13270 -26373
rect 13330 -26433 13590 -26373
rect 13650 -26433 13660 -26373
rect 13260 -26443 13660 -26433
rect 13716 -26373 14116 -26263
rect 13716 -26433 13726 -26373
rect 13786 -26433 14046 -26373
rect 14106 -26433 14116 -26373
rect 13716 -26443 14116 -26433
rect 14172 -26373 14572 -26263
rect 14172 -26433 14182 -26373
rect 14242 -26433 14502 -26373
rect 14562 -26433 14572 -26373
rect 14172 -26443 14572 -26433
rect 14630 -26373 15030 -26263
rect 14630 -26433 14640 -26373
rect 14700 -26433 14960 -26373
rect 15020 -26433 15030 -26373
rect 14630 -26443 15030 -26433
rect 15086 -26373 15486 -26263
rect 15086 -26433 15096 -26373
rect 15156 -26433 15416 -26373
rect 15476 -26433 15486 -26373
rect 15086 -26443 15486 -26433
rect 66 -26505 80 -26443
rect 456 -26505 527 -26443
rect 912 -26505 983 -26443
rect 1370 -26505 1441 -26443
rect 1826 -26505 1897 -26443
rect 2282 -26505 2353 -26443
rect 2740 -26505 2810 -26443
rect 3196 -26505 3266 -26443
rect 3652 -26505 3722 -26443
rect 66 -26515 400 -26505
rect 0 -26575 10 -26515
rect 70 -26575 330 -26515
rect 390 -26575 400 -26515
rect 0 -26865 14 -26575
rect 66 -26865 400 -26575
rect 0 -26925 10 -26865
rect 70 -26925 330 -26865
rect 390 -26925 400 -26865
rect 0 -27017 14 -26925
rect 66 -26935 400 -26925
rect 456 -26515 856 -26505
rect 456 -26575 466 -26515
rect 526 -26575 786 -26515
rect 846 -26575 856 -26515
rect 456 -26685 856 -26575
rect 912 -26515 1312 -26505
rect 912 -26575 922 -26515
rect 982 -26575 1242 -26515
rect 1302 -26575 1312 -26515
rect 912 -26685 1312 -26575
rect 1370 -26515 1770 -26505
rect 1370 -26575 1380 -26515
rect 1440 -26575 1700 -26515
rect 1760 -26575 1770 -26515
rect 1370 -26685 1770 -26575
rect 1826 -26515 2226 -26505
rect 1826 -26575 1836 -26515
rect 1896 -26575 2156 -26515
rect 2216 -26575 2226 -26515
rect 1826 -26685 2226 -26575
rect 2282 -26515 2682 -26505
rect 2282 -26575 2292 -26515
rect 2352 -26575 2612 -26515
rect 2672 -26575 2682 -26515
rect 2282 -26685 2682 -26575
rect 456 -26686 2682 -26685
rect 2740 -26515 3140 -26505
rect 2740 -26575 2750 -26515
rect 2810 -26575 3070 -26515
rect 3130 -26575 3140 -26515
rect 2740 -26685 3140 -26575
rect 3196 -26515 3596 -26505
rect 3196 -26575 3206 -26515
rect 3266 -26575 3526 -26515
rect 3586 -26575 3596 -26515
rect 3196 -26685 3596 -26575
rect 3652 -26515 4052 -26505
rect 3652 -26575 3662 -26515
rect 3722 -26575 3982 -26515
rect 4042 -26575 4052 -26515
rect 3652 -26685 4052 -26575
rect 4110 -26515 4510 -26505
rect 4110 -26575 4120 -26515
rect 4180 -26575 4440 -26515
rect 4500 -26575 4510 -26515
rect 4110 -26685 4510 -26575
rect 4566 -26515 4966 -26505
rect 4566 -26575 4576 -26515
rect 4636 -26575 4896 -26515
rect 4956 -26575 4966 -26515
rect 4566 -26685 4966 -26575
rect 5022 -26515 5422 -26505
rect 5022 -26575 5032 -26515
rect 5092 -26575 5352 -26515
rect 5412 -26575 5422 -26515
rect 5022 -26685 5422 -26575
rect 5480 -26515 5880 -26505
rect 5480 -26575 5490 -26515
rect 5550 -26575 5810 -26515
rect 5870 -26575 5880 -26515
rect 5480 -26685 5880 -26575
rect 5936 -26515 6336 -26505
rect 5936 -26575 5946 -26515
rect 6006 -26575 6266 -26515
rect 6326 -26575 6336 -26515
rect 5936 -26685 6336 -26575
rect 6392 -26515 6792 -26505
rect 6392 -26575 6402 -26515
rect 6462 -26575 6722 -26515
rect 6782 -26575 6792 -26515
rect 6392 -26685 6792 -26575
rect 6850 -26515 7250 -26505
rect 6850 -26575 6860 -26515
rect 6920 -26575 7180 -26515
rect 7240 -26575 7250 -26515
rect 6850 -26685 7250 -26575
rect 7306 -26515 7706 -26505
rect 7306 -26575 7316 -26515
rect 7376 -26575 7636 -26515
rect 7696 -26575 7706 -26515
rect 7306 -26685 7706 -26575
rect 7762 -26515 8162 -26505
rect 7762 -26575 7772 -26515
rect 7832 -26575 8092 -26515
rect 8152 -26575 8162 -26515
rect 7762 -26685 8162 -26575
rect 8236 -26515 8636 -26505
rect 8236 -26575 8246 -26515
rect 8306 -26575 8566 -26515
rect 8626 -26575 8636 -26515
rect 8236 -26685 8636 -26575
rect 8692 -26515 9092 -26505
rect 8692 -26575 8702 -26515
rect 8762 -26575 9022 -26515
rect 9082 -26575 9092 -26515
rect 8692 -26685 9092 -26575
rect 9150 -26515 9550 -26505
rect 9150 -26575 9160 -26515
rect 9220 -26575 9480 -26515
rect 9540 -26575 9550 -26515
rect 9150 -26685 9550 -26575
rect 9606 -26515 10006 -26505
rect 9606 -26575 9616 -26515
rect 9676 -26575 9936 -26515
rect 9996 -26575 10006 -26515
rect 9606 -26685 10006 -26575
rect 10062 -26515 10462 -26505
rect 10062 -26575 10072 -26515
rect 10132 -26575 10392 -26515
rect 10452 -26575 10462 -26515
rect 10062 -26685 10462 -26575
rect 2740 -26686 10462 -26685
rect 10520 -26515 10920 -26505
rect 10520 -26575 10530 -26515
rect 10590 -26575 10850 -26515
rect 10910 -26575 10920 -26515
rect 10520 -26685 10920 -26575
rect 10976 -26515 11376 -26505
rect 10976 -26575 10986 -26515
rect 11046 -26575 11306 -26515
rect 11366 -26575 11376 -26515
rect 10976 -26685 11376 -26575
rect 11432 -26515 11832 -26505
rect 11432 -26575 11442 -26515
rect 11502 -26575 11762 -26515
rect 11822 -26575 11832 -26515
rect 11432 -26685 11832 -26575
rect 11890 -26515 12290 -26505
rect 11890 -26575 11900 -26515
rect 11960 -26575 12220 -26515
rect 12280 -26575 12290 -26515
rect 11890 -26685 12290 -26575
rect 12346 -26515 12746 -26505
rect 12346 -26575 12356 -26515
rect 12416 -26575 12676 -26515
rect 12736 -26575 12746 -26515
rect 12346 -26685 12746 -26575
rect 12802 -26515 13202 -26505
rect 12802 -26575 12812 -26515
rect 12872 -26575 13132 -26515
rect 13192 -26575 13202 -26515
rect 12802 -26685 13202 -26575
rect 13260 -26515 13660 -26505
rect 13260 -26575 13270 -26515
rect 13330 -26575 13590 -26515
rect 13650 -26575 13660 -26515
rect 13260 -26685 13660 -26575
rect 13716 -26515 14116 -26505
rect 13716 -26575 13726 -26515
rect 13786 -26575 14046 -26515
rect 14106 -26575 14116 -26515
rect 13716 -26685 14116 -26575
rect 14172 -26515 14572 -26505
rect 14172 -26575 14182 -26515
rect 14242 -26575 14502 -26515
rect 14562 -26575 14572 -26515
rect 14172 -26685 14572 -26575
rect 14630 -26515 15030 -26505
rect 14630 -26575 14640 -26515
rect 14700 -26575 14960 -26515
rect 15020 -26575 15030 -26515
rect 14630 -26685 15030 -26575
rect 15086 -26515 15486 -26505
rect 15086 -26575 15096 -26515
rect 15156 -26575 15416 -26515
rect 15476 -26575 15486 -26515
rect 15086 -26685 15486 -26575
rect 10520 -26686 15486 -26685
rect 456 -26687 15486 -26686
rect 456 -26756 15721 -26687
rect 456 -26865 856 -26756
rect 456 -26925 466 -26865
rect 526 -26925 786 -26865
rect 846 -26925 856 -26865
rect 456 -26935 856 -26925
rect 912 -26865 1312 -26756
rect 912 -26925 922 -26865
rect 982 -26925 1242 -26865
rect 1302 -26925 1312 -26865
rect 912 -26935 1312 -26925
rect 1370 -26865 1770 -26756
rect 1370 -26925 1380 -26865
rect 1440 -26925 1700 -26865
rect 1760 -26925 1770 -26865
rect 1370 -26935 1770 -26925
rect 1826 -26865 2226 -26756
rect 1826 -26925 1836 -26865
rect 1896 -26925 2156 -26865
rect 2216 -26925 2226 -26865
rect 1826 -26935 2226 -26925
rect 2282 -26865 2682 -26756
rect 2282 -26925 2292 -26865
rect 2352 -26925 2612 -26865
rect 2672 -26925 2682 -26865
rect 2282 -26935 2682 -26925
rect 2740 -26865 3140 -26756
rect 2740 -26925 2750 -26865
rect 2810 -26925 3070 -26865
rect 3130 -26925 3140 -26865
rect 2740 -26935 3140 -26925
rect 3196 -26865 3596 -26756
rect 3196 -26925 3206 -26865
rect 3266 -26925 3526 -26865
rect 3586 -26925 3596 -26865
rect 3196 -26935 3596 -26925
rect 3652 -26865 4052 -26756
rect 3652 -26925 3662 -26865
rect 3722 -26925 3982 -26865
rect 4042 -26925 4052 -26865
rect 3652 -26935 4052 -26925
rect 4110 -26865 4510 -26756
rect 4110 -26925 4120 -26865
rect 4180 -26925 4440 -26865
rect 4500 -26925 4510 -26865
rect 4110 -26935 4510 -26925
rect 4566 -26865 4966 -26756
rect 4566 -26925 4576 -26865
rect 4636 -26925 4896 -26865
rect 4956 -26925 4966 -26865
rect 4566 -26935 4966 -26925
rect 5022 -26865 5422 -26756
rect 5022 -26925 5032 -26865
rect 5092 -26925 5352 -26865
rect 5412 -26925 5422 -26865
rect 5022 -26935 5422 -26925
rect 5480 -26865 5880 -26756
rect 5480 -26925 5490 -26865
rect 5550 -26925 5810 -26865
rect 5870 -26925 5880 -26865
rect 5480 -26935 5880 -26925
rect 5936 -26865 6336 -26756
rect 5936 -26925 5946 -26865
rect 6006 -26925 6266 -26865
rect 6326 -26925 6336 -26865
rect 5936 -26935 6336 -26925
rect 6392 -26865 6792 -26756
rect 6392 -26925 6402 -26865
rect 6462 -26925 6722 -26865
rect 6782 -26925 6792 -26865
rect 6392 -26935 6792 -26925
rect 6850 -26865 7250 -26756
rect 6850 -26925 6860 -26865
rect 6920 -26925 7180 -26865
rect 7240 -26925 7250 -26865
rect 6850 -26935 7250 -26925
rect 7306 -26865 7706 -26756
rect 7306 -26925 7316 -26865
rect 7376 -26925 7636 -26865
rect 7696 -26925 7706 -26865
rect 7306 -26935 7706 -26925
rect 7762 -26865 8162 -26756
rect 7762 -26925 7772 -26865
rect 7832 -26925 8092 -26865
rect 8152 -26925 8162 -26865
rect 7762 -26935 8162 -26925
rect 8236 -26865 8636 -26756
rect 8236 -26925 8246 -26865
rect 8306 -26925 8566 -26865
rect 8626 -26925 8636 -26865
rect 8236 -26935 8636 -26925
rect 8692 -26865 9092 -26756
rect 8692 -26925 8702 -26865
rect 8762 -26925 9022 -26865
rect 9082 -26925 9092 -26865
rect 8692 -26935 9092 -26925
rect 9150 -26865 9550 -26756
rect 9150 -26925 9160 -26865
rect 9220 -26925 9480 -26865
rect 9540 -26925 9550 -26865
rect 9150 -26935 9550 -26925
rect 9606 -26865 10006 -26756
rect 9606 -26925 9616 -26865
rect 9676 -26925 9936 -26865
rect 9996 -26925 10006 -26865
rect 9606 -26935 10006 -26925
rect 10062 -26865 10462 -26756
rect 10062 -26925 10072 -26865
rect 10132 -26925 10392 -26865
rect 10452 -26925 10462 -26865
rect 10062 -26935 10462 -26925
rect 10520 -26865 10920 -26756
rect 10520 -26925 10530 -26865
rect 10590 -26925 10850 -26865
rect 10910 -26925 10920 -26865
rect 10520 -26935 10920 -26925
rect 10976 -26865 11376 -26756
rect 10976 -26925 10986 -26865
rect 11046 -26925 11306 -26865
rect 11366 -26925 11376 -26865
rect 10976 -26935 11376 -26925
rect 11432 -26865 11832 -26756
rect 11432 -26925 11442 -26865
rect 11502 -26925 11762 -26865
rect 11822 -26925 11832 -26865
rect 11432 -26935 11832 -26925
rect 11890 -26865 12290 -26756
rect 11890 -26925 11900 -26865
rect 11960 -26925 12220 -26865
rect 12280 -26925 12290 -26865
rect 11890 -26935 12290 -26925
rect 12346 -26865 12746 -26756
rect 12346 -26925 12356 -26865
rect 12416 -26925 12676 -26865
rect 12736 -26925 12746 -26865
rect 12346 -26935 12746 -26925
rect 12802 -26865 13202 -26756
rect 12802 -26925 12812 -26865
rect 12872 -26925 13132 -26865
rect 13192 -26925 13202 -26865
rect 12802 -26935 13202 -26925
rect 13260 -26865 13660 -26756
rect 13260 -26925 13270 -26865
rect 13330 -26925 13590 -26865
rect 13650 -26925 13660 -26865
rect 13260 -26935 13660 -26925
rect 13716 -26865 14116 -26756
rect 13716 -26925 13726 -26865
rect 13786 -26925 14046 -26865
rect 14106 -26925 14116 -26865
rect 13716 -26935 14116 -26925
rect 14172 -26865 14572 -26756
rect 14172 -26925 14182 -26865
rect 14242 -26925 14502 -26865
rect 14562 -26925 14572 -26865
rect 14172 -26935 14572 -26925
rect 14630 -26865 15030 -26756
rect 14630 -26925 14640 -26865
rect 14700 -26925 14960 -26865
rect 15020 -26925 15030 -26865
rect 14630 -26935 15030 -26925
rect 15086 -26758 15721 -26756
rect 15086 -26865 15486 -26758
rect 15086 -26925 15096 -26865
rect 15156 -26925 15416 -26865
rect 15476 -26925 15486 -26865
rect 15086 -26935 15486 -26925
rect 66 -27007 80 -26935
rect 456 -27007 526 -26935
rect 912 -27007 983 -26935
rect 1370 -27007 1441 -26935
rect 1826 -27007 1897 -26935
rect 2282 -27007 2353 -26935
rect 2740 -27007 2811 -26935
rect 3196 -27007 3267 -26935
rect 3652 -27007 3723 -26935
rect 4110 -27007 4181 -26935
rect 4566 -27007 4637 -26935
rect 5022 -27007 5093 -26935
rect 5480 -27007 5551 -26935
rect 5936 -27007 6007 -26935
rect 6392 -27007 6463 -26935
rect 6850 -27007 6921 -26935
rect 7306 -27007 7377 -26935
rect 7762 -27007 7833 -26935
rect 8236 -27007 8307 -26935
rect 8692 -27007 8763 -26935
rect 9150 -27007 9221 -26935
rect 9606 -27007 9677 -26935
rect 10062 -27007 10133 -26935
rect 10520 -27007 10591 -26935
rect 10976 -27007 11047 -26935
rect 11432 -27007 11503 -26935
rect 11890 -27007 11961 -26935
rect 12346 -27007 12417 -26935
rect 12802 -27007 12873 -26935
rect 13260 -27007 13331 -26935
rect 13716 -27007 13787 -26935
rect 14172 -27007 14243 -26935
rect 14630 -27007 14701 -26935
rect 66 -27017 400 -27007
rect 0 -27077 10 -27017
rect 70 -27077 330 -27017
rect 390 -27077 400 -27017
rect 0 -27367 14 -27077
rect 66 -27367 400 -27077
rect 0 -27427 10 -27367
rect 70 -27427 330 -27367
rect 390 -27427 400 -27367
rect 0 -27533 14 -27427
rect 66 -27437 400 -27427
rect 456 -27017 856 -27007
rect 456 -27077 466 -27017
rect 526 -27077 786 -27017
rect 846 -27077 856 -27017
rect 456 -27187 856 -27077
rect 912 -27017 1312 -27007
rect 912 -27077 922 -27017
rect 982 -27077 1242 -27017
rect 1302 -27077 1312 -27017
rect 912 -27187 1312 -27077
rect 1370 -27017 1770 -27007
rect 1370 -27077 1380 -27017
rect 1440 -27077 1700 -27017
rect 1760 -27077 1770 -27017
rect 1370 -27187 1770 -27077
rect 1826 -27017 2226 -27007
rect 1826 -27077 1836 -27017
rect 1896 -27077 2156 -27017
rect 2216 -27077 2226 -27017
rect 1826 -27187 2226 -27077
rect 2282 -27017 2682 -27007
rect 2282 -27077 2292 -27017
rect 2352 -27077 2612 -27017
rect 2672 -27077 2682 -27017
rect 2282 -27187 2682 -27077
rect 2740 -27017 3140 -27007
rect 2740 -27077 2750 -27017
rect 2810 -27077 3070 -27017
rect 3130 -27077 3140 -27017
rect 2740 -27187 3140 -27077
rect 3196 -27017 3596 -27007
rect 3196 -27077 3206 -27017
rect 3266 -27077 3526 -27017
rect 3586 -27077 3596 -27017
rect 3196 -27187 3596 -27077
rect 3652 -27017 4052 -27007
rect 3652 -27077 3662 -27017
rect 3722 -27077 3982 -27017
rect 4042 -27077 4052 -27017
rect 3652 -27187 4052 -27077
rect 4110 -27017 4510 -27007
rect 4110 -27077 4120 -27017
rect 4180 -27077 4440 -27017
rect 4500 -27077 4510 -27017
rect 4110 -27187 4510 -27077
rect 4566 -27017 4966 -27007
rect 4566 -27077 4576 -27017
rect 4636 -27077 4896 -27017
rect 4956 -27077 4966 -27017
rect 4566 -27187 4966 -27077
rect 5022 -27017 5422 -27007
rect 5022 -27077 5032 -27017
rect 5092 -27077 5352 -27017
rect 5412 -27077 5422 -27017
rect 5022 -27187 5422 -27077
rect 5480 -27017 5880 -27007
rect 5480 -27077 5490 -27017
rect 5550 -27077 5810 -27017
rect 5870 -27077 5880 -27017
rect 5480 -27187 5880 -27077
rect 5936 -27017 6336 -27007
rect 5936 -27077 5946 -27017
rect 6006 -27077 6266 -27017
rect 6326 -27077 6336 -27017
rect 5936 -27187 6336 -27077
rect 6392 -27017 6792 -27007
rect 6392 -27077 6402 -27017
rect 6462 -27077 6722 -27017
rect 6782 -27077 6792 -27017
rect 6392 -27187 6792 -27077
rect 6850 -27017 7250 -27007
rect 6850 -27077 6860 -27017
rect 6920 -27077 7180 -27017
rect 7240 -27077 7250 -27017
rect 6850 -27187 7250 -27077
rect 7306 -27017 7706 -27007
rect 7306 -27077 7316 -27017
rect 7376 -27077 7636 -27017
rect 7696 -27077 7706 -27017
rect 7306 -27187 7706 -27077
rect 7762 -27017 8162 -27007
rect 7762 -27077 7772 -27017
rect 7832 -27077 8092 -27017
rect 8152 -27077 8162 -27017
rect 7762 -27187 8162 -27077
rect 8236 -27017 8636 -27007
rect 8236 -27077 8246 -27017
rect 8306 -27077 8566 -27017
rect 8626 -27077 8636 -27017
rect 8236 -27187 8636 -27077
rect 8692 -27017 9092 -27007
rect 8692 -27077 8702 -27017
rect 8762 -27077 9022 -27017
rect 9082 -27077 9092 -27017
rect 8692 -27187 9092 -27077
rect 9150 -27017 9550 -27007
rect 9150 -27077 9160 -27017
rect 9220 -27077 9480 -27017
rect 9540 -27077 9550 -27017
rect 9150 -27187 9550 -27077
rect 9606 -27017 10006 -27007
rect 9606 -27077 9616 -27017
rect 9676 -27077 9936 -27017
rect 9996 -27077 10006 -27017
rect 9606 -27187 10006 -27077
rect 10062 -27017 10462 -27007
rect 10062 -27077 10072 -27017
rect 10132 -27077 10392 -27017
rect 10452 -27077 10462 -27017
rect 10062 -27187 10462 -27077
rect 10520 -27017 10920 -27007
rect 10520 -27077 10530 -27017
rect 10590 -27077 10850 -27017
rect 10910 -27077 10920 -27017
rect 10520 -27187 10920 -27077
rect 10976 -27017 11376 -27007
rect 10976 -27077 10986 -27017
rect 11046 -27077 11306 -27017
rect 11366 -27077 11376 -27017
rect 10976 -27187 11376 -27077
rect 11432 -27017 11832 -27007
rect 11432 -27077 11442 -27017
rect 11502 -27077 11762 -27017
rect 11822 -27077 11832 -27017
rect 11432 -27187 11832 -27077
rect 11890 -27017 12290 -27007
rect 11890 -27077 11900 -27017
rect 11960 -27077 12220 -27017
rect 12280 -27077 12290 -27017
rect 11890 -27187 12290 -27077
rect 12346 -27017 12746 -27007
rect 12346 -27077 12356 -27017
rect 12416 -27077 12676 -27017
rect 12736 -27077 12746 -27017
rect 12346 -27187 12746 -27077
rect 12802 -27017 13202 -27007
rect 12802 -27077 12812 -27017
rect 12872 -27077 13132 -27017
rect 13192 -27077 13202 -27017
rect 12802 -27187 13202 -27077
rect 13260 -27017 13660 -27007
rect 13260 -27077 13270 -27017
rect 13330 -27077 13590 -27017
rect 13650 -27077 13660 -27017
rect 13260 -27187 13660 -27077
rect 13716 -27017 14116 -27007
rect 13716 -27077 13726 -27017
rect 13786 -27077 14046 -27017
rect 14106 -27077 14116 -27017
rect 13716 -27187 14116 -27077
rect 14172 -27017 14572 -27007
rect 14172 -27077 14182 -27017
rect 14242 -27077 14502 -27017
rect 14562 -27077 14572 -27017
rect 14172 -27187 14572 -27077
rect 14630 -27017 15030 -27007
rect 14630 -27077 14640 -27017
rect 14700 -27077 14960 -27017
rect 15020 -27077 15030 -27017
rect 14630 -27187 15030 -27077
rect 15086 -27017 15486 -27007
rect 15086 -27077 15096 -27017
rect 15156 -27077 15416 -27017
rect 15476 -27077 15486 -27017
rect 15086 -27187 15486 -27077
rect 456 -27257 15486 -27187
rect 456 -27367 856 -27257
rect 456 -27427 466 -27367
rect 526 -27427 786 -27367
rect 846 -27427 856 -27367
rect 456 -27437 856 -27427
rect 912 -27367 1312 -27257
rect 912 -27427 922 -27367
rect 982 -27427 1242 -27367
rect 1302 -27427 1312 -27367
rect 912 -27437 1312 -27427
rect 1370 -27367 1770 -27257
rect 1370 -27427 1380 -27367
rect 1440 -27427 1700 -27367
rect 1760 -27427 1770 -27367
rect 1370 -27437 1770 -27427
rect 1826 -27367 2226 -27257
rect 1826 -27427 1836 -27367
rect 1896 -27427 2156 -27367
rect 2216 -27427 2226 -27367
rect 1826 -27437 2226 -27427
rect 2282 -27367 2682 -27257
rect 2282 -27427 2292 -27367
rect 2352 -27427 2612 -27367
rect 2672 -27427 2682 -27367
rect 2282 -27437 2682 -27427
rect 2740 -27367 3140 -27257
rect 2740 -27427 2750 -27367
rect 2810 -27427 3070 -27367
rect 3130 -27427 3140 -27367
rect 2740 -27437 3140 -27427
rect 3196 -27367 3596 -27257
rect 3196 -27427 3206 -27367
rect 3266 -27427 3526 -27367
rect 3586 -27427 3596 -27367
rect 3196 -27437 3596 -27427
rect 3652 -27367 4052 -27257
rect 3652 -27427 3662 -27367
rect 3722 -27427 3982 -27367
rect 4042 -27427 4052 -27367
rect 3652 -27437 4052 -27427
rect 4110 -27367 4510 -27257
rect 4110 -27427 4120 -27367
rect 4180 -27427 4440 -27367
rect 4500 -27427 4510 -27367
rect 4110 -27437 4510 -27427
rect 4566 -27367 4966 -27257
rect 4566 -27427 4576 -27367
rect 4636 -27427 4896 -27367
rect 4956 -27427 4966 -27367
rect 4566 -27437 4966 -27427
rect 5022 -27367 5422 -27257
rect 5022 -27427 5032 -27367
rect 5092 -27427 5352 -27367
rect 5412 -27427 5422 -27367
rect 5022 -27437 5422 -27427
rect 5480 -27367 5880 -27257
rect 5480 -27427 5490 -27367
rect 5550 -27427 5810 -27367
rect 5870 -27427 5880 -27367
rect 5480 -27437 5880 -27427
rect 5936 -27367 6336 -27257
rect 5936 -27427 5946 -27367
rect 6006 -27427 6266 -27367
rect 6326 -27427 6336 -27367
rect 5936 -27437 6336 -27427
rect 6392 -27367 6792 -27257
rect 6392 -27427 6402 -27367
rect 6462 -27427 6722 -27367
rect 6782 -27427 6792 -27367
rect 6392 -27437 6792 -27427
rect 6850 -27367 7250 -27257
rect 6850 -27427 6860 -27367
rect 6920 -27427 7180 -27367
rect 7240 -27427 7250 -27367
rect 6850 -27437 7250 -27427
rect 7306 -27367 7706 -27257
rect 7306 -27427 7316 -27367
rect 7376 -27427 7636 -27367
rect 7696 -27427 7706 -27367
rect 7306 -27437 7706 -27427
rect 7762 -27367 8162 -27257
rect 7762 -27427 7772 -27367
rect 7832 -27427 8092 -27367
rect 8152 -27427 8162 -27367
rect 7762 -27437 8162 -27427
rect 8236 -27367 8636 -27257
rect 8236 -27427 8246 -27367
rect 8306 -27427 8566 -27367
rect 8626 -27427 8636 -27367
rect 8236 -27437 8636 -27427
rect 8692 -27367 9092 -27257
rect 8692 -27427 8702 -27367
rect 8762 -27427 9022 -27367
rect 9082 -27427 9092 -27367
rect 8692 -27437 9092 -27427
rect 9150 -27367 9550 -27257
rect 9150 -27427 9160 -27367
rect 9220 -27427 9480 -27367
rect 9540 -27427 9550 -27367
rect 9150 -27437 9550 -27427
rect 9606 -27367 10006 -27257
rect 9606 -27427 9616 -27367
rect 9676 -27427 9936 -27367
rect 9996 -27427 10006 -27367
rect 9606 -27437 10006 -27427
rect 10062 -27367 10462 -27257
rect 10062 -27427 10072 -27367
rect 10132 -27427 10392 -27367
rect 10452 -27427 10462 -27367
rect 10062 -27437 10462 -27427
rect 10520 -27367 10920 -27257
rect 10520 -27427 10530 -27367
rect 10590 -27427 10850 -27367
rect 10910 -27427 10920 -27367
rect 10520 -27437 10920 -27427
rect 10976 -27367 11376 -27257
rect 10976 -27427 10986 -27367
rect 11046 -27427 11306 -27367
rect 11366 -27427 11376 -27367
rect 10976 -27437 11376 -27427
rect 11432 -27367 11832 -27257
rect 11432 -27427 11442 -27367
rect 11502 -27427 11762 -27367
rect 11822 -27427 11832 -27367
rect 11432 -27437 11832 -27427
rect 11890 -27367 12290 -27257
rect 11890 -27427 11900 -27367
rect 11960 -27427 12220 -27367
rect 12280 -27427 12290 -27367
rect 11890 -27437 12290 -27427
rect 12346 -27367 12746 -27257
rect 12346 -27427 12356 -27367
rect 12416 -27427 12676 -27367
rect 12736 -27427 12746 -27367
rect 12346 -27437 12746 -27427
rect 12802 -27367 13202 -27257
rect 12802 -27427 12812 -27367
rect 12872 -27427 13132 -27367
rect 13192 -27427 13202 -27367
rect 12802 -27437 13202 -27427
rect 13260 -27367 13660 -27257
rect 13260 -27427 13270 -27367
rect 13330 -27427 13590 -27367
rect 13650 -27427 13660 -27367
rect 13260 -27437 13660 -27427
rect 13716 -27367 14116 -27257
rect 13716 -27427 13726 -27367
rect 13786 -27427 14046 -27367
rect 14106 -27427 14116 -27367
rect 13716 -27437 14116 -27427
rect 14172 -27367 14572 -27257
rect 14172 -27427 14182 -27367
rect 14242 -27427 14502 -27367
rect 14562 -27427 14572 -27367
rect 14172 -27437 14572 -27427
rect 14630 -27367 15030 -27257
rect 14630 -27427 14640 -27367
rect 14700 -27427 14960 -27367
rect 15020 -27427 15030 -27367
rect 14630 -27437 15030 -27427
rect 15086 -27367 15486 -27257
rect 15086 -27427 15096 -27367
rect 15156 -27427 15416 -27367
rect 15476 -27427 15486 -27367
rect 15086 -27437 15486 -27427
rect 66 -27523 80 -27437
rect 456 -27523 526 -27437
rect 912 -27523 982 -27437
rect 1370 -27523 1440 -27437
rect 1826 -27523 1896 -27437
rect 2282 -27523 2352 -27437
rect 2740 -27523 2810 -27437
rect 3196 -27523 3266 -27437
rect 3652 -27523 3722 -27437
rect 4110 -27523 4180 -27437
rect 4566 -27523 4636 -27437
rect 5022 -27523 5092 -27437
rect 5480 -27523 5550 -27437
rect 5936 -27523 6006 -27437
rect 6392 -27523 6462 -27437
rect 6850 -27523 6920 -27437
rect 7306 -27523 7376 -27437
rect 7762 -27523 7832 -27437
rect 8236 -27523 8306 -27437
rect 8692 -27523 8762 -27437
rect 9150 -27523 9220 -27437
rect 9606 -27523 9676 -27437
rect 10062 -27523 10132 -27437
rect 10520 -27523 10590 -27437
rect 10976 -27523 11046 -27437
rect 11432 -27523 11502 -27437
rect 11890 -27523 11960 -27437
rect 12346 -27523 12416 -27437
rect 12802 -27523 12872 -27437
rect 13260 -27523 13330 -27437
rect 13716 -27523 13786 -27437
rect 14172 -27523 14242 -27437
rect 14630 -27523 14700 -27437
rect 66 -27533 400 -27523
rect 0 -27593 10 -27533
rect 70 -27593 330 -27533
rect 390 -27593 400 -27533
rect 0 -27883 14 -27593
rect 66 -27883 400 -27593
rect 0 -27943 10 -27883
rect 70 -27943 330 -27883
rect 390 -27943 400 -27883
rect 0 -28025 14 -27943
rect 66 -27953 400 -27943
rect 456 -27533 856 -27523
rect 456 -27593 466 -27533
rect 526 -27593 786 -27533
rect 846 -27593 856 -27533
rect 456 -27701 856 -27593
rect 912 -27533 1312 -27523
rect 912 -27593 922 -27533
rect 982 -27593 1242 -27533
rect 1302 -27593 1312 -27533
rect 912 -27701 1312 -27593
rect 1370 -27533 1770 -27523
rect 1370 -27593 1380 -27533
rect 1440 -27593 1700 -27533
rect 1760 -27593 1770 -27533
rect 1370 -27701 1770 -27593
rect 1826 -27533 2226 -27523
rect 1826 -27593 1836 -27533
rect 1896 -27593 2156 -27533
rect 2216 -27593 2226 -27533
rect 1826 -27701 2226 -27593
rect 2282 -27533 2682 -27523
rect 2282 -27593 2292 -27533
rect 2352 -27593 2612 -27533
rect 2672 -27593 2682 -27533
rect 2282 -27701 2682 -27593
rect 2740 -27533 3140 -27523
rect 2740 -27593 2750 -27533
rect 2810 -27593 3070 -27533
rect 3130 -27593 3140 -27533
rect 2740 -27701 3140 -27593
rect 3196 -27533 3596 -27523
rect 3196 -27593 3206 -27533
rect 3266 -27593 3526 -27533
rect 3586 -27593 3596 -27533
rect 3196 -27701 3596 -27593
rect 3652 -27533 4052 -27523
rect 3652 -27593 3662 -27533
rect 3722 -27593 3982 -27533
rect 4042 -27593 4052 -27533
rect 3652 -27701 4052 -27593
rect 4110 -27533 4510 -27523
rect 4110 -27593 4120 -27533
rect 4180 -27593 4440 -27533
rect 4500 -27593 4510 -27533
rect 4110 -27701 4510 -27593
rect 4566 -27533 4966 -27523
rect 4566 -27593 4576 -27533
rect 4636 -27593 4896 -27533
rect 4956 -27593 4966 -27533
rect 4566 -27701 4966 -27593
rect 5022 -27533 5422 -27523
rect 5022 -27593 5032 -27533
rect 5092 -27593 5352 -27533
rect 5412 -27593 5422 -27533
rect 5022 -27701 5422 -27593
rect 5480 -27533 5880 -27523
rect 5480 -27593 5490 -27533
rect 5550 -27593 5810 -27533
rect 5870 -27593 5880 -27533
rect 5480 -27701 5880 -27593
rect 5936 -27533 6336 -27523
rect 5936 -27593 5946 -27533
rect 6006 -27593 6266 -27533
rect 6326 -27593 6336 -27533
rect 5936 -27701 6336 -27593
rect 6392 -27533 6792 -27523
rect 6392 -27593 6402 -27533
rect 6462 -27593 6722 -27533
rect 6782 -27593 6792 -27533
rect 6392 -27701 6792 -27593
rect 6850 -27533 7250 -27523
rect 6850 -27593 6860 -27533
rect 6920 -27593 7180 -27533
rect 7240 -27593 7250 -27533
rect 6850 -27701 7250 -27593
rect 7306 -27533 7706 -27523
rect 7306 -27593 7316 -27533
rect 7376 -27593 7636 -27533
rect 7696 -27593 7706 -27533
rect 7306 -27701 7706 -27593
rect 7762 -27533 8162 -27523
rect 7762 -27593 7772 -27533
rect 7832 -27593 8092 -27533
rect 8152 -27593 8162 -27533
rect 7762 -27701 8162 -27593
rect 8236 -27533 8636 -27523
rect 8236 -27593 8246 -27533
rect 8306 -27593 8566 -27533
rect 8626 -27593 8636 -27533
rect 8236 -27701 8636 -27593
rect 8692 -27533 9092 -27523
rect 8692 -27593 8702 -27533
rect 8762 -27593 9022 -27533
rect 9082 -27593 9092 -27533
rect 8692 -27701 9092 -27593
rect 9150 -27533 9550 -27523
rect 9150 -27593 9160 -27533
rect 9220 -27593 9480 -27533
rect 9540 -27593 9550 -27533
rect 9150 -27701 9550 -27593
rect 9606 -27533 10006 -27523
rect 9606 -27593 9616 -27533
rect 9676 -27593 9936 -27533
rect 9996 -27593 10006 -27533
rect 9606 -27701 10006 -27593
rect 10062 -27533 10462 -27523
rect 10062 -27593 10072 -27533
rect 10132 -27593 10392 -27533
rect 10452 -27593 10462 -27533
rect 10062 -27701 10462 -27593
rect 10520 -27533 10920 -27523
rect 10520 -27593 10530 -27533
rect 10590 -27593 10850 -27533
rect 10910 -27593 10920 -27533
rect 10520 -27701 10920 -27593
rect 10976 -27533 11376 -27523
rect 10976 -27593 10986 -27533
rect 11046 -27593 11306 -27533
rect 11366 -27593 11376 -27533
rect 10976 -27701 11376 -27593
rect 11432 -27533 11832 -27523
rect 11432 -27593 11442 -27533
rect 11502 -27593 11762 -27533
rect 11822 -27593 11832 -27533
rect 11432 -27701 11832 -27593
rect 11890 -27533 12290 -27523
rect 11890 -27593 11900 -27533
rect 11960 -27593 12220 -27533
rect 12280 -27593 12290 -27533
rect 11890 -27701 12290 -27593
rect 12346 -27533 12746 -27523
rect 12346 -27593 12356 -27533
rect 12416 -27593 12676 -27533
rect 12736 -27593 12746 -27533
rect 12346 -27701 12746 -27593
rect 12802 -27533 13202 -27523
rect 12802 -27593 12812 -27533
rect 12872 -27593 13132 -27533
rect 13192 -27593 13202 -27533
rect 12802 -27701 13202 -27593
rect 13260 -27533 13660 -27523
rect 13260 -27593 13270 -27533
rect 13330 -27593 13590 -27533
rect 13650 -27593 13660 -27533
rect 13260 -27701 13660 -27593
rect 13716 -27533 14116 -27523
rect 13716 -27593 13726 -27533
rect 13786 -27593 14046 -27533
rect 14106 -27593 14116 -27533
rect 13716 -27701 14116 -27593
rect 14172 -27533 14572 -27523
rect 14172 -27593 14182 -27533
rect 14242 -27593 14502 -27533
rect 14562 -27593 14572 -27533
rect 14172 -27701 14572 -27593
rect 14630 -27533 15030 -27523
rect 14630 -27593 14640 -27533
rect 14700 -27593 14960 -27533
rect 15020 -27593 15030 -27533
rect 14630 -27701 15030 -27593
rect 15086 -27533 15486 -27523
rect 15086 -27593 15096 -27533
rect 15156 -27593 15416 -27533
rect 15476 -27593 15486 -27533
rect 15086 -27701 15486 -27593
rect 456 -27771 15486 -27701
rect 456 -27773 2682 -27771
rect 456 -27883 856 -27773
rect 456 -27943 466 -27883
rect 526 -27943 786 -27883
rect 846 -27943 856 -27883
rect 456 -27953 856 -27943
rect 912 -27883 1312 -27773
rect 912 -27943 922 -27883
rect 982 -27943 1242 -27883
rect 1302 -27943 1312 -27883
rect 912 -27953 1312 -27943
rect 1370 -27883 1770 -27773
rect 1370 -27943 1380 -27883
rect 1440 -27943 1700 -27883
rect 1760 -27943 1770 -27883
rect 1370 -27953 1770 -27943
rect 1826 -27883 2226 -27773
rect 1826 -27943 1836 -27883
rect 1896 -27943 2156 -27883
rect 2216 -27943 2226 -27883
rect 1826 -27953 2226 -27943
rect 2282 -27883 2682 -27773
rect 2282 -27943 2292 -27883
rect 2352 -27943 2612 -27883
rect 2672 -27943 2682 -27883
rect 2282 -27953 2682 -27943
rect 2740 -27773 10462 -27771
rect 2740 -27883 3140 -27773
rect 2740 -27943 2750 -27883
rect 2810 -27943 3070 -27883
rect 3130 -27943 3140 -27883
rect 2740 -27953 3140 -27943
rect 3196 -27883 3596 -27773
rect 3196 -27943 3206 -27883
rect 3266 -27943 3526 -27883
rect 3586 -27943 3596 -27883
rect 3196 -27953 3596 -27943
rect 3652 -27883 4052 -27773
rect 3652 -27943 3662 -27883
rect 3722 -27943 3982 -27883
rect 4042 -27943 4052 -27883
rect 3652 -27953 4052 -27943
rect 4110 -27883 4510 -27773
rect 4110 -27943 4120 -27883
rect 4180 -27943 4440 -27883
rect 4500 -27943 4510 -27883
rect 4110 -27953 4510 -27943
rect 4566 -27883 4966 -27773
rect 4566 -27943 4576 -27883
rect 4636 -27943 4896 -27883
rect 4956 -27943 4966 -27883
rect 4566 -27953 4966 -27943
rect 5022 -27883 5422 -27773
rect 5022 -27943 5032 -27883
rect 5092 -27943 5352 -27883
rect 5412 -27943 5422 -27883
rect 5022 -27953 5422 -27943
rect 5480 -27883 5880 -27773
rect 5480 -27943 5490 -27883
rect 5550 -27943 5810 -27883
rect 5870 -27943 5880 -27883
rect 5480 -27953 5880 -27943
rect 5936 -27883 6336 -27773
rect 5936 -27943 5946 -27883
rect 6006 -27943 6266 -27883
rect 6326 -27943 6336 -27883
rect 5936 -27953 6336 -27943
rect 6392 -27883 6792 -27773
rect 6392 -27943 6402 -27883
rect 6462 -27943 6722 -27883
rect 6782 -27943 6792 -27883
rect 6392 -27953 6792 -27943
rect 6850 -27883 7250 -27773
rect 6850 -27943 6860 -27883
rect 6920 -27943 7180 -27883
rect 7240 -27943 7250 -27883
rect 6850 -27953 7250 -27943
rect 7306 -27883 7706 -27773
rect 7306 -27943 7316 -27883
rect 7376 -27943 7636 -27883
rect 7696 -27943 7706 -27883
rect 7306 -27953 7706 -27943
rect 7762 -27883 8162 -27773
rect 7762 -27943 7772 -27883
rect 7832 -27943 8092 -27883
rect 8152 -27943 8162 -27883
rect 7762 -27953 8162 -27943
rect 8236 -27883 8636 -27773
rect 8236 -27943 8246 -27883
rect 8306 -27943 8566 -27883
rect 8626 -27943 8636 -27883
rect 8236 -27953 8636 -27943
rect 8692 -27883 9092 -27773
rect 8692 -27943 8702 -27883
rect 8762 -27943 9022 -27883
rect 9082 -27943 9092 -27883
rect 8692 -27953 9092 -27943
rect 9150 -27883 9550 -27773
rect 9150 -27943 9160 -27883
rect 9220 -27943 9480 -27883
rect 9540 -27943 9550 -27883
rect 9150 -27953 9550 -27943
rect 9606 -27883 10006 -27773
rect 9606 -27943 9616 -27883
rect 9676 -27943 9936 -27883
rect 9996 -27943 10006 -27883
rect 9606 -27953 10006 -27943
rect 10062 -27883 10462 -27773
rect 10062 -27943 10072 -27883
rect 10132 -27943 10392 -27883
rect 10452 -27943 10462 -27883
rect 10062 -27953 10462 -27943
rect 10520 -27773 15486 -27771
rect 10520 -27883 10920 -27773
rect 10520 -27943 10530 -27883
rect 10590 -27943 10850 -27883
rect 10910 -27943 10920 -27883
rect 10520 -27953 10920 -27943
rect 10976 -27883 11376 -27773
rect 10976 -27943 10986 -27883
rect 11046 -27943 11306 -27883
rect 11366 -27943 11376 -27883
rect 10976 -27953 11376 -27943
rect 11432 -27883 11832 -27773
rect 11432 -27943 11442 -27883
rect 11502 -27943 11762 -27883
rect 11822 -27943 11832 -27883
rect 11432 -27953 11832 -27943
rect 11890 -27883 12290 -27773
rect 11890 -27943 11900 -27883
rect 11960 -27943 12220 -27883
rect 12280 -27943 12290 -27883
rect 11890 -27953 12290 -27943
rect 12346 -27883 12746 -27773
rect 12346 -27943 12356 -27883
rect 12416 -27943 12676 -27883
rect 12736 -27943 12746 -27883
rect 12346 -27953 12746 -27943
rect 12802 -27883 13202 -27773
rect 12802 -27943 12812 -27883
rect 12872 -27943 13132 -27883
rect 13192 -27943 13202 -27883
rect 12802 -27953 13202 -27943
rect 13260 -27883 13660 -27773
rect 13260 -27943 13270 -27883
rect 13330 -27943 13590 -27883
rect 13650 -27943 13660 -27883
rect 13260 -27953 13660 -27943
rect 13716 -27883 14116 -27773
rect 13716 -27943 13726 -27883
rect 13786 -27943 14046 -27883
rect 14106 -27943 14116 -27883
rect 13716 -27953 14116 -27943
rect 14172 -27883 14572 -27773
rect 14172 -27943 14182 -27883
rect 14242 -27943 14502 -27883
rect 14562 -27943 14572 -27883
rect 14172 -27953 14572 -27943
rect 14630 -27883 15030 -27773
rect 14630 -27943 14640 -27883
rect 14700 -27943 14960 -27883
rect 15020 -27943 15030 -27883
rect 14630 -27953 15030 -27943
rect 15086 -27883 15486 -27773
rect 15086 -27943 15096 -27883
rect 15156 -27943 15416 -27883
rect 15476 -27943 15486 -27883
rect 15086 -27953 15486 -27943
rect 66 -28015 80 -27953
rect 456 -28015 527 -27953
rect 912 -28015 983 -27953
rect 1370 -28015 1441 -27953
rect 1826 -28015 1897 -27953
rect 2282 -28015 2353 -27953
rect 2740 -28015 2810 -27953
rect 3196 -28015 3266 -27953
rect 3652 -28015 3722 -27953
rect 4110 -28015 4180 -27953
rect 4566 -28015 4636 -27953
rect 5022 -28015 5092 -27953
rect 5480 -28015 5550 -27953
rect 5936 -28015 6006 -27953
rect 6392 -28015 6462 -27953
rect 6850 -28015 6920 -27953
rect 7306 -28015 7376 -27953
rect 7762 -28015 7832 -27953
rect 8236 -28015 8306 -27953
rect 8692 -28015 8762 -27953
rect 9150 -28015 9220 -27953
rect 9606 -28015 9676 -27953
rect 10062 -28015 10132 -27953
rect 10520 -28015 10590 -27953
rect 10976 -28015 11046 -27953
rect 11432 -28015 11502 -27953
rect 11890 -28015 11960 -27953
rect 12346 -28015 12416 -27953
rect 12802 -28015 12872 -27953
rect 13260 -28015 13330 -27953
rect 13716 -28015 13786 -27953
rect 14172 -28015 14242 -27953
rect 14630 -28015 14700 -27953
rect 66 -28025 400 -28015
rect 0 -28085 10 -28025
rect 70 -28085 330 -28025
rect 390 -28085 400 -28025
rect 0 -28375 14 -28085
rect 66 -28375 400 -28085
rect 0 -28435 10 -28375
rect 70 -28435 330 -28375
rect 390 -28435 400 -28375
rect 0 -28527 14 -28435
rect 66 -28445 400 -28435
rect 456 -28025 856 -28015
rect 456 -28085 466 -28025
rect 526 -28085 786 -28025
rect 846 -28085 856 -28025
rect 456 -28193 856 -28085
rect 912 -28025 1312 -28015
rect 912 -28085 922 -28025
rect 982 -28085 1242 -28025
rect 1302 -28085 1312 -28025
rect 912 -28193 1312 -28085
rect 1370 -28025 1770 -28015
rect 1370 -28085 1380 -28025
rect 1440 -28085 1700 -28025
rect 1760 -28085 1770 -28025
rect 1370 -28193 1770 -28085
rect 1826 -28025 2226 -28015
rect 1826 -28085 1836 -28025
rect 1896 -28085 2156 -28025
rect 2216 -28085 2226 -28025
rect 1826 -28193 2226 -28085
rect 2282 -28025 2682 -28015
rect 2282 -28085 2292 -28025
rect 2352 -28085 2612 -28025
rect 2672 -28085 2682 -28025
rect 2282 -28193 2682 -28085
rect 2740 -28025 3140 -28015
rect 2740 -28085 2750 -28025
rect 2810 -28085 3070 -28025
rect 3130 -28085 3140 -28025
rect 2740 -28193 3140 -28085
rect 3196 -28025 3596 -28015
rect 3196 -28085 3206 -28025
rect 3266 -28085 3526 -28025
rect 3586 -28085 3596 -28025
rect 3196 -28193 3596 -28085
rect 3652 -28025 4052 -28015
rect 3652 -28085 3662 -28025
rect 3722 -28085 3982 -28025
rect 4042 -28085 4052 -28025
rect 3652 -28193 4052 -28085
rect 4110 -28025 4510 -28015
rect 4110 -28085 4120 -28025
rect 4180 -28085 4440 -28025
rect 4500 -28085 4510 -28025
rect 4110 -28193 4510 -28085
rect 4566 -28025 4966 -28015
rect 4566 -28085 4576 -28025
rect 4636 -28085 4896 -28025
rect 4956 -28085 4966 -28025
rect 4566 -28193 4966 -28085
rect 5022 -28025 5422 -28015
rect 5022 -28085 5032 -28025
rect 5092 -28085 5352 -28025
rect 5412 -28085 5422 -28025
rect 5022 -28193 5422 -28085
rect 5480 -28025 5880 -28015
rect 5480 -28085 5490 -28025
rect 5550 -28085 5810 -28025
rect 5870 -28085 5880 -28025
rect 5480 -28193 5880 -28085
rect 5936 -28025 6336 -28015
rect 5936 -28085 5946 -28025
rect 6006 -28085 6266 -28025
rect 6326 -28085 6336 -28025
rect 5936 -28193 6336 -28085
rect 6392 -28025 6792 -28015
rect 6392 -28085 6402 -28025
rect 6462 -28085 6722 -28025
rect 6782 -28085 6792 -28025
rect 6392 -28193 6792 -28085
rect 6850 -28025 7250 -28015
rect 6850 -28085 6860 -28025
rect 6920 -28085 7180 -28025
rect 7240 -28085 7250 -28025
rect 6850 -28193 7250 -28085
rect 7306 -28025 7706 -28015
rect 7306 -28085 7316 -28025
rect 7376 -28085 7636 -28025
rect 7696 -28085 7706 -28025
rect 7306 -28193 7706 -28085
rect 7762 -28025 8162 -28015
rect 7762 -28085 7772 -28025
rect 7832 -28085 8092 -28025
rect 8152 -28085 8162 -28025
rect 7762 -28193 8162 -28085
rect 8236 -28025 8636 -28015
rect 8236 -28085 8246 -28025
rect 8306 -28085 8566 -28025
rect 8626 -28085 8636 -28025
rect 8236 -28193 8636 -28085
rect 8692 -28025 9092 -28015
rect 8692 -28085 8702 -28025
rect 8762 -28085 9022 -28025
rect 9082 -28085 9092 -28025
rect 8692 -28193 9092 -28085
rect 9150 -28025 9550 -28015
rect 9150 -28085 9160 -28025
rect 9220 -28085 9480 -28025
rect 9540 -28085 9550 -28025
rect 9150 -28193 9550 -28085
rect 9606 -28025 10006 -28015
rect 9606 -28085 9616 -28025
rect 9676 -28085 9936 -28025
rect 9996 -28085 10006 -28025
rect 9606 -28193 10006 -28085
rect 10062 -28025 10462 -28015
rect 10062 -28085 10072 -28025
rect 10132 -28085 10392 -28025
rect 10452 -28085 10462 -28025
rect 10062 -28193 10462 -28085
rect 10520 -28025 10920 -28015
rect 10520 -28085 10530 -28025
rect 10590 -28085 10850 -28025
rect 10910 -28085 10920 -28025
rect 10520 -28193 10920 -28085
rect 10976 -28025 11376 -28015
rect 10976 -28085 10986 -28025
rect 11046 -28085 11306 -28025
rect 11366 -28085 11376 -28025
rect 10976 -28193 11376 -28085
rect 11432 -28025 11832 -28015
rect 11432 -28085 11442 -28025
rect 11502 -28085 11762 -28025
rect 11822 -28085 11832 -28025
rect 11432 -28193 11832 -28085
rect 11890 -28025 12290 -28015
rect 11890 -28085 11900 -28025
rect 11960 -28085 12220 -28025
rect 12280 -28085 12290 -28025
rect 11890 -28193 12290 -28085
rect 12346 -28025 12746 -28015
rect 12346 -28085 12356 -28025
rect 12416 -28085 12676 -28025
rect 12736 -28085 12746 -28025
rect 12346 -28193 12746 -28085
rect 12802 -28025 13202 -28015
rect 12802 -28085 12812 -28025
rect 12872 -28085 13132 -28025
rect 13192 -28085 13202 -28025
rect 12802 -28193 13202 -28085
rect 13260 -28025 13660 -28015
rect 13260 -28085 13270 -28025
rect 13330 -28085 13590 -28025
rect 13650 -28085 13660 -28025
rect 13260 -28193 13660 -28085
rect 13716 -28025 14116 -28015
rect 13716 -28085 13726 -28025
rect 13786 -28085 14046 -28025
rect 14106 -28085 14116 -28025
rect 13716 -28193 14116 -28085
rect 14172 -28025 14572 -28015
rect 14172 -28085 14182 -28025
rect 14242 -28085 14502 -28025
rect 14562 -28085 14572 -28025
rect 14172 -28193 14572 -28085
rect 14630 -28025 15030 -28015
rect 14630 -28085 14640 -28025
rect 14700 -28085 14960 -28025
rect 15020 -28085 15030 -28025
rect 14630 -28193 15030 -28085
rect 15086 -28025 15486 -28015
rect 15086 -28085 15096 -28025
rect 15156 -28085 15416 -28025
rect 15476 -28085 15486 -28025
rect 15086 -28193 15486 -28085
rect 456 -28263 15486 -28193
rect 456 -28265 2682 -28263
rect 456 -28375 856 -28265
rect 456 -28435 466 -28375
rect 526 -28435 786 -28375
rect 846 -28435 856 -28375
rect 456 -28445 856 -28435
rect 912 -28375 1312 -28265
rect 912 -28435 922 -28375
rect 982 -28435 1242 -28375
rect 1302 -28435 1312 -28375
rect 912 -28445 1312 -28435
rect 1370 -28375 1770 -28265
rect 1370 -28435 1380 -28375
rect 1440 -28435 1700 -28375
rect 1760 -28435 1770 -28375
rect 1370 -28445 1770 -28435
rect 1826 -28375 2226 -28265
rect 1826 -28435 1836 -28375
rect 1896 -28435 2156 -28375
rect 2216 -28435 2226 -28375
rect 1826 -28445 2226 -28435
rect 2282 -28375 2682 -28265
rect 2282 -28435 2292 -28375
rect 2352 -28435 2612 -28375
rect 2672 -28435 2682 -28375
rect 2282 -28445 2682 -28435
rect 2740 -28265 10462 -28263
rect 2740 -28375 3140 -28265
rect 2740 -28435 2750 -28375
rect 2810 -28435 3070 -28375
rect 3130 -28435 3140 -28375
rect 2740 -28445 3140 -28435
rect 3196 -28375 3596 -28265
rect 3196 -28435 3206 -28375
rect 3266 -28435 3526 -28375
rect 3586 -28435 3596 -28375
rect 3196 -28445 3596 -28435
rect 3652 -28375 4052 -28265
rect 3652 -28435 3662 -28375
rect 3722 -28435 3982 -28375
rect 4042 -28435 4052 -28375
rect 3652 -28445 4052 -28435
rect 4110 -28375 4510 -28265
rect 4110 -28435 4120 -28375
rect 4180 -28435 4440 -28375
rect 4500 -28435 4510 -28375
rect 4110 -28445 4510 -28435
rect 4566 -28375 4966 -28265
rect 4566 -28435 4576 -28375
rect 4636 -28435 4896 -28375
rect 4956 -28435 4966 -28375
rect 4566 -28445 4966 -28435
rect 5022 -28375 5422 -28265
rect 5022 -28435 5032 -28375
rect 5092 -28435 5352 -28375
rect 5412 -28435 5422 -28375
rect 5022 -28445 5422 -28435
rect 5480 -28375 5880 -28265
rect 5480 -28435 5490 -28375
rect 5550 -28435 5810 -28375
rect 5870 -28435 5880 -28375
rect 5480 -28445 5880 -28435
rect 5936 -28375 6336 -28265
rect 5936 -28435 5946 -28375
rect 6006 -28435 6266 -28375
rect 6326 -28435 6336 -28375
rect 5936 -28445 6336 -28435
rect 6392 -28375 6792 -28265
rect 6392 -28435 6402 -28375
rect 6462 -28435 6722 -28375
rect 6782 -28435 6792 -28375
rect 6392 -28445 6792 -28435
rect 6850 -28375 7250 -28265
rect 6850 -28435 6860 -28375
rect 6920 -28435 7180 -28375
rect 7240 -28435 7250 -28375
rect 6850 -28445 7250 -28435
rect 7306 -28375 7706 -28265
rect 7306 -28435 7316 -28375
rect 7376 -28435 7636 -28375
rect 7696 -28435 7706 -28375
rect 7306 -28445 7706 -28435
rect 7762 -28375 8162 -28265
rect 7762 -28435 7772 -28375
rect 7832 -28435 8092 -28375
rect 8152 -28435 8162 -28375
rect 7762 -28445 8162 -28435
rect 8236 -28375 8636 -28265
rect 8236 -28435 8246 -28375
rect 8306 -28435 8566 -28375
rect 8626 -28435 8636 -28375
rect 8236 -28445 8636 -28435
rect 8692 -28375 9092 -28265
rect 8692 -28435 8702 -28375
rect 8762 -28435 9022 -28375
rect 9082 -28435 9092 -28375
rect 8692 -28445 9092 -28435
rect 9150 -28375 9550 -28265
rect 9150 -28435 9160 -28375
rect 9220 -28435 9480 -28375
rect 9540 -28435 9550 -28375
rect 9150 -28445 9550 -28435
rect 9606 -28375 10006 -28265
rect 9606 -28435 9616 -28375
rect 9676 -28435 9936 -28375
rect 9996 -28435 10006 -28375
rect 9606 -28445 10006 -28435
rect 10062 -28375 10462 -28265
rect 10062 -28435 10072 -28375
rect 10132 -28435 10392 -28375
rect 10452 -28435 10462 -28375
rect 10062 -28445 10462 -28435
rect 10520 -28265 15486 -28263
rect 10520 -28375 10920 -28265
rect 10520 -28435 10530 -28375
rect 10590 -28435 10850 -28375
rect 10910 -28435 10920 -28375
rect 10520 -28445 10920 -28435
rect 10976 -28375 11376 -28265
rect 10976 -28435 10986 -28375
rect 11046 -28435 11306 -28375
rect 11366 -28435 11376 -28375
rect 10976 -28445 11376 -28435
rect 11432 -28375 11832 -28265
rect 11432 -28435 11442 -28375
rect 11502 -28435 11762 -28375
rect 11822 -28435 11832 -28375
rect 11432 -28445 11832 -28435
rect 11890 -28375 12290 -28265
rect 11890 -28435 11900 -28375
rect 11960 -28435 12220 -28375
rect 12280 -28435 12290 -28375
rect 11890 -28445 12290 -28435
rect 12346 -28375 12746 -28265
rect 12346 -28435 12356 -28375
rect 12416 -28435 12676 -28375
rect 12736 -28435 12746 -28375
rect 12346 -28445 12746 -28435
rect 12802 -28375 13202 -28265
rect 12802 -28435 12812 -28375
rect 12872 -28435 13132 -28375
rect 13192 -28435 13202 -28375
rect 12802 -28445 13202 -28435
rect 13260 -28375 13660 -28265
rect 13260 -28435 13270 -28375
rect 13330 -28435 13590 -28375
rect 13650 -28435 13660 -28375
rect 13260 -28445 13660 -28435
rect 13716 -28375 14116 -28265
rect 13716 -28435 13726 -28375
rect 13786 -28435 14046 -28375
rect 14106 -28435 14116 -28375
rect 13716 -28445 14116 -28435
rect 14172 -28375 14572 -28265
rect 14172 -28435 14182 -28375
rect 14242 -28435 14502 -28375
rect 14562 -28435 14572 -28375
rect 14172 -28445 14572 -28435
rect 14630 -28375 15030 -28265
rect 14630 -28435 14640 -28375
rect 14700 -28435 14960 -28375
rect 15020 -28435 15030 -28375
rect 14630 -28445 15030 -28435
rect 15086 -28375 15486 -28265
rect 15086 -28435 15096 -28375
rect 15156 -28435 15416 -28375
rect 15476 -28435 15486 -28375
rect 15086 -28445 15486 -28435
rect 66 -28517 80 -28445
rect 456 -28517 526 -28445
rect 912 -28517 983 -28445
rect 1370 -28517 1441 -28445
rect 1826 -28517 1897 -28445
rect 2282 -28517 2353 -28445
rect 2740 -28517 2811 -28445
rect 3196 -28517 3267 -28445
rect 3652 -28517 3723 -28445
rect 4110 -28517 4181 -28445
rect 4566 -28517 4637 -28445
rect 5022 -28517 5093 -28445
rect 5480 -28517 5551 -28445
rect 5936 -28517 6007 -28445
rect 6392 -28517 6463 -28445
rect 6850 -28517 6921 -28445
rect 7306 -28517 7377 -28445
rect 7762 -28517 7833 -28445
rect 8236 -28517 8307 -28445
rect 8692 -28517 8763 -28445
rect 9150 -28517 9221 -28445
rect 9606 -28517 9677 -28445
rect 10062 -28517 10133 -28445
rect 10520 -28517 10591 -28445
rect 10976 -28517 11047 -28445
rect 11432 -28517 11503 -28445
rect 11890 -28517 11961 -28445
rect 12346 -28517 12417 -28445
rect 12802 -28517 12873 -28445
rect 13260 -28517 13331 -28445
rect 13716 -28517 13787 -28445
rect 14172 -28517 14243 -28445
rect 14630 -28517 14701 -28445
rect 66 -28527 400 -28517
rect 0 -28587 10 -28527
rect 70 -28587 330 -28527
rect 390 -28587 400 -28527
rect 0 -28877 14 -28587
rect 66 -28877 400 -28587
rect 0 -28937 10 -28877
rect 70 -28937 330 -28877
rect 390 -28937 400 -28877
rect 0 -29021 14 -28937
rect 66 -28947 400 -28937
rect 456 -28527 856 -28517
rect 456 -28587 466 -28527
rect 526 -28587 786 -28527
rect 846 -28587 856 -28527
rect 456 -28696 856 -28587
rect 912 -28527 1312 -28517
rect 912 -28587 922 -28527
rect 982 -28587 1242 -28527
rect 1302 -28587 1312 -28527
rect 912 -28696 1312 -28587
rect 1370 -28527 1770 -28517
rect 1370 -28587 1380 -28527
rect 1440 -28587 1700 -28527
rect 1760 -28587 1770 -28527
rect 1370 -28696 1770 -28587
rect 1826 -28527 2226 -28517
rect 1826 -28587 1836 -28527
rect 1896 -28587 2156 -28527
rect 2216 -28587 2226 -28527
rect 1826 -28696 2226 -28587
rect 2282 -28527 2682 -28517
rect 2282 -28587 2292 -28527
rect 2352 -28587 2612 -28527
rect 2672 -28587 2682 -28527
rect 2282 -28696 2682 -28587
rect 2740 -28527 3140 -28517
rect 2740 -28587 2750 -28527
rect 2810 -28587 3070 -28527
rect 3130 -28587 3140 -28527
rect 2740 -28696 3140 -28587
rect 3196 -28527 3596 -28517
rect 3196 -28587 3206 -28527
rect 3266 -28587 3526 -28527
rect 3586 -28587 3596 -28527
rect 3196 -28696 3596 -28587
rect 3652 -28527 4052 -28517
rect 3652 -28587 3662 -28527
rect 3722 -28587 3982 -28527
rect 4042 -28587 4052 -28527
rect 3652 -28696 4052 -28587
rect 4110 -28527 4510 -28517
rect 4110 -28587 4120 -28527
rect 4180 -28587 4440 -28527
rect 4500 -28587 4510 -28527
rect 4110 -28696 4510 -28587
rect 4566 -28527 4966 -28517
rect 4566 -28587 4576 -28527
rect 4636 -28587 4896 -28527
rect 4956 -28587 4966 -28527
rect 4566 -28696 4966 -28587
rect 5022 -28527 5422 -28517
rect 5022 -28587 5032 -28527
rect 5092 -28587 5352 -28527
rect 5412 -28587 5422 -28527
rect 5022 -28696 5422 -28587
rect 5480 -28527 5880 -28517
rect 5480 -28587 5490 -28527
rect 5550 -28587 5810 -28527
rect 5870 -28587 5880 -28527
rect 5480 -28696 5880 -28587
rect 5936 -28527 6336 -28517
rect 5936 -28587 5946 -28527
rect 6006 -28587 6266 -28527
rect 6326 -28587 6336 -28527
rect 5936 -28696 6336 -28587
rect 6392 -28527 6792 -28517
rect 6392 -28587 6402 -28527
rect 6462 -28587 6722 -28527
rect 6782 -28587 6792 -28527
rect 6392 -28696 6792 -28587
rect 6850 -28527 7250 -28517
rect 6850 -28587 6860 -28527
rect 6920 -28587 7180 -28527
rect 7240 -28587 7250 -28527
rect 6850 -28696 7250 -28587
rect 7306 -28527 7706 -28517
rect 7306 -28587 7316 -28527
rect 7376 -28587 7636 -28527
rect 7696 -28587 7706 -28527
rect 7306 -28696 7706 -28587
rect 7762 -28527 8162 -28517
rect 7762 -28587 7772 -28527
rect 7832 -28587 8092 -28527
rect 8152 -28587 8162 -28527
rect 7762 -28696 8162 -28587
rect 8236 -28527 8636 -28517
rect 8236 -28587 8246 -28527
rect 8306 -28587 8566 -28527
rect 8626 -28587 8636 -28527
rect 8236 -28696 8636 -28587
rect 8692 -28527 9092 -28517
rect 8692 -28587 8702 -28527
rect 8762 -28587 9022 -28527
rect 9082 -28587 9092 -28527
rect 8692 -28696 9092 -28587
rect 9150 -28527 9550 -28517
rect 9150 -28587 9160 -28527
rect 9220 -28587 9480 -28527
rect 9540 -28587 9550 -28527
rect 9150 -28696 9550 -28587
rect 9606 -28527 10006 -28517
rect 9606 -28587 9616 -28527
rect 9676 -28587 9936 -28527
rect 9996 -28587 10006 -28527
rect 9606 -28696 10006 -28587
rect 10062 -28527 10462 -28517
rect 10062 -28587 10072 -28527
rect 10132 -28587 10392 -28527
rect 10452 -28587 10462 -28527
rect 10062 -28696 10462 -28587
rect 10520 -28527 10920 -28517
rect 10520 -28587 10530 -28527
rect 10590 -28587 10850 -28527
rect 10910 -28587 10920 -28527
rect 10520 -28696 10920 -28587
rect 10976 -28527 11376 -28517
rect 10976 -28587 10986 -28527
rect 11046 -28587 11306 -28527
rect 11366 -28587 11376 -28527
rect 10976 -28696 11376 -28587
rect 11432 -28527 11832 -28517
rect 11432 -28587 11442 -28527
rect 11502 -28587 11762 -28527
rect 11822 -28587 11832 -28527
rect 11432 -28696 11832 -28587
rect 11890 -28527 12290 -28517
rect 11890 -28587 11900 -28527
rect 11960 -28587 12220 -28527
rect 12280 -28587 12290 -28527
rect 11890 -28696 12290 -28587
rect 12346 -28527 12746 -28517
rect 12346 -28587 12356 -28527
rect 12416 -28587 12676 -28527
rect 12736 -28587 12746 -28527
rect 12346 -28696 12746 -28587
rect 12802 -28527 13202 -28517
rect 12802 -28587 12812 -28527
rect 12872 -28587 13132 -28527
rect 13192 -28587 13202 -28527
rect 12802 -28696 13202 -28587
rect 13260 -28527 13660 -28517
rect 13260 -28587 13270 -28527
rect 13330 -28587 13590 -28527
rect 13650 -28587 13660 -28527
rect 13260 -28696 13660 -28587
rect 13716 -28527 14116 -28517
rect 13716 -28587 13726 -28527
rect 13786 -28587 14046 -28527
rect 14106 -28587 14116 -28527
rect 13716 -28696 14116 -28587
rect 14172 -28527 14572 -28517
rect 14172 -28587 14182 -28527
rect 14242 -28587 14502 -28527
rect 14562 -28587 14572 -28527
rect 14172 -28696 14572 -28587
rect 14630 -28527 15030 -28517
rect 14630 -28587 14640 -28527
rect 14700 -28587 14960 -28527
rect 15020 -28587 15030 -28527
rect 14630 -28696 15030 -28587
rect 15086 -28527 15486 -28517
rect 15086 -28587 15096 -28527
rect 15156 -28587 15416 -28527
rect 15476 -28587 15486 -28527
rect 15086 -28696 15486 -28587
rect 456 -28766 15486 -28696
rect 456 -28877 856 -28766
rect 456 -28937 466 -28877
rect 526 -28937 786 -28877
rect 846 -28937 856 -28877
rect 456 -28947 856 -28937
rect 912 -28877 1312 -28766
rect 912 -28937 922 -28877
rect 982 -28937 1242 -28877
rect 1302 -28937 1312 -28877
rect 912 -28947 1312 -28937
rect 1370 -28877 1770 -28766
rect 1370 -28937 1380 -28877
rect 1440 -28937 1700 -28877
rect 1760 -28937 1770 -28877
rect 1370 -28947 1770 -28937
rect 1826 -28877 2226 -28766
rect 1826 -28937 1836 -28877
rect 1896 -28937 2156 -28877
rect 2216 -28937 2226 -28877
rect 1826 -28947 2226 -28937
rect 2282 -28877 2682 -28766
rect 2282 -28937 2292 -28877
rect 2352 -28937 2612 -28877
rect 2672 -28937 2682 -28877
rect 2282 -28947 2682 -28937
rect 2740 -28877 3140 -28766
rect 2740 -28937 2750 -28877
rect 2810 -28937 3070 -28877
rect 3130 -28937 3140 -28877
rect 2740 -28947 3140 -28937
rect 3196 -28877 3596 -28766
rect 3196 -28937 3206 -28877
rect 3266 -28937 3526 -28877
rect 3586 -28937 3596 -28877
rect 3196 -28947 3596 -28937
rect 3652 -28877 4052 -28766
rect 3652 -28937 3662 -28877
rect 3722 -28937 3982 -28877
rect 4042 -28937 4052 -28877
rect 3652 -28947 4052 -28937
rect 4110 -28877 4510 -28766
rect 4110 -28937 4120 -28877
rect 4180 -28937 4440 -28877
rect 4500 -28937 4510 -28877
rect 4110 -28947 4510 -28937
rect 4566 -28877 4966 -28766
rect 4566 -28937 4576 -28877
rect 4636 -28937 4896 -28877
rect 4956 -28937 4966 -28877
rect 4566 -28947 4966 -28937
rect 5022 -28877 5422 -28766
rect 5022 -28937 5032 -28877
rect 5092 -28937 5352 -28877
rect 5412 -28937 5422 -28877
rect 5022 -28947 5422 -28937
rect 5480 -28877 5880 -28766
rect 5480 -28937 5490 -28877
rect 5550 -28937 5810 -28877
rect 5870 -28937 5880 -28877
rect 5480 -28947 5880 -28937
rect 5936 -28877 6336 -28766
rect 5936 -28937 5946 -28877
rect 6006 -28937 6266 -28877
rect 6326 -28937 6336 -28877
rect 5936 -28947 6336 -28937
rect 6392 -28877 6792 -28766
rect 6392 -28937 6402 -28877
rect 6462 -28937 6722 -28877
rect 6782 -28937 6792 -28877
rect 6392 -28947 6792 -28937
rect 6850 -28877 7250 -28766
rect 6850 -28937 6860 -28877
rect 6920 -28937 7180 -28877
rect 7240 -28937 7250 -28877
rect 6850 -28947 7250 -28937
rect 7306 -28877 7706 -28766
rect 7306 -28937 7316 -28877
rect 7376 -28937 7636 -28877
rect 7696 -28937 7706 -28877
rect 7306 -28947 7706 -28937
rect 7762 -28877 8162 -28766
rect 7762 -28937 7772 -28877
rect 7832 -28937 8092 -28877
rect 8152 -28937 8162 -28877
rect 7762 -28947 8162 -28937
rect 8236 -28877 8636 -28766
rect 8236 -28937 8246 -28877
rect 8306 -28937 8566 -28877
rect 8626 -28937 8636 -28877
rect 8236 -28947 8636 -28937
rect 8692 -28877 9092 -28766
rect 8692 -28937 8702 -28877
rect 8762 -28937 9022 -28877
rect 9082 -28937 9092 -28877
rect 8692 -28947 9092 -28937
rect 9150 -28877 9550 -28766
rect 9150 -28937 9160 -28877
rect 9220 -28937 9480 -28877
rect 9540 -28937 9550 -28877
rect 9150 -28947 9550 -28937
rect 9606 -28877 10006 -28766
rect 9606 -28937 9616 -28877
rect 9676 -28937 9936 -28877
rect 9996 -28937 10006 -28877
rect 9606 -28947 10006 -28937
rect 10062 -28877 10462 -28766
rect 10062 -28937 10072 -28877
rect 10132 -28937 10392 -28877
rect 10452 -28937 10462 -28877
rect 10062 -28947 10462 -28937
rect 10520 -28877 10920 -28766
rect 10520 -28937 10530 -28877
rect 10590 -28937 10850 -28877
rect 10910 -28937 10920 -28877
rect 10520 -28947 10920 -28937
rect 10976 -28877 11376 -28766
rect 10976 -28937 10986 -28877
rect 11046 -28937 11306 -28877
rect 11366 -28937 11376 -28877
rect 10976 -28947 11376 -28937
rect 11432 -28877 11832 -28766
rect 11432 -28937 11442 -28877
rect 11502 -28937 11762 -28877
rect 11822 -28937 11832 -28877
rect 11432 -28947 11832 -28937
rect 11890 -28877 12290 -28766
rect 11890 -28937 11900 -28877
rect 11960 -28937 12220 -28877
rect 12280 -28937 12290 -28877
rect 11890 -28947 12290 -28937
rect 12346 -28877 12746 -28766
rect 12346 -28937 12356 -28877
rect 12416 -28937 12676 -28877
rect 12736 -28937 12746 -28877
rect 12346 -28947 12746 -28937
rect 12802 -28877 13202 -28766
rect 12802 -28937 12812 -28877
rect 12872 -28937 13132 -28877
rect 13192 -28937 13202 -28877
rect 12802 -28947 13202 -28937
rect 13260 -28877 13660 -28766
rect 13260 -28937 13270 -28877
rect 13330 -28937 13590 -28877
rect 13650 -28937 13660 -28877
rect 13260 -28947 13660 -28937
rect 13716 -28877 14116 -28766
rect 13716 -28937 13726 -28877
rect 13786 -28937 14046 -28877
rect 14106 -28937 14116 -28877
rect 13716 -28947 14116 -28937
rect 14172 -28877 14572 -28766
rect 14172 -28937 14182 -28877
rect 14242 -28937 14502 -28877
rect 14562 -28937 14572 -28877
rect 14172 -28947 14572 -28937
rect 14630 -28877 15030 -28766
rect 14630 -28937 14640 -28877
rect 14700 -28937 14960 -28877
rect 15020 -28937 15030 -28877
rect 14630 -28947 15030 -28937
rect 15086 -28877 15486 -28766
rect 15086 -28937 15096 -28877
rect 15156 -28937 15416 -28877
rect 15476 -28937 15486 -28877
rect 15086 -28947 15486 -28937
rect 66 -29011 80 -28947
rect 456 -29011 526 -28947
rect 912 -29011 982 -28947
rect 1370 -29011 1440 -28947
rect 1826 -29011 1896 -28947
rect 2282 -29011 2352 -28947
rect 2740 -29011 2810 -28947
rect 3196 -29011 3266 -28947
rect 3652 -29011 3722 -28947
rect 4110 -29011 4180 -28947
rect 4566 -29011 4636 -28947
rect 5022 -29011 5092 -28947
rect 5480 -29011 5550 -28947
rect 5936 -29011 6006 -28947
rect 6392 -29011 6462 -28947
rect 6850 -29011 6920 -28947
rect 7306 -29011 7376 -28947
rect 7762 -29011 7832 -28947
rect 8236 -29011 8306 -28947
rect 8692 -29011 8762 -28947
rect 9150 -29011 9220 -28947
rect 9606 -29011 9676 -28947
rect 10062 -29011 10132 -28947
rect 10520 -29011 10590 -28947
rect 10976 -29011 11047 -28947
rect 11432 -29011 11503 -28947
rect 11890 -29011 11961 -28947
rect 12346 -29011 12417 -28947
rect 12802 -29011 12873 -28947
rect 13260 -29011 13331 -28947
rect 13716 -29011 13787 -28947
rect 14172 -29011 14243 -28947
rect 14630 -29011 14701 -28947
rect 66 -29021 400 -29011
rect 0 -29081 10 -29021
rect 70 -29081 330 -29021
rect 390 -29081 400 -29021
rect 0 -29371 14 -29081
rect 66 -29371 400 -29081
rect 0 -29431 10 -29371
rect 70 -29431 330 -29371
rect 390 -29431 400 -29371
rect 0 -29513 14 -29431
rect 66 -29441 400 -29431
rect 456 -29021 856 -29011
rect 456 -29081 466 -29021
rect 526 -29081 786 -29021
rect 846 -29081 856 -29021
rect 456 -29191 856 -29081
rect 912 -29021 1312 -29011
rect 912 -29081 922 -29021
rect 982 -29081 1242 -29021
rect 1302 -29081 1312 -29021
rect 912 -29191 1312 -29081
rect 1370 -29021 1770 -29011
rect 1370 -29081 1380 -29021
rect 1440 -29081 1700 -29021
rect 1760 -29081 1770 -29021
rect 1370 -29191 1770 -29081
rect 1826 -29021 2226 -29011
rect 1826 -29081 1836 -29021
rect 1896 -29081 2156 -29021
rect 2216 -29081 2226 -29021
rect 1826 -29191 2226 -29081
rect 2282 -29021 2682 -29011
rect 2282 -29081 2292 -29021
rect 2352 -29081 2612 -29021
rect 2672 -29081 2682 -29021
rect 2282 -29191 2682 -29081
rect 456 -29192 2682 -29191
rect 2740 -29021 3140 -29011
rect 2740 -29081 2750 -29021
rect 2810 -29081 3070 -29021
rect 3130 -29081 3140 -29021
rect 2740 -29191 3140 -29081
rect 3196 -29021 3596 -29011
rect 3196 -29081 3206 -29021
rect 3266 -29081 3526 -29021
rect 3586 -29081 3596 -29021
rect 3196 -29191 3596 -29081
rect 3652 -29021 4052 -29011
rect 3652 -29081 3662 -29021
rect 3722 -29081 3982 -29021
rect 4042 -29081 4052 -29021
rect 3652 -29191 4052 -29081
rect 4110 -29021 4510 -29011
rect 4110 -29081 4120 -29021
rect 4180 -29081 4440 -29021
rect 4500 -29081 4510 -29021
rect 4110 -29191 4510 -29081
rect 4566 -29021 4966 -29011
rect 4566 -29081 4576 -29021
rect 4636 -29081 4896 -29021
rect 4956 -29081 4966 -29021
rect 4566 -29191 4966 -29081
rect 5022 -29021 5422 -29011
rect 5022 -29081 5032 -29021
rect 5092 -29081 5352 -29021
rect 5412 -29081 5422 -29021
rect 5022 -29191 5422 -29081
rect 5480 -29021 5880 -29011
rect 5480 -29081 5490 -29021
rect 5550 -29081 5810 -29021
rect 5870 -29081 5880 -29021
rect 5480 -29191 5880 -29081
rect 5936 -29021 6336 -29011
rect 5936 -29081 5946 -29021
rect 6006 -29081 6266 -29021
rect 6326 -29081 6336 -29021
rect 5936 -29191 6336 -29081
rect 6392 -29021 6792 -29011
rect 6392 -29081 6402 -29021
rect 6462 -29081 6722 -29021
rect 6782 -29081 6792 -29021
rect 6392 -29191 6792 -29081
rect 6850 -29021 7250 -29011
rect 6850 -29081 6860 -29021
rect 6920 -29081 7180 -29021
rect 7240 -29081 7250 -29021
rect 6850 -29191 7250 -29081
rect 7306 -29021 7706 -29011
rect 7306 -29081 7316 -29021
rect 7376 -29081 7636 -29021
rect 7696 -29081 7706 -29021
rect 7306 -29191 7706 -29081
rect 7762 -29021 8162 -29011
rect 7762 -29081 7772 -29021
rect 7832 -29081 8092 -29021
rect 8152 -29081 8162 -29021
rect 7762 -29191 8162 -29081
rect 8236 -29021 8636 -29011
rect 8236 -29081 8246 -29021
rect 8306 -29081 8566 -29021
rect 8626 -29081 8636 -29021
rect 8236 -29191 8636 -29081
rect 8692 -29021 9092 -29011
rect 8692 -29081 8702 -29021
rect 8762 -29081 9022 -29021
rect 9082 -29081 9092 -29021
rect 8692 -29191 9092 -29081
rect 9150 -29021 9550 -29011
rect 9150 -29081 9160 -29021
rect 9220 -29081 9480 -29021
rect 9540 -29081 9550 -29021
rect 9150 -29191 9550 -29081
rect 9606 -29021 10006 -29011
rect 9606 -29081 9616 -29021
rect 9676 -29081 9936 -29021
rect 9996 -29081 10006 -29021
rect 9606 -29191 10006 -29081
rect 10062 -29021 10462 -29011
rect 10062 -29081 10072 -29021
rect 10132 -29081 10392 -29021
rect 10452 -29081 10462 -29021
rect 10062 -29191 10462 -29081
rect 2740 -29192 10462 -29191
rect 10520 -29021 10920 -29011
rect 10520 -29081 10530 -29021
rect 10590 -29081 10850 -29021
rect 10910 -29081 10920 -29021
rect 10520 -29191 10920 -29081
rect 10976 -29021 11376 -29011
rect 10976 -29081 10986 -29021
rect 11046 -29081 11306 -29021
rect 11366 -29081 11376 -29021
rect 10976 -29191 11376 -29081
rect 11432 -29021 11832 -29011
rect 11432 -29081 11442 -29021
rect 11502 -29081 11762 -29021
rect 11822 -29081 11832 -29021
rect 11432 -29191 11832 -29081
rect 11890 -29021 12290 -29011
rect 11890 -29081 11900 -29021
rect 11960 -29081 12220 -29021
rect 12280 -29081 12290 -29021
rect 11890 -29191 12290 -29081
rect 12346 -29021 12746 -29011
rect 12346 -29081 12356 -29021
rect 12416 -29081 12676 -29021
rect 12736 -29081 12746 -29021
rect 12346 -29191 12746 -29081
rect 12802 -29021 13202 -29011
rect 12802 -29081 12812 -29021
rect 12872 -29081 13132 -29021
rect 13192 -29081 13202 -29021
rect 12802 -29191 13202 -29081
rect 13260 -29021 13660 -29011
rect 13260 -29081 13270 -29021
rect 13330 -29081 13590 -29021
rect 13650 -29081 13660 -29021
rect 13260 -29191 13660 -29081
rect 13716 -29021 14116 -29011
rect 13716 -29081 13726 -29021
rect 13786 -29081 14046 -29021
rect 14106 -29081 14116 -29021
rect 13716 -29191 14116 -29081
rect 14172 -29021 14572 -29011
rect 14172 -29081 14182 -29021
rect 14242 -29081 14502 -29021
rect 14562 -29081 14572 -29021
rect 14172 -29191 14572 -29081
rect 14630 -29021 15030 -29011
rect 14630 -29081 14640 -29021
rect 14700 -29081 14960 -29021
rect 15020 -29081 15030 -29021
rect 14630 -29191 15030 -29081
rect 15086 -29021 15486 -29011
rect 15086 -29081 15096 -29021
rect 15156 -29081 15416 -29021
rect 15476 -29081 15486 -29021
rect 15086 -29191 15486 -29081
rect 10520 -29192 15486 -29191
rect 456 -29262 15486 -29192
rect 456 -29371 856 -29262
rect 456 -29431 466 -29371
rect 526 -29431 786 -29371
rect 846 -29431 856 -29371
rect 456 -29441 856 -29431
rect 912 -29371 1312 -29262
rect 912 -29431 922 -29371
rect 982 -29431 1242 -29371
rect 1302 -29431 1312 -29371
rect 912 -29441 1312 -29431
rect 1370 -29371 1770 -29262
rect 1370 -29431 1380 -29371
rect 1440 -29431 1700 -29371
rect 1760 -29431 1770 -29371
rect 1370 -29441 1770 -29431
rect 1826 -29371 2226 -29262
rect 1826 -29431 1836 -29371
rect 1896 -29431 2156 -29371
rect 2216 -29431 2226 -29371
rect 1826 -29441 2226 -29431
rect 2282 -29371 2682 -29262
rect 2282 -29431 2292 -29371
rect 2352 -29431 2612 -29371
rect 2672 -29431 2682 -29371
rect 2282 -29441 2682 -29431
rect 2740 -29371 3140 -29262
rect 2740 -29431 2750 -29371
rect 2810 -29431 3070 -29371
rect 3130 -29431 3140 -29371
rect 2740 -29441 3140 -29431
rect 3196 -29371 3596 -29262
rect 3196 -29431 3206 -29371
rect 3266 -29431 3526 -29371
rect 3586 -29431 3596 -29371
rect 3196 -29441 3596 -29431
rect 3652 -29371 4052 -29262
rect 3652 -29431 3662 -29371
rect 3722 -29431 3982 -29371
rect 4042 -29431 4052 -29371
rect 3652 -29441 4052 -29431
rect 4110 -29371 4510 -29262
rect 4110 -29431 4120 -29371
rect 4180 -29431 4440 -29371
rect 4500 -29431 4510 -29371
rect 4110 -29441 4510 -29431
rect 4566 -29371 4966 -29262
rect 4566 -29431 4576 -29371
rect 4636 -29431 4896 -29371
rect 4956 -29431 4966 -29371
rect 4566 -29441 4966 -29431
rect 5022 -29371 5422 -29262
rect 5022 -29431 5032 -29371
rect 5092 -29431 5352 -29371
rect 5412 -29431 5422 -29371
rect 5022 -29441 5422 -29431
rect 5480 -29371 5880 -29262
rect 5480 -29431 5490 -29371
rect 5550 -29431 5810 -29371
rect 5870 -29431 5880 -29371
rect 5480 -29441 5880 -29431
rect 5936 -29371 6336 -29262
rect 5936 -29431 5946 -29371
rect 6006 -29431 6266 -29371
rect 6326 -29431 6336 -29371
rect 5936 -29441 6336 -29431
rect 6392 -29371 6792 -29262
rect 6392 -29431 6402 -29371
rect 6462 -29431 6722 -29371
rect 6782 -29431 6792 -29371
rect 6392 -29441 6792 -29431
rect 6850 -29371 7250 -29262
rect 6850 -29431 6860 -29371
rect 6920 -29431 7180 -29371
rect 7240 -29431 7250 -29371
rect 6850 -29441 7250 -29431
rect 7306 -29371 7706 -29262
rect 7306 -29431 7316 -29371
rect 7376 -29431 7636 -29371
rect 7696 -29431 7706 -29371
rect 7306 -29441 7706 -29431
rect 7762 -29371 8162 -29262
rect 7762 -29431 7772 -29371
rect 7832 -29431 8092 -29371
rect 8152 -29431 8162 -29371
rect 7762 -29441 8162 -29431
rect 8236 -29371 8636 -29262
rect 8236 -29431 8246 -29371
rect 8306 -29431 8566 -29371
rect 8626 -29431 8636 -29371
rect 8236 -29441 8636 -29431
rect 8692 -29371 9092 -29262
rect 8692 -29431 8702 -29371
rect 8762 -29431 9022 -29371
rect 9082 -29431 9092 -29371
rect 8692 -29441 9092 -29431
rect 9150 -29371 9550 -29262
rect 9150 -29431 9160 -29371
rect 9220 -29431 9480 -29371
rect 9540 -29431 9550 -29371
rect 9150 -29441 9550 -29431
rect 9606 -29371 10006 -29262
rect 9606 -29431 9616 -29371
rect 9676 -29431 9936 -29371
rect 9996 -29431 10006 -29371
rect 9606 -29441 10006 -29431
rect 10062 -29371 10462 -29262
rect 10062 -29431 10072 -29371
rect 10132 -29431 10392 -29371
rect 10452 -29431 10462 -29371
rect 10062 -29441 10462 -29431
rect 10520 -29371 10920 -29262
rect 10520 -29431 10530 -29371
rect 10590 -29431 10850 -29371
rect 10910 -29431 10920 -29371
rect 10520 -29441 10920 -29431
rect 10976 -29371 11376 -29262
rect 10976 -29431 10986 -29371
rect 11046 -29431 11306 -29371
rect 11366 -29431 11376 -29371
rect 10976 -29441 11376 -29431
rect 11432 -29371 11832 -29262
rect 11432 -29431 11442 -29371
rect 11502 -29431 11762 -29371
rect 11822 -29431 11832 -29371
rect 11432 -29441 11832 -29431
rect 11890 -29371 12290 -29262
rect 11890 -29431 11900 -29371
rect 11960 -29431 12220 -29371
rect 12280 -29431 12290 -29371
rect 11890 -29441 12290 -29431
rect 12346 -29371 12746 -29262
rect 12346 -29431 12356 -29371
rect 12416 -29431 12676 -29371
rect 12736 -29431 12746 -29371
rect 12346 -29441 12746 -29431
rect 12802 -29371 13202 -29262
rect 12802 -29431 12812 -29371
rect 12872 -29431 13132 -29371
rect 13192 -29431 13202 -29371
rect 12802 -29441 13202 -29431
rect 13260 -29371 13660 -29262
rect 13260 -29431 13270 -29371
rect 13330 -29431 13590 -29371
rect 13650 -29431 13660 -29371
rect 13260 -29441 13660 -29431
rect 13716 -29371 14116 -29262
rect 13716 -29431 13726 -29371
rect 13786 -29431 14046 -29371
rect 14106 -29431 14116 -29371
rect 13716 -29441 14116 -29431
rect 14172 -29371 14572 -29262
rect 14172 -29431 14182 -29371
rect 14242 -29431 14502 -29371
rect 14562 -29431 14572 -29371
rect 14172 -29441 14572 -29431
rect 14630 -29371 15030 -29262
rect 14630 -29431 14640 -29371
rect 14700 -29431 14960 -29371
rect 15020 -29431 15030 -29371
rect 14630 -29441 15030 -29431
rect 15086 -29371 15486 -29262
rect 15086 -29431 15096 -29371
rect 15156 -29431 15416 -29371
rect 15476 -29431 15486 -29371
rect 15086 -29441 15486 -29431
rect 66 -29503 80 -29441
rect 456 -29503 527 -29441
rect 912 -29503 983 -29441
rect 1370 -29503 1441 -29441
rect 1826 -29503 1897 -29441
rect 2282 -29503 2353 -29441
rect 2740 -29503 2810 -29441
rect 3196 -29503 3266 -29441
rect 3652 -29503 3722 -29441
rect 4110 -29503 4180 -29441
rect 4566 -29503 4636 -29441
rect 5022 -29503 5092 -29441
rect 5480 -29503 5550 -29441
rect 5936 -29503 6006 -29441
rect 6392 -29503 6462 -29441
rect 6850 -29503 6920 -29441
rect 7306 -29503 7376 -29441
rect 7762 -29503 7832 -29441
rect 8236 -29503 8306 -29441
rect 8692 -29503 8762 -29441
rect 9150 -29503 9220 -29441
rect 9606 -29503 9676 -29441
rect 10062 -29503 10132 -29441
rect 10520 -29503 10590 -29441
rect 10976 -29503 11046 -29441
rect 11432 -29503 11502 -29441
rect 11890 -29503 11960 -29441
rect 12346 -29503 12416 -29441
rect 12802 -29503 12872 -29441
rect 13260 -29503 13330 -29441
rect 13716 -29503 13786 -29441
rect 14172 -29503 14242 -29441
rect 14630 -29503 14700 -29441
rect 66 -29513 400 -29503
rect 0 -29573 10 -29513
rect 70 -29573 330 -29513
rect 390 -29573 400 -29513
rect 0 -29863 14 -29573
rect 66 -29863 400 -29573
rect 0 -29923 10 -29863
rect 70 -29923 330 -29863
rect 390 -29923 400 -29863
rect 0 -30015 14 -29923
rect 66 -29933 400 -29923
rect 456 -29513 856 -29503
rect 456 -29573 466 -29513
rect 526 -29573 786 -29513
rect 846 -29573 856 -29513
rect 456 -29683 856 -29573
rect 912 -29513 1312 -29503
rect 912 -29573 922 -29513
rect 982 -29573 1242 -29513
rect 1302 -29573 1312 -29513
rect 912 -29683 1312 -29573
rect 1370 -29513 1770 -29503
rect 1370 -29573 1380 -29513
rect 1440 -29573 1700 -29513
rect 1760 -29573 1770 -29513
rect 1370 -29683 1770 -29573
rect 1826 -29513 2226 -29503
rect 1826 -29573 1836 -29513
rect 1896 -29573 2156 -29513
rect 2216 -29573 2226 -29513
rect 1826 -29683 2226 -29573
rect 2282 -29513 2682 -29503
rect 2282 -29573 2292 -29513
rect 2352 -29573 2612 -29513
rect 2672 -29573 2682 -29513
rect 2282 -29683 2682 -29573
rect 2740 -29513 3140 -29503
rect 2740 -29573 2750 -29513
rect 2810 -29573 3070 -29513
rect 3130 -29573 3140 -29513
rect 2740 -29683 3140 -29573
rect 3196 -29513 3596 -29503
rect 3196 -29573 3206 -29513
rect 3266 -29573 3526 -29513
rect 3586 -29573 3596 -29513
rect 3196 -29683 3596 -29573
rect 3652 -29513 4052 -29503
rect 3652 -29573 3662 -29513
rect 3722 -29573 3982 -29513
rect 4042 -29573 4052 -29513
rect 3652 -29683 4052 -29573
rect 4110 -29513 4510 -29503
rect 4110 -29573 4120 -29513
rect 4180 -29573 4440 -29513
rect 4500 -29573 4510 -29513
rect 4110 -29683 4510 -29573
rect 4566 -29513 4966 -29503
rect 4566 -29573 4576 -29513
rect 4636 -29573 4896 -29513
rect 4956 -29573 4966 -29513
rect 4566 -29683 4966 -29573
rect 5022 -29513 5422 -29503
rect 5022 -29573 5032 -29513
rect 5092 -29573 5352 -29513
rect 5412 -29573 5422 -29513
rect 5022 -29683 5422 -29573
rect 5480 -29513 5880 -29503
rect 5480 -29573 5490 -29513
rect 5550 -29573 5810 -29513
rect 5870 -29573 5880 -29513
rect 5480 -29683 5880 -29573
rect 5936 -29513 6336 -29503
rect 5936 -29573 5946 -29513
rect 6006 -29573 6266 -29513
rect 6326 -29573 6336 -29513
rect 5936 -29683 6336 -29573
rect 6392 -29513 6792 -29503
rect 6392 -29573 6402 -29513
rect 6462 -29573 6722 -29513
rect 6782 -29573 6792 -29513
rect 6392 -29683 6792 -29573
rect 6850 -29513 7250 -29503
rect 6850 -29573 6860 -29513
rect 6920 -29573 7180 -29513
rect 7240 -29573 7250 -29513
rect 6850 -29683 7250 -29573
rect 7306 -29513 7706 -29503
rect 7306 -29573 7316 -29513
rect 7376 -29573 7636 -29513
rect 7696 -29573 7706 -29513
rect 7306 -29683 7706 -29573
rect 7762 -29513 8162 -29503
rect 7762 -29573 7772 -29513
rect 7832 -29573 8092 -29513
rect 8152 -29573 8162 -29513
rect 7762 -29683 8162 -29573
rect 8236 -29513 8636 -29503
rect 8236 -29573 8246 -29513
rect 8306 -29573 8566 -29513
rect 8626 -29573 8636 -29513
rect 8236 -29683 8636 -29573
rect 8692 -29513 9092 -29503
rect 8692 -29573 8702 -29513
rect 8762 -29573 9022 -29513
rect 9082 -29573 9092 -29513
rect 8692 -29683 9092 -29573
rect 9150 -29513 9550 -29503
rect 9150 -29573 9160 -29513
rect 9220 -29573 9480 -29513
rect 9540 -29573 9550 -29513
rect 9150 -29683 9550 -29573
rect 9606 -29513 10006 -29503
rect 9606 -29573 9616 -29513
rect 9676 -29573 9936 -29513
rect 9996 -29573 10006 -29513
rect 9606 -29683 10006 -29573
rect 10062 -29513 10462 -29503
rect 10062 -29573 10072 -29513
rect 10132 -29573 10392 -29513
rect 10452 -29573 10462 -29513
rect 10062 -29683 10462 -29573
rect 10520 -29513 10920 -29503
rect 10520 -29573 10530 -29513
rect 10590 -29573 10850 -29513
rect 10910 -29573 10920 -29513
rect 10520 -29683 10920 -29573
rect 10976 -29513 11376 -29503
rect 10976 -29573 10986 -29513
rect 11046 -29573 11306 -29513
rect 11366 -29573 11376 -29513
rect 10976 -29683 11376 -29573
rect 11432 -29513 11832 -29503
rect 11432 -29573 11442 -29513
rect 11502 -29573 11762 -29513
rect 11822 -29573 11832 -29513
rect 11432 -29683 11832 -29573
rect 11890 -29513 12290 -29503
rect 11890 -29573 11900 -29513
rect 11960 -29573 12220 -29513
rect 12280 -29573 12290 -29513
rect 11890 -29683 12290 -29573
rect 12346 -29513 12746 -29503
rect 12346 -29573 12356 -29513
rect 12416 -29573 12676 -29513
rect 12736 -29573 12746 -29513
rect 12346 -29683 12746 -29573
rect 12802 -29513 13202 -29503
rect 12802 -29573 12812 -29513
rect 12872 -29573 13132 -29513
rect 13192 -29573 13202 -29513
rect 12802 -29683 13202 -29573
rect 13260 -29513 13660 -29503
rect 13260 -29573 13270 -29513
rect 13330 -29573 13590 -29513
rect 13650 -29573 13660 -29513
rect 13260 -29683 13660 -29573
rect 13716 -29513 14116 -29503
rect 13716 -29573 13726 -29513
rect 13786 -29573 14046 -29513
rect 14106 -29573 14116 -29513
rect 13716 -29683 14116 -29573
rect 14172 -29513 14572 -29503
rect 14172 -29573 14182 -29513
rect 14242 -29573 14502 -29513
rect 14562 -29573 14572 -29513
rect 14172 -29683 14572 -29573
rect 14630 -29513 15030 -29503
rect 14630 -29573 14640 -29513
rect 14700 -29573 14960 -29513
rect 15020 -29573 15030 -29513
rect 14630 -29683 15030 -29573
rect 15086 -29513 15486 -29503
rect 15086 -29573 15096 -29513
rect 15156 -29573 15416 -29513
rect 15476 -29573 15486 -29513
rect 15086 -29683 15486 -29573
rect 456 -29753 15486 -29683
rect 456 -29863 856 -29753
rect 456 -29923 466 -29863
rect 526 -29923 786 -29863
rect 846 -29923 856 -29863
rect 456 -29933 856 -29923
rect 912 -29863 1312 -29753
rect 912 -29923 922 -29863
rect 982 -29923 1242 -29863
rect 1302 -29923 1312 -29863
rect 912 -29933 1312 -29923
rect 1370 -29863 1770 -29753
rect 1370 -29923 1380 -29863
rect 1440 -29923 1700 -29863
rect 1760 -29923 1770 -29863
rect 1370 -29933 1770 -29923
rect 1826 -29863 2226 -29753
rect 1826 -29923 1836 -29863
rect 1896 -29923 2156 -29863
rect 2216 -29923 2226 -29863
rect 1826 -29933 2226 -29923
rect 2282 -29863 2682 -29753
rect 2282 -29923 2292 -29863
rect 2352 -29923 2612 -29863
rect 2672 -29923 2682 -29863
rect 2282 -29933 2682 -29923
rect 2740 -29863 3140 -29753
rect 2740 -29923 2750 -29863
rect 2810 -29923 3070 -29863
rect 3130 -29923 3140 -29863
rect 2740 -29933 3140 -29923
rect 3196 -29863 3596 -29753
rect 3196 -29923 3206 -29863
rect 3266 -29923 3526 -29863
rect 3586 -29923 3596 -29863
rect 3196 -29933 3596 -29923
rect 3652 -29863 4052 -29753
rect 3652 -29923 3662 -29863
rect 3722 -29923 3982 -29863
rect 4042 -29923 4052 -29863
rect 3652 -29933 4052 -29923
rect 4110 -29863 4510 -29753
rect 4110 -29923 4120 -29863
rect 4180 -29923 4440 -29863
rect 4500 -29923 4510 -29863
rect 4110 -29933 4510 -29923
rect 4566 -29863 4966 -29753
rect 4566 -29923 4576 -29863
rect 4636 -29923 4896 -29863
rect 4956 -29923 4966 -29863
rect 4566 -29933 4966 -29923
rect 5022 -29863 5422 -29753
rect 5022 -29923 5032 -29863
rect 5092 -29923 5352 -29863
rect 5412 -29923 5422 -29863
rect 5022 -29933 5422 -29923
rect 5480 -29863 5880 -29753
rect 5480 -29923 5490 -29863
rect 5550 -29923 5810 -29863
rect 5870 -29923 5880 -29863
rect 5480 -29933 5880 -29923
rect 5936 -29863 6336 -29753
rect 5936 -29923 5946 -29863
rect 6006 -29923 6266 -29863
rect 6326 -29923 6336 -29863
rect 5936 -29933 6336 -29923
rect 6392 -29863 6792 -29753
rect 6392 -29923 6402 -29863
rect 6462 -29923 6722 -29863
rect 6782 -29923 6792 -29863
rect 6392 -29933 6792 -29923
rect 6850 -29863 7250 -29753
rect 6850 -29923 6860 -29863
rect 6920 -29923 7180 -29863
rect 7240 -29923 7250 -29863
rect 6850 -29933 7250 -29923
rect 7306 -29863 7706 -29753
rect 7306 -29923 7316 -29863
rect 7376 -29923 7636 -29863
rect 7696 -29923 7706 -29863
rect 7306 -29933 7706 -29923
rect 7762 -29863 8162 -29753
rect 7762 -29923 7772 -29863
rect 7832 -29923 8092 -29863
rect 8152 -29923 8162 -29863
rect 7762 -29933 8162 -29923
rect 8236 -29863 8636 -29753
rect 8236 -29923 8246 -29863
rect 8306 -29923 8566 -29863
rect 8626 -29923 8636 -29863
rect 8236 -29933 8636 -29923
rect 8692 -29863 9092 -29753
rect 8692 -29923 8702 -29863
rect 8762 -29923 9022 -29863
rect 9082 -29923 9092 -29863
rect 8692 -29933 9092 -29923
rect 9150 -29863 9550 -29753
rect 9150 -29923 9160 -29863
rect 9220 -29923 9480 -29863
rect 9540 -29923 9550 -29863
rect 9150 -29933 9550 -29923
rect 9606 -29863 10006 -29753
rect 9606 -29923 9616 -29863
rect 9676 -29923 9936 -29863
rect 9996 -29923 10006 -29863
rect 9606 -29933 10006 -29923
rect 10062 -29863 10462 -29753
rect 10062 -29923 10072 -29863
rect 10132 -29923 10392 -29863
rect 10452 -29923 10462 -29863
rect 10062 -29933 10462 -29923
rect 10520 -29863 10920 -29753
rect 10520 -29923 10530 -29863
rect 10590 -29923 10850 -29863
rect 10910 -29923 10920 -29863
rect 10520 -29933 10920 -29923
rect 10976 -29863 11376 -29753
rect 10976 -29923 10986 -29863
rect 11046 -29923 11306 -29863
rect 11366 -29923 11376 -29863
rect 10976 -29933 11376 -29923
rect 11432 -29863 11832 -29753
rect 11432 -29923 11442 -29863
rect 11502 -29923 11762 -29863
rect 11822 -29923 11832 -29863
rect 11432 -29933 11832 -29923
rect 11890 -29863 12290 -29753
rect 11890 -29923 11900 -29863
rect 11960 -29923 12220 -29863
rect 12280 -29923 12290 -29863
rect 11890 -29933 12290 -29923
rect 12346 -29863 12746 -29753
rect 12346 -29923 12356 -29863
rect 12416 -29923 12676 -29863
rect 12736 -29923 12746 -29863
rect 12346 -29933 12746 -29923
rect 12802 -29863 13202 -29753
rect 12802 -29923 12812 -29863
rect 12872 -29923 13132 -29863
rect 13192 -29923 13202 -29863
rect 12802 -29933 13202 -29923
rect 13260 -29863 13660 -29753
rect 13260 -29923 13270 -29863
rect 13330 -29923 13590 -29863
rect 13650 -29923 13660 -29863
rect 13260 -29933 13660 -29923
rect 13716 -29863 14116 -29753
rect 13716 -29923 13726 -29863
rect 13786 -29923 14046 -29863
rect 14106 -29923 14116 -29863
rect 13716 -29933 14116 -29923
rect 14172 -29863 14572 -29753
rect 14172 -29923 14182 -29863
rect 14242 -29923 14502 -29863
rect 14562 -29923 14572 -29863
rect 14172 -29933 14572 -29923
rect 14630 -29863 15030 -29753
rect 14630 -29923 14640 -29863
rect 14700 -29923 14960 -29863
rect 15020 -29923 15030 -29863
rect 14630 -29933 15030 -29923
rect 15086 -29863 15486 -29753
rect 15086 -29923 15096 -29863
rect 15156 -29923 15416 -29863
rect 15476 -29923 15486 -29863
rect 15086 -29933 15486 -29923
rect 66 -30005 80 -29933
rect 456 -30005 526 -29933
rect 912 -30005 983 -29933
rect 1370 -30005 1441 -29933
rect 1826 -30005 1897 -29933
rect 2282 -30005 2353 -29933
rect 2740 -30005 2811 -29933
rect 3196 -30005 3267 -29933
rect 3652 -30005 3723 -29933
rect 4110 -30005 4181 -29933
rect 4566 -30005 4637 -29933
rect 5022 -30005 5093 -29933
rect 5480 -30005 5551 -29933
rect 5936 -30005 6007 -29933
rect 6392 -30005 6463 -29933
rect 6850 -30005 6921 -29933
rect 7306 -30005 7377 -29933
rect 7762 -30005 7833 -29933
rect 8236 -30005 8307 -29933
rect 8692 -30005 8763 -29933
rect 9150 -30005 9221 -29933
rect 9606 -30005 9677 -29933
rect 10062 -30005 10133 -29933
rect 10520 -30005 10591 -29933
rect 10976 -30005 11047 -29933
rect 11432 -30005 11503 -29933
rect 11890 -30005 11961 -29933
rect 12346 -30005 12417 -29933
rect 12802 -30005 12873 -29933
rect 13260 -30005 13331 -29933
rect 13716 -30005 13787 -29933
rect 14172 -30005 14243 -29933
rect 14630 -30005 14701 -29933
rect 66 -30015 400 -30005
rect 0 -30075 10 -30015
rect 70 -30075 330 -30015
rect 390 -30075 400 -30015
rect 0 -30365 14 -30075
rect 66 -30365 400 -30075
rect 0 -30425 10 -30365
rect 70 -30425 330 -30365
rect 390 -30425 400 -30365
rect 0 -30531 14 -30425
rect 66 -30435 400 -30425
rect 456 -30015 856 -30005
rect 456 -30075 466 -30015
rect 526 -30075 786 -30015
rect 846 -30075 856 -30015
rect 456 -30184 856 -30075
rect 912 -30015 1312 -30005
rect 912 -30075 922 -30015
rect 982 -30075 1242 -30015
rect 1302 -30075 1312 -30015
rect 912 -30184 1312 -30075
rect 1370 -30015 1770 -30005
rect 1370 -30075 1380 -30015
rect 1440 -30075 1700 -30015
rect 1760 -30075 1770 -30015
rect 1370 -30184 1770 -30075
rect 1826 -30015 2226 -30005
rect 1826 -30075 1836 -30015
rect 1896 -30075 2156 -30015
rect 2216 -30075 2226 -30015
rect 1826 -30184 2226 -30075
rect 2282 -30015 2682 -30005
rect 2282 -30075 2292 -30015
rect 2352 -30075 2612 -30015
rect 2672 -30075 2682 -30015
rect 2282 -30184 2682 -30075
rect 2740 -30015 3140 -30005
rect 2740 -30075 2750 -30015
rect 2810 -30075 3070 -30015
rect 3130 -30075 3140 -30015
rect 2740 -30184 3140 -30075
rect 3196 -30015 3596 -30005
rect 3196 -30075 3206 -30015
rect 3266 -30075 3526 -30015
rect 3586 -30075 3596 -30015
rect 3196 -30184 3596 -30075
rect 3652 -30015 4052 -30005
rect 3652 -30075 3662 -30015
rect 3722 -30075 3982 -30015
rect 4042 -30075 4052 -30015
rect 3652 -30184 4052 -30075
rect 4110 -30015 4510 -30005
rect 4110 -30075 4120 -30015
rect 4180 -30075 4440 -30015
rect 4500 -30075 4510 -30015
rect 4110 -30184 4510 -30075
rect 4566 -30015 4966 -30005
rect 4566 -30075 4576 -30015
rect 4636 -30075 4896 -30015
rect 4956 -30075 4966 -30015
rect 4566 -30184 4966 -30075
rect 5022 -30015 5422 -30005
rect 5022 -30075 5032 -30015
rect 5092 -30075 5352 -30015
rect 5412 -30075 5422 -30015
rect 5022 -30184 5422 -30075
rect 5480 -30015 5880 -30005
rect 5480 -30075 5490 -30015
rect 5550 -30075 5810 -30015
rect 5870 -30075 5880 -30015
rect 5480 -30184 5880 -30075
rect 5936 -30015 6336 -30005
rect 5936 -30075 5946 -30015
rect 6006 -30075 6266 -30015
rect 6326 -30075 6336 -30015
rect 5936 -30184 6336 -30075
rect 6392 -30015 6792 -30005
rect 6392 -30075 6402 -30015
rect 6462 -30075 6722 -30015
rect 6782 -30075 6792 -30015
rect 6392 -30184 6792 -30075
rect 6850 -30015 7250 -30005
rect 6850 -30075 6860 -30015
rect 6920 -30075 7180 -30015
rect 7240 -30075 7250 -30015
rect 6850 -30184 7250 -30075
rect 7306 -30015 7706 -30005
rect 7306 -30075 7316 -30015
rect 7376 -30075 7636 -30015
rect 7696 -30075 7706 -30015
rect 7306 -30184 7706 -30075
rect 7762 -30015 8162 -30005
rect 7762 -30075 7772 -30015
rect 7832 -30075 8092 -30015
rect 8152 -30075 8162 -30015
rect 7762 -30184 8162 -30075
rect 8236 -30015 8636 -30005
rect 8236 -30075 8246 -30015
rect 8306 -30075 8566 -30015
rect 8626 -30075 8636 -30015
rect 8236 -30184 8636 -30075
rect 8692 -30015 9092 -30005
rect 8692 -30075 8702 -30015
rect 8762 -30075 9022 -30015
rect 9082 -30075 9092 -30015
rect 8692 -30184 9092 -30075
rect 9150 -30015 9550 -30005
rect 9150 -30075 9160 -30015
rect 9220 -30075 9480 -30015
rect 9540 -30075 9550 -30015
rect 9150 -30184 9550 -30075
rect 9606 -30015 10006 -30005
rect 9606 -30075 9616 -30015
rect 9676 -30075 9936 -30015
rect 9996 -30075 10006 -30015
rect 9606 -30184 10006 -30075
rect 10062 -30015 10462 -30005
rect 10062 -30075 10072 -30015
rect 10132 -30075 10392 -30015
rect 10452 -30075 10462 -30015
rect 10062 -30184 10462 -30075
rect 10520 -30015 10920 -30005
rect 10520 -30075 10530 -30015
rect 10590 -30075 10850 -30015
rect 10910 -30075 10920 -30015
rect 10520 -30184 10920 -30075
rect 10976 -30015 11376 -30005
rect 10976 -30075 10986 -30015
rect 11046 -30075 11306 -30015
rect 11366 -30075 11376 -30015
rect 10976 -30184 11376 -30075
rect 11432 -30015 11832 -30005
rect 11432 -30075 11442 -30015
rect 11502 -30075 11762 -30015
rect 11822 -30075 11832 -30015
rect 11432 -30184 11832 -30075
rect 11890 -30015 12290 -30005
rect 11890 -30075 11900 -30015
rect 11960 -30075 12220 -30015
rect 12280 -30075 12290 -30015
rect 11890 -30184 12290 -30075
rect 12346 -30015 12746 -30005
rect 12346 -30075 12356 -30015
rect 12416 -30075 12676 -30015
rect 12736 -30075 12746 -30015
rect 12346 -30184 12746 -30075
rect 12802 -30015 13202 -30005
rect 12802 -30075 12812 -30015
rect 12872 -30075 13132 -30015
rect 13192 -30075 13202 -30015
rect 12802 -30184 13202 -30075
rect 13260 -30015 13660 -30005
rect 13260 -30075 13270 -30015
rect 13330 -30075 13590 -30015
rect 13650 -30075 13660 -30015
rect 13260 -30184 13660 -30075
rect 13716 -30015 14116 -30005
rect 13716 -30075 13726 -30015
rect 13786 -30075 14046 -30015
rect 14106 -30075 14116 -30015
rect 13716 -30184 14116 -30075
rect 14172 -30015 14572 -30005
rect 14172 -30075 14182 -30015
rect 14242 -30075 14502 -30015
rect 14562 -30075 14572 -30015
rect 14172 -30184 14572 -30075
rect 14630 -30015 15030 -30005
rect 14630 -30075 14640 -30015
rect 14700 -30075 14960 -30015
rect 15020 -30075 15030 -30015
rect 14630 -30184 15030 -30075
rect 15086 -30015 15486 -30005
rect 15086 -30075 15096 -30015
rect 15156 -30075 15416 -30015
rect 15476 -30075 15486 -30015
rect 15086 -30184 15486 -30075
rect 456 -30254 15486 -30184
rect 456 -30255 2682 -30254
rect 456 -30365 856 -30255
rect 456 -30425 466 -30365
rect 526 -30425 786 -30365
rect 846 -30425 856 -30365
rect 456 -30435 856 -30425
rect 912 -30365 1312 -30255
rect 912 -30425 922 -30365
rect 982 -30425 1242 -30365
rect 1302 -30425 1312 -30365
rect 912 -30435 1312 -30425
rect 1370 -30365 1770 -30255
rect 1370 -30425 1380 -30365
rect 1440 -30425 1700 -30365
rect 1760 -30425 1770 -30365
rect 1370 -30435 1770 -30425
rect 1826 -30365 2226 -30255
rect 1826 -30425 1836 -30365
rect 1896 -30425 2156 -30365
rect 2216 -30425 2226 -30365
rect 1826 -30435 2226 -30425
rect 2282 -30365 2682 -30255
rect 2282 -30425 2292 -30365
rect 2352 -30425 2612 -30365
rect 2672 -30425 2682 -30365
rect 2282 -30435 2682 -30425
rect 2740 -30255 10462 -30254
rect 2740 -30365 3140 -30255
rect 2740 -30425 2750 -30365
rect 2810 -30425 3070 -30365
rect 3130 -30425 3140 -30365
rect 2740 -30435 3140 -30425
rect 3196 -30365 3596 -30255
rect 3196 -30425 3206 -30365
rect 3266 -30425 3526 -30365
rect 3586 -30425 3596 -30365
rect 3196 -30435 3596 -30425
rect 3652 -30365 4052 -30255
rect 3652 -30425 3662 -30365
rect 3722 -30425 3982 -30365
rect 4042 -30425 4052 -30365
rect 3652 -30435 4052 -30425
rect 4110 -30365 4510 -30255
rect 4110 -30425 4120 -30365
rect 4180 -30425 4440 -30365
rect 4500 -30425 4510 -30365
rect 4110 -30435 4510 -30425
rect 4566 -30365 4966 -30255
rect 4566 -30425 4576 -30365
rect 4636 -30425 4896 -30365
rect 4956 -30425 4966 -30365
rect 4566 -30435 4966 -30425
rect 5022 -30365 5422 -30255
rect 5022 -30425 5032 -30365
rect 5092 -30425 5352 -30365
rect 5412 -30425 5422 -30365
rect 5022 -30435 5422 -30425
rect 5480 -30365 5880 -30255
rect 5480 -30425 5490 -30365
rect 5550 -30425 5810 -30365
rect 5870 -30425 5880 -30365
rect 5480 -30435 5880 -30425
rect 5936 -30365 6336 -30255
rect 5936 -30425 5946 -30365
rect 6006 -30425 6266 -30365
rect 6326 -30425 6336 -30365
rect 5936 -30435 6336 -30425
rect 6392 -30365 6792 -30255
rect 6392 -30425 6402 -30365
rect 6462 -30425 6722 -30365
rect 6782 -30425 6792 -30365
rect 6392 -30435 6792 -30425
rect 6850 -30365 7250 -30255
rect 6850 -30425 6860 -30365
rect 6920 -30425 7180 -30365
rect 7240 -30425 7250 -30365
rect 6850 -30435 7250 -30425
rect 7306 -30365 7706 -30255
rect 7306 -30425 7316 -30365
rect 7376 -30425 7636 -30365
rect 7696 -30425 7706 -30365
rect 7306 -30435 7706 -30425
rect 7762 -30365 8162 -30255
rect 7762 -30425 7772 -30365
rect 7832 -30425 8092 -30365
rect 8152 -30425 8162 -30365
rect 7762 -30435 8162 -30425
rect 8236 -30365 8636 -30255
rect 8236 -30425 8246 -30365
rect 8306 -30425 8566 -30365
rect 8626 -30425 8636 -30365
rect 8236 -30435 8636 -30425
rect 8692 -30365 9092 -30255
rect 8692 -30425 8702 -30365
rect 8762 -30425 9022 -30365
rect 9082 -30425 9092 -30365
rect 8692 -30435 9092 -30425
rect 9150 -30365 9550 -30255
rect 9150 -30425 9160 -30365
rect 9220 -30425 9480 -30365
rect 9540 -30425 9550 -30365
rect 9150 -30435 9550 -30425
rect 9606 -30365 10006 -30255
rect 9606 -30425 9616 -30365
rect 9676 -30425 9936 -30365
rect 9996 -30425 10006 -30365
rect 9606 -30435 10006 -30425
rect 10062 -30365 10462 -30255
rect 10062 -30425 10072 -30365
rect 10132 -30425 10392 -30365
rect 10452 -30425 10462 -30365
rect 10062 -30435 10462 -30425
rect 10520 -30255 15486 -30254
rect 10520 -30365 10920 -30255
rect 10520 -30425 10530 -30365
rect 10590 -30425 10850 -30365
rect 10910 -30425 10920 -30365
rect 10520 -30435 10920 -30425
rect 10976 -30365 11376 -30255
rect 10976 -30425 10986 -30365
rect 11046 -30425 11306 -30365
rect 11366 -30425 11376 -30365
rect 10976 -30435 11376 -30425
rect 11432 -30365 11832 -30255
rect 11432 -30425 11442 -30365
rect 11502 -30425 11762 -30365
rect 11822 -30425 11832 -30365
rect 11432 -30435 11832 -30425
rect 11890 -30365 12290 -30255
rect 11890 -30425 11900 -30365
rect 11960 -30425 12220 -30365
rect 12280 -30425 12290 -30365
rect 11890 -30435 12290 -30425
rect 12346 -30365 12746 -30255
rect 12346 -30425 12356 -30365
rect 12416 -30425 12676 -30365
rect 12736 -30425 12746 -30365
rect 12346 -30435 12746 -30425
rect 12802 -30365 13202 -30255
rect 12802 -30425 12812 -30365
rect 12872 -30425 13132 -30365
rect 13192 -30425 13202 -30365
rect 12802 -30435 13202 -30425
rect 13260 -30365 13660 -30255
rect 13260 -30425 13270 -30365
rect 13330 -30425 13590 -30365
rect 13650 -30425 13660 -30365
rect 13260 -30435 13660 -30425
rect 13716 -30365 14116 -30255
rect 13716 -30425 13726 -30365
rect 13786 -30425 14046 -30365
rect 14106 -30425 14116 -30365
rect 13716 -30435 14116 -30425
rect 14172 -30365 14572 -30255
rect 14172 -30425 14182 -30365
rect 14242 -30425 14502 -30365
rect 14562 -30425 14572 -30365
rect 14172 -30435 14572 -30425
rect 14630 -30365 15030 -30255
rect 14630 -30425 14640 -30365
rect 14700 -30425 14960 -30365
rect 15020 -30425 15030 -30365
rect 14630 -30435 15030 -30425
rect 15086 -30365 15486 -30255
rect 15086 -30425 15096 -30365
rect 15156 -30425 15416 -30365
rect 15476 -30425 15486 -30365
rect 15086 -30435 15486 -30425
rect 66 -30521 80 -30435
rect 456 -30521 526 -30435
rect 912 -30521 982 -30435
rect 1370 -30521 1440 -30435
rect 1826 -30521 1896 -30435
rect 2282 -30521 2352 -30435
rect 2740 -30521 2810 -30435
rect 3196 -30521 3266 -30435
rect 3652 -30521 3722 -30435
rect 4110 -30521 4180 -30435
rect 4566 -30521 4636 -30435
rect 5022 -30521 5092 -30435
rect 5480 -30521 5550 -30435
rect 5936 -30521 6006 -30435
rect 6392 -30521 6462 -30435
rect 6850 -30521 6920 -30435
rect 7306 -30521 7376 -30435
rect 7762 -30521 7832 -30435
rect 8236 -30521 8306 -30435
rect 8692 -30521 8762 -30435
rect 9150 -30521 9220 -30435
rect 9606 -30521 9676 -30435
rect 10062 -30521 10132 -30435
rect 10520 -30521 10590 -30435
rect 10976 -30521 11046 -30435
rect 11432 -30521 11502 -30435
rect 11890 -30521 11960 -30435
rect 12346 -30521 12416 -30435
rect 12802 -30521 12872 -30435
rect 13260 -30521 13330 -30435
rect 13716 -30521 13786 -30435
rect 14172 -30521 14242 -30435
rect 14630 -30521 14700 -30435
rect 66 -30531 400 -30521
rect 0 -30591 10 -30531
rect 70 -30591 330 -30531
rect 390 -30591 400 -30531
rect 0 -30881 14 -30591
rect 66 -30881 400 -30591
rect 0 -30941 10 -30881
rect 70 -30941 330 -30881
rect 390 -30941 400 -30881
rect 0 -31023 14 -30941
rect 66 -30951 400 -30941
rect 456 -30531 856 -30521
rect 456 -30591 466 -30531
rect 526 -30591 786 -30531
rect 846 -30591 856 -30531
rect 456 -30699 856 -30591
rect 912 -30531 1312 -30521
rect 912 -30591 922 -30531
rect 982 -30591 1242 -30531
rect 1302 -30591 1312 -30531
rect 912 -30699 1312 -30591
rect 1370 -30531 1770 -30521
rect 1370 -30591 1380 -30531
rect 1440 -30591 1700 -30531
rect 1760 -30591 1770 -30531
rect 1370 -30699 1770 -30591
rect 1826 -30531 2226 -30521
rect 1826 -30591 1836 -30531
rect 1896 -30591 2156 -30531
rect 2216 -30591 2226 -30531
rect 1826 -30699 2226 -30591
rect 2282 -30531 2682 -30521
rect 2282 -30591 2292 -30531
rect 2352 -30591 2612 -30531
rect 2672 -30591 2682 -30531
rect 2282 -30699 2682 -30591
rect 2740 -30531 3140 -30521
rect 2740 -30591 2750 -30531
rect 2810 -30591 3070 -30531
rect 3130 -30591 3140 -30531
rect 2740 -30699 3140 -30591
rect 3196 -30531 3596 -30521
rect 3196 -30591 3206 -30531
rect 3266 -30591 3526 -30531
rect 3586 -30591 3596 -30531
rect 3196 -30699 3596 -30591
rect 3652 -30531 4052 -30521
rect 3652 -30591 3662 -30531
rect 3722 -30591 3982 -30531
rect 4042 -30591 4052 -30531
rect 3652 -30699 4052 -30591
rect 4110 -30531 4510 -30521
rect 4110 -30591 4120 -30531
rect 4180 -30591 4440 -30531
rect 4500 -30591 4510 -30531
rect 4110 -30699 4510 -30591
rect 4566 -30531 4966 -30521
rect 4566 -30591 4576 -30531
rect 4636 -30591 4896 -30531
rect 4956 -30591 4966 -30531
rect 4566 -30699 4966 -30591
rect 5022 -30531 5422 -30521
rect 5022 -30591 5032 -30531
rect 5092 -30591 5352 -30531
rect 5412 -30591 5422 -30531
rect 5022 -30699 5422 -30591
rect 5480 -30531 5880 -30521
rect 5480 -30591 5490 -30531
rect 5550 -30591 5810 -30531
rect 5870 -30591 5880 -30531
rect 5480 -30699 5880 -30591
rect 5936 -30531 6336 -30521
rect 5936 -30591 5946 -30531
rect 6006 -30591 6266 -30531
rect 6326 -30591 6336 -30531
rect 5936 -30699 6336 -30591
rect 6392 -30531 6792 -30521
rect 6392 -30591 6402 -30531
rect 6462 -30591 6722 -30531
rect 6782 -30591 6792 -30531
rect 6392 -30699 6792 -30591
rect 6850 -30531 7250 -30521
rect 6850 -30591 6860 -30531
rect 6920 -30591 7180 -30531
rect 7240 -30591 7250 -30531
rect 6850 -30699 7250 -30591
rect 7306 -30531 7706 -30521
rect 7306 -30591 7316 -30531
rect 7376 -30591 7636 -30531
rect 7696 -30591 7706 -30531
rect 7306 -30699 7706 -30591
rect 7762 -30531 8162 -30521
rect 7762 -30591 7772 -30531
rect 7832 -30591 8092 -30531
rect 8152 -30591 8162 -30531
rect 7762 -30699 8162 -30591
rect 8236 -30531 8636 -30521
rect 8236 -30591 8246 -30531
rect 8306 -30591 8566 -30531
rect 8626 -30591 8636 -30531
rect 8236 -30699 8636 -30591
rect 8692 -30531 9092 -30521
rect 8692 -30591 8702 -30531
rect 8762 -30591 9022 -30531
rect 9082 -30591 9092 -30531
rect 8692 -30699 9092 -30591
rect 9150 -30531 9550 -30521
rect 9150 -30591 9160 -30531
rect 9220 -30591 9480 -30531
rect 9540 -30591 9550 -30531
rect 9150 -30699 9550 -30591
rect 9606 -30531 10006 -30521
rect 9606 -30591 9616 -30531
rect 9676 -30591 9936 -30531
rect 9996 -30591 10006 -30531
rect 9606 -30699 10006 -30591
rect 10062 -30531 10462 -30521
rect 10062 -30591 10072 -30531
rect 10132 -30591 10392 -30531
rect 10452 -30591 10462 -30531
rect 10062 -30699 10462 -30591
rect 10520 -30531 10920 -30521
rect 10520 -30591 10530 -30531
rect 10590 -30591 10850 -30531
rect 10910 -30591 10920 -30531
rect 10520 -30699 10920 -30591
rect 10976 -30531 11376 -30521
rect 10976 -30591 10986 -30531
rect 11046 -30591 11306 -30531
rect 11366 -30591 11376 -30531
rect 10976 -30699 11376 -30591
rect 11432 -30531 11832 -30521
rect 11432 -30591 11442 -30531
rect 11502 -30591 11762 -30531
rect 11822 -30591 11832 -30531
rect 11432 -30699 11832 -30591
rect 11890 -30531 12290 -30521
rect 11890 -30591 11900 -30531
rect 11960 -30591 12220 -30531
rect 12280 -30591 12290 -30531
rect 11890 -30699 12290 -30591
rect 12346 -30531 12746 -30521
rect 12346 -30591 12356 -30531
rect 12416 -30591 12676 -30531
rect 12736 -30591 12746 -30531
rect 12346 -30699 12746 -30591
rect 12802 -30531 13202 -30521
rect 12802 -30591 12812 -30531
rect 12872 -30591 13132 -30531
rect 13192 -30591 13202 -30531
rect 12802 -30699 13202 -30591
rect 13260 -30531 13660 -30521
rect 13260 -30591 13270 -30531
rect 13330 -30591 13590 -30531
rect 13650 -30591 13660 -30531
rect 13260 -30699 13660 -30591
rect 13716 -30531 14116 -30521
rect 13716 -30591 13726 -30531
rect 13786 -30591 14046 -30531
rect 14106 -30591 14116 -30531
rect 13716 -30699 14116 -30591
rect 14172 -30531 14572 -30521
rect 14172 -30591 14182 -30531
rect 14242 -30591 14502 -30531
rect 14562 -30591 14572 -30531
rect 14172 -30699 14572 -30591
rect 14630 -30531 15030 -30521
rect 14630 -30591 14640 -30531
rect 14700 -30591 14960 -30531
rect 15020 -30591 15030 -30531
rect 14630 -30699 15030 -30591
rect 15086 -30531 15486 -30521
rect 15086 -30591 15096 -30531
rect 15156 -30591 15416 -30531
rect 15476 -30591 15486 -30531
rect 15086 -30699 15486 -30591
rect 456 -30769 15486 -30699
rect 456 -30771 2682 -30769
rect 456 -30881 856 -30771
rect 456 -30941 466 -30881
rect 526 -30941 786 -30881
rect 846 -30941 856 -30881
rect 456 -30951 856 -30941
rect 912 -30881 1312 -30771
rect 912 -30941 922 -30881
rect 982 -30941 1242 -30881
rect 1302 -30941 1312 -30881
rect 912 -30951 1312 -30941
rect 1370 -30881 1770 -30771
rect 1370 -30941 1380 -30881
rect 1440 -30941 1700 -30881
rect 1760 -30941 1770 -30881
rect 1370 -30951 1770 -30941
rect 1826 -30881 2226 -30771
rect 1826 -30941 1836 -30881
rect 1896 -30941 2156 -30881
rect 2216 -30941 2226 -30881
rect 1826 -30951 2226 -30941
rect 2282 -30881 2682 -30771
rect 2282 -30941 2292 -30881
rect 2352 -30941 2612 -30881
rect 2672 -30941 2682 -30881
rect 2282 -30951 2682 -30941
rect 2740 -30771 10462 -30769
rect 2740 -30881 3140 -30771
rect 2740 -30941 2750 -30881
rect 2810 -30941 3070 -30881
rect 3130 -30941 3140 -30881
rect 2740 -30951 3140 -30941
rect 3196 -30881 3596 -30771
rect 3196 -30941 3206 -30881
rect 3266 -30941 3526 -30881
rect 3586 -30941 3596 -30881
rect 3196 -30951 3596 -30941
rect 3652 -30881 4052 -30771
rect 3652 -30941 3662 -30881
rect 3722 -30941 3982 -30881
rect 4042 -30941 4052 -30881
rect 3652 -30951 4052 -30941
rect 4110 -30881 4510 -30771
rect 4110 -30941 4120 -30881
rect 4180 -30941 4440 -30881
rect 4500 -30941 4510 -30881
rect 4110 -30951 4510 -30941
rect 4566 -30881 4966 -30771
rect 4566 -30941 4576 -30881
rect 4636 -30941 4896 -30881
rect 4956 -30941 4966 -30881
rect 4566 -30951 4966 -30941
rect 5022 -30881 5422 -30771
rect 5022 -30941 5032 -30881
rect 5092 -30941 5352 -30881
rect 5412 -30941 5422 -30881
rect 5022 -30951 5422 -30941
rect 5480 -30881 5880 -30771
rect 5480 -30941 5490 -30881
rect 5550 -30941 5810 -30881
rect 5870 -30941 5880 -30881
rect 5480 -30951 5880 -30941
rect 5936 -30881 6336 -30771
rect 5936 -30941 5946 -30881
rect 6006 -30941 6266 -30881
rect 6326 -30941 6336 -30881
rect 5936 -30951 6336 -30941
rect 6392 -30881 6792 -30771
rect 6392 -30941 6402 -30881
rect 6462 -30941 6722 -30881
rect 6782 -30941 6792 -30881
rect 6392 -30951 6792 -30941
rect 6850 -30881 7250 -30771
rect 6850 -30941 6860 -30881
rect 6920 -30941 7180 -30881
rect 7240 -30941 7250 -30881
rect 6850 -30951 7250 -30941
rect 7306 -30881 7706 -30771
rect 7306 -30941 7316 -30881
rect 7376 -30941 7636 -30881
rect 7696 -30941 7706 -30881
rect 7306 -30951 7706 -30941
rect 7762 -30881 8162 -30771
rect 7762 -30941 7772 -30881
rect 7832 -30941 8092 -30881
rect 8152 -30941 8162 -30881
rect 7762 -30951 8162 -30941
rect 8236 -30881 8636 -30771
rect 8236 -30941 8246 -30881
rect 8306 -30941 8566 -30881
rect 8626 -30941 8636 -30881
rect 8236 -30951 8636 -30941
rect 8692 -30881 9092 -30771
rect 8692 -30941 8702 -30881
rect 8762 -30941 9022 -30881
rect 9082 -30941 9092 -30881
rect 8692 -30951 9092 -30941
rect 9150 -30881 9550 -30771
rect 9150 -30941 9160 -30881
rect 9220 -30941 9480 -30881
rect 9540 -30941 9550 -30881
rect 9150 -30951 9550 -30941
rect 9606 -30881 10006 -30771
rect 9606 -30941 9616 -30881
rect 9676 -30941 9936 -30881
rect 9996 -30941 10006 -30881
rect 9606 -30951 10006 -30941
rect 10062 -30881 10462 -30771
rect 10062 -30941 10072 -30881
rect 10132 -30941 10392 -30881
rect 10452 -30941 10462 -30881
rect 10062 -30951 10462 -30941
rect 10520 -30771 15486 -30769
rect 10520 -30881 10920 -30771
rect 10520 -30941 10530 -30881
rect 10590 -30941 10850 -30881
rect 10910 -30941 10920 -30881
rect 10520 -30951 10920 -30941
rect 10976 -30881 11376 -30771
rect 10976 -30941 10986 -30881
rect 11046 -30941 11306 -30881
rect 11366 -30941 11376 -30881
rect 10976 -30951 11376 -30941
rect 11432 -30881 11832 -30771
rect 11432 -30941 11442 -30881
rect 11502 -30941 11762 -30881
rect 11822 -30941 11832 -30881
rect 11432 -30951 11832 -30941
rect 11890 -30881 12290 -30771
rect 11890 -30941 11900 -30881
rect 11960 -30941 12220 -30881
rect 12280 -30941 12290 -30881
rect 11890 -30951 12290 -30941
rect 12346 -30881 12746 -30771
rect 12346 -30941 12356 -30881
rect 12416 -30941 12676 -30881
rect 12736 -30941 12746 -30881
rect 12346 -30951 12746 -30941
rect 12802 -30881 13202 -30771
rect 12802 -30941 12812 -30881
rect 12872 -30941 13132 -30881
rect 13192 -30941 13202 -30881
rect 12802 -30951 13202 -30941
rect 13260 -30881 13660 -30771
rect 13260 -30941 13270 -30881
rect 13330 -30941 13590 -30881
rect 13650 -30941 13660 -30881
rect 13260 -30951 13660 -30941
rect 13716 -30881 14116 -30771
rect 13716 -30941 13726 -30881
rect 13786 -30941 14046 -30881
rect 14106 -30941 14116 -30881
rect 13716 -30951 14116 -30941
rect 14172 -30881 14572 -30771
rect 14172 -30941 14182 -30881
rect 14242 -30941 14502 -30881
rect 14562 -30941 14572 -30881
rect 14172 -30951 14572 -30941
rect 14630 -30881 15030 -30771
rect 14630 -30941 14640 -30881
rect 14700 -30941 14960 -30881
rect 15020 -30941 15030 -30881
rect 14630 -30951 15030 -30941
rect 15086 -30881 15486 -30771
rect 15086 -30941 15096 -30881
rect 15156 -30941 15416 -30881
rect 15476 -30941 15486 -30881
rect 15086 -30951 15486 -30941
rect 66 -31013 80 -30951
rect 456 -31013 527 -30951
rect 912 -31013 983 -30951
rect 1370 -31013 1441 -30951
rect 1826 -31013 1897 -30951
rect 2282 -31013 2353 -30951
rect 2740 -31013 2810 -30951
rect 3196 -31013 3266 -30951
rect 3652 -31013 3722 -30951
rect 4110 -31013 4180 -30951
rect 4566 -31013 4636 -30951
rect 5022 -31013 5092 -30951
rect 5480 -31013 5550 -30951
rect 5936 -31013 6006 -30951
rect 6392 -31013 6462 -30951
rect 6850 -31013 6920 -30951
rect 7306 -31013 7376 -30951
rect 7762 -31013 7832 -30951
rect 8236 -31013 8306 -30951
rect 8692 -31013 8762 -30951
rect 9150 -31013 9220 -30951
rect 9606 -31013 9676 -30951
rect 10062 -31013 10132 -30951
rect 10520 -31013 10590 -30951
rect 10976 -31013 11046 -30951
rect 11432 -31013 11502 -30951
rect 11890 -31013 11960 -30951
rect 12346 -31013 12416 -30951
rect 12802 -31013 12872 -30951
rect 13260 -31013 13330 -30951
rect 13716 -31013 13786 -30951
rect 14172 -31013 14242 -30951
rect 14630 -31013 14700 -30951
rect 66 -31023 400 -31013
rect 0 -31083 10 -31023
rect 70 -31083 330 -31023
rect 390 -31083 400 -31023
rect 0 -31373 14 -31083
rect 66 -31373 400 -31083
rect 0 -31433 10 -31373
rect 70 -31433 330 -31373
rect 390 -31433 400 -31373
rect 0 -31525 14 -31433
rect 66 -31443 400 -31433
rect 456 -31023 856 -31013
rect 456 -31083 466 -31023
rect 526 -31083 786 -31023
rect 846 -31083 856 -31023
rect 456 -31191 856 -31083
rect 912 -31023 1312 -31013
rect 912 -31083 922 -31023
rect 982 -31083 1242 -31023
rect 1302 -31083 1312 -31023
rect 912 -31191 1312 -31083
rect 1370 -31023 1770 -31013
rect 1370 -31083 1380 -31023
rect 1440 -31083 1700 -31023
rect 1760 -31083 1770 -31023
rect 1370 -31191 1770 -31083
rect 1826 -31023 2226 -31013
rect 1826 -31083 1836 -31023
rect 1896 -31083 2156 -31023
rect 2216 -31083 2226 -31023
rect 1826 -31191 2226 -31083
rect 2282 -31023 2682 -31013
rect 2282 -31083 2292 -31023
rect 2352 -31083 2612 -31023
rect 2672 -31083 2682 -31023
rect 2282 -31191 2682 -31083
rect 2740 -31023 3140 -31013
rect 2740 -31083 2750 -31023
rect 2810 -31083 3070 -31023
rect 3130 -31083 3140 -31023
rect 2740 -31191 3140 -31083
rect 3196 -31023 3596 -31013
rect 3196 -31083 3206 -31023
rect 3266 -31083 3526 -31023
rect 3586 -31083 3596 -31023
rect 3196 -31191 3596 -31083
rect 3652 -31023 4052 -31013
rect 3652 -31083 3662 -31023
rect 3722 -31083 3982 -31023
rect 4042 -31083 4052 -31023
rect 3652 -31191 4052 -31083
rect 4110 -31023 4510 -31013
rect 4110 -31083 4120 -31023
rect 4180 -31083 4440 -31023
rect 4500 -31083 4510 -31023
rect 4110 -31191 4510 -31083
rect 4566 -31023 4966 -31013
rect 4566 -31083 4576 -31023
rect 4636 -31083 4896 -31023
rect 4956 -31083 4966 -31023
rect 4566 -31191 4966 -31083
rect 5022 -31023 5422 -31013
rect 5022 -31083 5032 -31023
rect 5092 -31083 5352 -31023
rect 5412 -31083 5422 -31023
rect 5022 -31191 5422 -31083
rect 5480 -31023 5880 -31013
rect 5480 -31083 5490 -31023
rect 5550 -31083 5810 -31023
rect 5870 -31083 5880 -31023
rect 5480 -31191 5880 -31083
rect 5936 -31023 6336 -31013
rect 5936 -31083 5946 -31023
rect 6006 -31083 6266 -31023
rect 6326 -31083 6336 -31023
rect 5936 -31191 6336 -31083
rect 6392 -31023 6792 -31013
rect 6392 -31083 6402 -31023
rect 6462 -31083 6722 -31023
rect 6782 -31083 6792 -31023
rect 6392 -31191 6792 -31083
rect 6850 -31023 7250 -31013
rect 6850 -31083 6860 -31023
rect 6920 -31083 7180 -31023
rect 7240 -31083 7250 -31023
rect 6850 -31191 7250 -31083
rect 7306 -31023 7706 -31013
rect 7306 -31083 7316 -31023
rect 7376 -31083 7636 -31023
rect 7696 -31083 7706 -31023
rect 7306 -31191 7706 -31083
rect 7762 -31023 8162 -31013
rect 7762 -31083 7772 -31023
rect 7832 -31083 8092 -31023
rect 8152 -31083 8162 -31023
rect 7762 -31191 8162 -31083
rect 8236 -31023 8636 -31013
rect 8236 -31083 8246 -31023
rect 8306 -31083 8566 -31023
rect 8626 -31083 8636 -31023
rect 8236 -31191 8636 -31083
rect 8692 -31023 9092 -31013
rect 8692 -31083 8702 -31023
rect 8762 -31083 9022 -31023
rect 9082 -31083 9092 -31023
rect 8692 -31191 9092 -31083
rect 9150 -31023 9550 -31013
rect 9150 -31083 9160 -31023
rect 9220 -31083 9480 -31023
rect 9540 -31083 9550 -31023
rect 9150 -31191 9550 -31083
rect 9606 -31023 10006 -31013
rect 9606 -31083 9616 -31023
rect 9676 -31083 9936 -31023
rect 9996 -31083 10006 -31023
rect 9606 -31191 10006 -31083
rect 10062 -31023 10462 -31013
rect 10062 -31083 10072 -31023
rect 10132 -31083 10392 -31023
rect 10452 -31083 10462 -31023
rect 10062 -31191 10462 -31083
rect 10520 -31023 10920 -31013
rect 10520 -31083 10530 -31023
rect 10590 -31083 10850 -31023
rect 10910 -31083 10920 -31023
rect 10520 -31191 10920 -31083
rect 10976 -31023 11376 -31013
rect 10976 -31083 10986 -31023
rect 11046 -31083 11306 -31023
rect 11366 -31083 11376 -31023
rect 10976 -31191 11376 -31083
rect 11432 -31023 11832 -31013
rect 11432 -31083 11442 -31023
rect 11502 -31083 11762 -31023
rect 11822 -31083 11832 -31023
rect 11432 -31191 11832 -31083
rect 11890 -31023 12290 -31013
rect 11890 -31083 11900 -31023
rect 11960 -31083 12220 -31023
rect 12280 -31083 12290 -31023
rect 11890 -31191 12290 -31083
rect 12346 -31023 12746 -31013
rect 12346 -31083 12356 -31023
rect 12416 -31083 12676 -31023
rect 12736 -31083 12746 -31023
rect 12346 -31191 12746 -31083
rect 12802 -31023 13202 -31013
rect 12802 -31083 12812 -31023
rect 12872 -31083 13132 -31023
rect 13192 -31083 13202 -31023
rect 12802 -31191 13202 -31083
rect 13260 -31023 13660 -31013
rect 13260 -31083 13270 -31023
rect 13330 -31083 13590 -31023
rect 13650 -31083 13660 -31023
rect 13260 -31191 13660 -31083
rect 13716 -31023 14116 -31013
rect 13716 -31083 13726 -31023
rect 13786 -31083 14046 -31023
rect 14106 -31083 14116 -31023
rect 13716 -31191 14116 -31083
rect 14172 -31023 14572 -31013
rect 14172 -31083 14182 -31023
rect 14242 -31083 14502 -31023
rect 14562 -31083 14572 -31023
rect 14172 -31191 14572 -31083
rect 14630 -31023 15030 -31013
rect 14630 -31083 14640 -31023
rect 14700 -31083 14960 -31023
rect 15020 -31083 15030 -31023
rect 14630 -31191 15030 -31083
rect 15086 -31023 15486 -31013
rect 15086 -31083 15096 -31023
rect 15156 -31083 15416 -31023
rect 15476 -31083 15486 -31023
rect 15086 -31191 15486 -31083
rect 456 -31261 15486 -31191
rect 456 -31263 2682 -31261
rect 456 -31373 856 -31263
rect 456 -31433 466 -31373
rect 526 -31433 786 -31373
rect 846 -31433 856 -31373
rect 456 -31443 856 -31433
rect 912 -31373 1312 -31263
rect 912 -31433 922 -31373
rect 982 -31433 1242 -31373
rect 1302 -31433 1312 -31373
rect 912 -31443 1312 -31433
rect 1370 -31373 1770 -31263
rect 1370 -31433 1380 -31373
rect 1440 -31433 1700 -31373
rect 1760 -31433 1770 -31373
rect 1370 -31443 1770 -31433
rect 1826 -31373 2226 -31263
rect 1826 -31433 1836 -31373
rect 1896 -31433 2156 -31373
rect 2216 -31433 2226 -31373
rect 1826 -31443 2226 -31433
rect 2282 -31373 2682 -31263
rect 2282 -31433 2292 -31373
rect 2352 -31433 2612 -31373
rect 2672 -31433 2682 -31373
rect 2282 -31443 2682 -31433
rect 2740 -31263 10462 -31261
rect 2740 -31373 3140 -31263
rect 2740 -31433 2750 -31373
rect 2810 -31433 3070 -31373
rect 3130 -31433 3140 -31373
rect 2740 -31443 3140 -31433
rect 3196 -31373 3596 -31263
rect 3196 -31433 3206 -31373
rect 3266 -31433 3526 -31373
rect 3586 -31433 3596 -31373
rect 3196 -31443 3596 -31433
rect 3652 -31373 4052 -31263
rect 3652 -31433 3662 -31373
rect 3722 -31433 3982 -31373
rect 4042 -31433 4052 -31373
rect 3652 -31443 4052 -31433
rect 4110 -31373 4510 -31263
rect 4110 -31433 4120 -31373
rect 4180 -31433 4440 -31373
rect 4500 -31433 4510 -31373
rect 4110 -31443 4510 -31433
rect 4566 -31373 4966 -31263
rect 4566 -31433 4576 -31373
rect 4636 -31433 4896 -31373
rect 4956 -31433 4966 -31373
rect 4566 -31443 4966 -31433
rect 5022 -31373 5422 -31263
rect 5022 -31433 5032 -31373
rect 5092 -31433 5352 -31373
rect 5412 -31433 5422 -31373
rect 5022 -31443 5422 -31433
rect 5480 -31373 5880 -31263
rect 5480 -31433 5490 -31373
rect 5550 -31433 5810 -31373
rect 5870 -31433 5880 -31373
rect 5480 -31443 5880 -31433
rect 5936 -31373 6336 -31263
rect 5936 -31433 5946 -31373
rect 6006 -31433 6266 -31373
rect 6326 -31433 6336 -31373
rect 5936 -31443 6336 -31433
rect 6392 -31373 6792 -31263
rect 6392 -31433 6402 -31373
rect 6462 -31433 6722 -31373
rect 6782 -31433 6792 -31373
rect 6392 -31443 6792 -31433
rect 6850 -31373 7250 -31263
rect 6850 -31433 6860 -31373
rect 6920 -31433 7180 -31373
rect 7240 -31433 7250 -31373
rect 6850 -31443 7250 -31433
rect 7306 -31373 7706 -31263
rect 7306 -31433 7316 -31373
rect 7376 -31433 7636 -31373
rect 7696 -31433 7706 -31373
rect 7306 -31443 7706 -31433
rect 7762 -31373 8162 -31263
rect 7762 -31433 7772 -31373
rect 7832 -31433 8092 -31373
rect 8152 -31433 8162 -31373
rect 7762 -31443 8162 -31433
rect 8236 -31373 8636 -31263
rect 8236 -31433 8246 -31373
rect 8306 -31433 8566 -31373
rect 8626 -31433 8636 -31373
rect 8236 -31443 8636 -31433
rect 8692 -31373 9092 -31263
rect 8692 -31433 8702 -31373
rect 8762 -31433 9022 -31373
rect 9082 -31433 9092 -31373
rect 8692 -31443 9092 -31433
rect 9150 -31373 9550 -31263
rect 9150 -31433 9160 -31373
rect 9220 -31433 9480 -31373
rect 9540 -31433 9550 -31373
rect 9150 -31443 9550 -31433
rect 9606 -31373 10006 -31263
rect 9606 -31433 9616 -31373
rect 9676 -31433 9936 -31373
rect 9996 -31433 10006 -31373
rect 9606 -31443 10006 -31433
rect 10062 -31373 10462 -31263
rect 10062 -31433 10072 -31373
rect 10132 -31433 10392 -31373
rect 10452 -31433 10462 -31373
rect 10062 -31443 10462 -31433
rect 10520 -31263 15486 -31261
rect 10520 -31373 10920 -31263
rect 10520 -31433 10530 -31373
rect 10590 -31433 10850 -31373
rect 10910 -31433 10920 -31373
rect 10520 -31443 10920 -31433
rect 10976 -31373 11376 -31263
rect 10976 -31433 10986 -31373
rect 11046 -31433 11306 -31373
rect 11366 -31433 11376 -31373
rect 10976 -31443 11376 -31433
rect 11432 -31373 11832 -31263
rect 11432 -31433 11442 -31373
rect 11502 -31433 11762 -31373
rect 11822 -31433 11832 -31373
rect 11432 -31443 11832 -31433
rect 11890 -31373 12290 -31263
rect 11890 -31433 11900 -31373
rect 11960 -31433 12220 -31373
rect 12280 -31433 12290 -31373
rect 11890 -31443 12290 -31433
rect 12346 -31373 12746 -31263
rect 12346 -31433 12356 -31373
rect 12416 -31433 12676 -31373
rect 12736 -31433 12746 -31373
rect 12346 -31443 12746 -31433
rect 12802 -31373 13202 -31263
rect 12802 -31433 12812 -31373
rect 12872 -31433 13132 -31373
rect 13192 -31433 13202 -31373
rect 12802 -31443 13202 -31433
rect 13260 -31373 13660 -31263
rect 13260 -31433 13270 -31373
rect 13330 -31433 13590 -31373
rect 13650 -31433 13660 -31373
rect 13260 -31443 13660 -31433
rect 13716 -31373 14116 -31263
rect 13716 -31433 13726 -31373
rect 13786 -31433 14046 -31373
rect 14106 -31433 14116 -31373
rect 13716 -31443 14116 -31433
rect 14172 -31373 14572 -31263
rect 14172 -31433 14182 -31373
rect 14242 -31433 14502 -31373
rect 14562 -31433 14572 -31373
rect 14172 -31443 14572 -31433
rect 14630 -31373 15030 -31263
rect 14630 -31433 14640 -31373
rect 14700 -31433 14960 -31373
rect 15020 -31433 15030 -31373
rect 14630 -31443 15030 -31433
rect 15086 -31373 15486 -31263
rect 15086 -31433 15096 -31373
rect 15156 -31433 15416 -31373
rect 15476 -31433 15486 -31373
rect 15086 -31443 15486 -31433
rect 66 -31515 80 -31443
rect 456 -31515 526 -31443
rect 912 -31515 983 -31443
rect 1370 -31515 1441 -31443
rect 1826 -31515 1897 -31443
rect 2282 -31515 2353 -31443
rect 2740 -31515 2811 -31443
rect 3196 -31515 3267 -31443
rect 3652 -31515 3723 -31443
rect 4110 -31515 4181 -31443
rect 4566 -31515 4637 -31443
rect 5022 -31515 5093 -31443
rect 5480 -31515 5551 -31443
rect 5936 -31515 6007 -31443
rect 6392 -31515 6463 -31443
rect 6850 -31515 6921 -31443
rect 7306 -31515 7377 -31443
rect 7762 -31515 7833 -31443
rect 8236 -31515 8307 -31443
rect 8692 -31515 8763 -31443
rect 9150 -31515 9221 -31443
rect 9606 -31515 9677 -31443
rect 10062 -31515 10133 -31443
rect 10520 -31515 10591 -31443
rect 10976 -31515 11047 -31443
rect 11432 -31515 11503 -31443
rect 11890 -31515 11961 -31443
rect 12346 -31515 12417 -31443
rect 12802 -31515 12873 -31443
rect 13260 -31515 13331 -31443
rect 13716 -31515 13787 -31443
rect 14172 -31515 14243 -31443
rect 14630 -31515 14701 -31443
rect 66 -31525 400 -31515
rect 0 -31585 10 -31525
rect 70 -31585 330 -31525
rect 390 -31585 400 -31525
rect 0 -31875 14 -31585
rect 66 -31875 400 -31585
rect 0 -31935 10 -31875
rect 70 -31935 330 -31875
rect 390 -31935 400 -31875
rect 0 -32017 14 -31935
rect 66 -31945 400 -31935
rect 456 -31525 856 -31515
rect 456 -31585 466 -31525
rect 526 -31585 786 -31525
rect 846 -31585 856 -31525
rect 456 -31694 856 -31585
rect 912 -31525 1312 -31515
rect 912 -31585 922 -31525
rect 982 -31585 1242 -31525
rect 1302 -31585 1312 -31525
rect 912 -31694 1312 -31585
rect 1370 -31525 1770 -31515
rect 1370 -31585 1380 -31525
rect 1440 -31585 1700 -31525
rect 1760 -31585 1770 -31525
rect 1370 -31694 1770 -31585
rect 1826 -31525 2226 -31515
rect 1826 -31585 1836 -31525
rect 1896 -31585 2156 -31525
rect 2216 -31585 2226 -31525
rect 1826 -31694 2226 -31585
rect 2282 -31525 2682 -31515
rect 2282 -31585 2292 -31525
rect 2352 -31585 2612 -31525
rect 2672 -31585 2682 -31525
rect 2282 -31694 2682 -31585
rect 2740 -31525 3140 -31515
rect 2740 -31585 2750 -31525
rect 2810 -31585 3070 -31525
rect 3130 -31585 3140 -31525
rect 2740 -31694 3140 -31585
rect 3196 -31525 3596 -31515
rect 3196 -31585 3206 -31525
rect 3266 -31585 3526 -31525
rect 3586 -31585 3596 -31525
rect 3196 -31694 3596 -31585
rect 3652 -31525 4052 -31515
rect 3652 -31585 3662 -31525
rect 3722 -31585 3982 -31525
rect 4042 -31585 4052 -31525
rect 3652 -31694 4052 -31585
rect 4110 -31525 4510 -31515
rect 4110 -31585 4120 -31525
rect 4180 -31585 4440 -31525
rect 4500 -31585 4510 -31525
rect 4110 -31694 4510 -31585
rect 4566 -31525 4966 -31515
rect 4566 -31585 4576 -31525
rect 4636 -31585 4896 -31525
rect 4956 -31585 4966 -31525
rect 4566 -31694 4966 -31585
rect 5022 -31525 5422 -31515
rect 5022 -31585 5032 -31525
rect 5092 -31585 5352 -31525
rect 5412 -31585 5422 -31525
rect 5022 -31694 5422 -31585
rect 5480 -31525 5880 -31515
rect 5480 -31585 5490 -31525
rect 5550 -31585 5810 -31525
rect 5870 -31585 5880 -31525
rect 5480 -31694 5880 -31585
rect 5936 -31525 6336 -31515
rect 5936 -31585 5946 -31525
rect 6006 -31585 6266 -31525
rect 6326 -31585 6336 -31525
rect 5936 -31694 6336 -31585
rect 6392 -31525 6792 -31515
rect 6392 -31585 6402 -31525
rect 6462 -31585 6722 -31525
rect 6782 -31585 6792 -31525
rect 6392 -31694 6792 -31585
rect 6850 -31525 7250 -31515
rect 6850 -31585 6860 -31525
rect 6920 -31585 7180 -31525
rect 7240 -31585 7250 -31525
rect 6850 -31694 7250 -31585
rect 7306 -31525 7706 -31515
rect 7306 -31585 7316 -31525
rect 7376 -31585 7636 -31525
rect 7696 -31585 7706 -31525
rect 7306 -31694 7706 -31585
rect 7762 -31525 8162 -31515
rect 7762 -31585 7772 -31525
rect 7832 -31585 8092 -31525
rect 8152 -31585 8162 -31525
rect 7762 -31694 8162 -31585
rect 8236 -31525 8636 -31515
rect 8236 -31585 8246 -31525
rect 8306 -31585 8566 -31525
rect 8626 -31585 8636 -31525
rect 8236 -31694 8636 -31585
rect 8692 -31525 9092 -31515
rect 8692 -31585 8702 -31525
rect 8762 -31585 9022 -31525
rect 9082 -31585 9092 -31525
rect 8692 -31694 9092 -31585
rect 9150 -31525 9550 -31515
rect 9150 -31585 9160 -31525
rect 9220 -31585 9480 -31525
rect 9540 -31585 9550 -31525
rect 9150 -31694 9550 -31585
rect 9606 -31525 10006 -31515
rect 9606 -31585 9616 -31525
rect 9676 -31585 9936 -31525
rect 9996 -31585 10006 -31525
rect 9606 -31694 10006 -31585
rect 10062 -31525 10462 -31515
rect 10062 -31585 10072 -31525
rect 10132 -31585 10392 -31525
rect 10452 -31585 10462 -31525
rect 10062 -31694 10462 -31585
rect 10520 -31525 10920 -31515
rect 10520 -31585 10530 -31525
rect 10590 -31585 10850 -31525
rect 10910 -31585 10920 -31525
rect 10520 -31694 10920 -31585
rect 10976 -31525 11376 -31515
rect 10976 -31585 10986 -31525
rect 11046 -31585 11306 -31525
rect 11366 -31585 11376 -31525
rect 10976 -31694 11376 -31585
rect 11432 -31525 11832 -31515
rect 11432 -31585 11442 -31525
rect 11502 -31585 11762 -31525
rect 11822 -31585 11832 -31525
rect 11432 -31694 11832 -31585
rect 11890 -31525 12290 -31515
rect 11890 -31585 11900 -31525
rect 11960 -31585 12220 -31525
rect 12280 -31585 12290 -31525
rect 11890 -31694 12290 -31585
rect 12346 -31525 12746 -31515
rect 12346 -31585 12356 -31525
rect 12416 -31585 12676 -31525
rect 12736 -31585 12746 -31525
rect 12346 -31694 12746 -31585
rect 12802 -31525 13202 -31515
rect 12802 -31585 12812 -31525
rect 12872 -31585 13132 -31525
rect 13192 -31585 13202 -31525
rect 12802 -31694 13202 -31585
rect 13260 -31525 13660 -31515
rect 13260 -31585 13270 -31525
rect 13330 -31585 13590 -31525
rect 13650 -31585 13660 -31525
rect 13260 -31694 13660 -31585
rect 13716 -31525 14116 -31515
rect 13716 -31585 13726 -31525
rect 13786 -31585 14046 -31525
rect 14106 -31585 14116 -31525
rect 13716 -31694 14116 -31585
rect 14172 -31525 14572 -31515
rect 14172 -31585 14182 -31525
rect 14242 -31585 14502 -31525
rect 14562 -31585 14572 -31525
rect 14172 -31694 14572 -31585
rect 14630 -31525 15030 -31515
rect 14630 -31585 14640 -31525
rect 14700 -31585 14960 -31525
rect 15020 -31585 15030 -31525
rect 14630 -31694 15030 -31585
rect 15086 -31525 15486 -31515
rect 15086 -31585 15096 -31525
rect 15156 -31585 15416 -31525
rect 15476 -31585 15486 -31525
rect 15086 -31694 15486 -31585
rect 456 -31764 15486 -31694
rect 456 -31765 2682 -31764
rect 456 -31875 856 -31765
rect 456 -31935 466 -31875
rect 526 -31935 786 -31875
rect 846 -31935 856 -31875
rect 456 -31945 856 -31935
rect 912 -31875 1312 -31765
rect 912 -31935 922 -31875
rect 982 -31935 1242 -31875
rect 1302 -31935 1312 -31875
rect 912 -31945 1312 -31935
rect 1370 -31875 1770 -31765
rect 1370 -31935 1380 -31875
rect 1440 -31935 1700 -31875
rect 1760 -31935 1770 -31875
rect 1370 -31945 1770 -31935
rect 1826 -31875 2226 -31765
rect 1826 -31935 1836 -31875
rect 1896 -31935 2156 -31875
rect 2216 -31935 2226 -31875
rect 1826 -31945 2226 -31935
rect 2282 -31875 2682 -31765
rect 2282 -31935 2292 -31875
rect 2352 -31935 2612 -31875
rect 2672 -31935 2682 -31875
rect 2282 -31945 2682 -31935
rect 2740 -31765 10462 -31764
rect 2740 -31875 3140 -31765
rect 2740 -31935 2750 -31875
rect 2810 -31935 3070 -31875
rect 3130 -31935 3140 -31875
rect 2740 -31945 3140 -31935
rect 3196 -31875 3596 -31765
rect 3196 -31935 3206 -31875
rect 3266 -31935 3526 -31875
rect 3586 -31935 3596 -31875
rect 3196 -31945 3596 -31935
rect 3652 -31875 4052 -31765
rect 3652 -31935 3662 -31875
rect 3722 -31935 3982 -31875
rect 4042 -31935 4052 -31875
rect 3652 -31945 4052 -31935
rect 4110 -31875 4510 -31765
rect 4110 -31935 4120 -31875
rect 4180 -31935 4440 -31875
rect 4500 -31935 4510 -31875
rect 4110 -31945 4510 -31935
rect 4566 -31875 4966 -31765
rect 4566 -31935 4576 -31875
rect 4636 -31935 4896 -31875
rect 4956 -31935 4966 -31875
rect 4566 -31945 4966 -31935
rect 5022 -31875 5422 -31765
rect 5022 -31935 5032 -31875
rect 5092 -31935 5352 -31875
rect 5412 -31935 5422 -31875
rect 5022 -31945 5422 -31935
rect 5480 -31875 5880 -31765
rect 5480 -31935 5490 -31875
rect 5550 -31935 5810 -31875
rect 5870 -31935 5880 -31875
rect 5480 -31945 5880 -31935
rect 5936 -31875 6336 -31765
rect 5936 -31935 5946 -31875
rect 6006 -31935 6266 -31875
rect 6326 -31935 6336 -31875
rect 5936 -31945 6336 -31935
rect 6392 -31875 6792 -31765
rect 6392 -31935 6402 -31875
rect 6462 -31935 6722 -31875
rect 6782 -31935 6792 -31875
rect 6392 -31945 6792 -31935
rect 6850 -31875 7250 -31765
rect 6850 -31935 6860 -31875
rect 6920 -31935 7180 -31875
rect 7240 -31935 7250 -31875
rect 6850 -31945 7250 -31935
rect 7306 -31875 7706 -31765
rect 7306 -31935 7316 -31875
rect 7376 -31935 7636 -31875
rect 7696 -31935 7706 -31875
rect 7306 -31945 7706 -31935
rect 7762 -31875 8162 -31765
rect 7762 -31935 7772 -31875
rect 7832 -31935 8092 -31875
rect 8152 -31935 8162 -31875
rect 7762 -31945 8162 -31935
rect 8236 -31875 8636 -31765
rect 8236 -31935 8246 -31875
rect 8306 -31935 8566 -31875
rect 8626 -31935 8636 -31875
rect 8236 -31945 8636 -31935
rect 8692 -31875 9092 -31765
rect 8692 -31935 8702 -31875
rect 8762 -31935 9022 -31875
rect 9082 -31935 9092 -31875
rect 8692 -31945 9092 -31935
rect 9150 -31875 9550 -31765
rect 9150 -31935 9160 -31875
rect 9220 -31935 9480 -31875
rect 9540 -31935 9550 -31875
rect 9150 -31945 9550 -31935
rect 9606 -31875 10006 -31765
rect 9606 -31935 9616 -31875
rect 9676 -31935 9936 -31875
rect 9996 -31935 10006 -31875
rect 9606 -31945 10006 -31935
rect 10062 -31875 10462 -31765
rect 10062 -31935 10072 -31875
rect 10132 -31935 10392 -31875
rect 10452 -31935 10462 -31875
rect 10062 -31945 10462 -31935
rect 10520 -31765 15486 -31764
rect 10520 -31875 10920 -31765
rect 10520 -31935 10530 -31875
rect 10590 -31935 10850 -31875
rect 10910 -31935 10920 -31875
rect 10520 -31945 10920 -31935
rect 10976 -31875 11376 -31765
rect 10976 -31935 10986 -31875
rect 11046 -31935 11306 -31875
rect 11366 -31935 11376 -31875
rect 10976 -31945 11376 -31935
rect 11432 -31875 11832 -31765
rect 11432 -31935 11442 -31875
rect 11502 -31935 11762 -31875
rect 11822 -31935 11832 -31875
rect 11432 -31945 11832 -31935
rect 11890 -31875 12290 -31765
rect 11890 -31935 11900 -31875
rect 11960 -31935 12220 -31875
rect 12280 -31935 12290 -31875
rect 11890 -31945 12290 -31935
rect 12346 -31875 12746 -31765
rect 12346 -31935 12356 -31875
rect 12416 -31935 12676 -31875
rect 12736 -31935 12746 -31875
rect 12346 -31945 12746 -31935
rect 12802 -31875 13202 -31765
rect 12802 -31935 12812 -31875
rect 12872 -31935 13132 -31875
rect 13192 -31935 13202 -31875
rect 12802 -31945 13202 -31935
rect 13260 -31875 13660 -31765
rect 13260 -31935 13270 -31875
rect 13330 -31935 13590 -31875
rect 13650 -31935 13660 -31875
rect 13260 -31945 13660 -31935
rect 13716 -31875 14116 -31765
rect 13716 -31935 13726 -31875
rect 13786 -31935 14046 -31875
rect 14106 -31935 14116 -31875
rect 13716 -31945 14116 -31935
rect 14172 -31875 14572 -31765
rect 14172 -31935 14182 -31875
rect 14242 -31935 14502 -31875
rect 14562 -31935 14572 -31875
rect 14172 -31945 14572 -31935
rect 14630 -31875 15030 -31765
rect 14630 -31935 14640 -31875
rect 14700 -31935 14960 -31875
rect 15020 -31935 15030 -31875
rect 14630 -31945 15030 -31935
rect 15086 -31875 15486 -31765
rect 15086 -31935 15096 -31875
rect 15156 -31935 15416 -31875
rect 15476 -31935 15486 -31875
rect 15086 -31945 15486 -31935
rect 66 -32007 80 -31945
rect 66 -32017 400 -32007
rect 0 -32077 10 -32017
rect 70 -32077 330 -32017
rect 390 -32077 400 -32017
rect 0 -32110 14 -32077
rect 66 -32110 400 -32077
rect 0 -32180 400 -32110
rect 456 -32017 856 -32007
rect 456 -32077 466 -32017
rect 526 -32077 786 -32017
rect 846 -32077 856 -32017
rect 456 -32180 856 -32077
rect 912 -32017 1312 -32007
rect 912 -32077 922 -32017
rect 982 -32077 1242 -32017
rect 1302 -32077 1312 -32017
rect 912 -32180 1312 -32077
rect 1370 -32017 1770 -32007
rect 1370 -32077 1380 -32017
rect 1440 -32077 1700 -32017
rect 1760 -32077 1770 -32017
rect 1370 -32180 1770 -32077
rect 1826 -32017 2226 -32007
rect 1826 -32077 1836 -32017
rect 1896 -32077 2156 -32017
rect 2216 -32077 2226 -32017
rect 1826 -32180 2226 -32077
rect 2282 -32017 2682 -32007
rect 2282 -32077 2292 -32017
rect 2352 -32077 2612 -32017
rect 2672 -32077 2682 -32017
rect 2282 -32180 2682 -32077
rect 2740 -32017 3140 -32007
rect 2740 -32077 2750 -32017
rect 2810 -32077 3070 -32017
rect 3130 -32077 3140 -32017
rect 2740 -32180 3140 -32077
rect 3196 -32017 3596 -32007
rect 3196 -32077 3206 -32017
rect 3266 -32077 3526 -32017
rect 3586 -32077 3596 -32017
rect 3196 -32180 3596 -32077
rect 3652 -32017 4052 -32007
rect 3652 -32077 3662 -32017
rect 3722 -32077 3982 -32017
rect 4042 -32077 4052 -32017
rect 3652 -32180 4052 -32077
rect 4110 -32017 4510 -32007
rect 4110 -32077 4120 -32017
rect 4180 -32077 4440 -32017
rect 4500 -32077 4510 -32017
rect 4110 -32180 4510 -32077
rect 4566 -32017 4966 -32007
rect 4566 -32077 4576 -32017
rect 4636 -32077 4896 -32017
rect 4956 -32077 4966 -32017
rect 4566 -32180 4966 -32077
rect 5022 -32017 5422 -32007
rect 5022 -32077 5032 -32017
rect 5092 -32077 5352 -32017
rect 5412 -32077 5422 -32017
rect 5022 -32180 5422 -32077
rect 5480 -32017 5880 -32007
rect 5480 -32077 5490 -32017
rect 5550 -32077 5810 -32017
rect 5870 -32077 5880 -32017
rect 5480 -32180 5880 -32077
rect 5936 -32017 6336 -32007
rect 5936 -32077 5946 -32017
rect 6006 -32077 6266 -32017
rect 6326 -32077 6336 -32017
rect 5936 -32180 6336 -32077
rect 6392 -32017 6792 -32007
rect 6392 -32077 6402 -32017
rect 6462 -32077 6722 -32017
rect 6782 -32077 6792 -32017
rect 6392 -32180 6792 -32077
rect 6850 -32017 7250 -32007
rect 6850 -32077 6860 -32017
rect 6920 -32077 7180 -32017
rect 7240 -32077 7250 -32017
rect 6850 -32180 7250 -32077
rect 7306 -32017 7706 -32007
rect 7306 -32077 7316 -32017
rect 7376 -32077 7636 -32017
rect 7696 -32077 7706 -32017
rect 7306 -32180 7706 -32077
rect 7762 -32017 8162 -32007
rect 7762 -32077 7772 -32017
rect 7832 -32077 8092 -32017
rect 8152 -32077 8162 -32017
rect 7762 -32180 8162 -32077
rect 8236 -32017 8636 -32007
rect 8236 -32077 8246 -32017
rect 8306 -32077 8566 -32017
rect 8626 -32077 8636 -32017
rect 8236 -32180 8636 -32077
rect 8692 -32017 9092 -32007
rect 8692 -32077 8702 -32017
rect 8762 -32077 9022 -32017
rect 9082 -32077 9092 -32017
rect 8692 -32180 9092 -32077
rect 9150 -32017 9550 -32007
rect 9150 -32077 9160 -32017
rect 9220 -32077 9480 -32017
rect 9540 -32077 9550 -32017
rect 9150 -32180 9550 -32077
rect 9606 -32017 10006 -32007
rect 9606 -32077 9616 -32017
rect 9676 -32077 9936 -32017
rect 9996 -32077 10006 -32017
rect 9606 -32180 10006 -32077
rect 10062 -32017 10462 -32007
rect 10062 -32077 10072 -32017
rect 10132 -32077 10392 -32017
rect 10452 -32077 10462 -32017
rect 10062 -32180 10462 -32077
rect 10520 -32017 10920 -32007
rect 10520 -32077 10530 -32017
rect 10590 -32077 10850 -32017
rect 10910 -32077 10920 -32017
rect 10520 -32180 10920 -32077
rect 10976 -32017 11376 -32007
rect 10976 -32077 10986 -32017
rect 11046 -32077 11306 -32017
rect 11366 -32077 11376 -32017
rect 10976 -32180 11376 -32077
rect 11432 -32017 11832 -32007
rect 11432 -32077 11442 -32017
rect 11502 -32077 11762 -32017
rect 11822 -32077 11832 -32017
rect 11432 -32180 11832 -32077
rect 11890 -32017 12290 -32007
rect 11890 -32077 11900 -32017
rect 11960 -32077 12220 -32017
rect 12280 -32077 12290 -32017
rect 11890 -32180 12290 -32077
rect 12346 -32017 12746 -32007
rect 12346 -32077 12356 -32017
rect 12416 -32077 12676 -32017
rect 12736 -32077 12746 -32017
rect 12346 -32180 12746 -32077
rect 12802 -32017 13202 -32007
rect 12802 -32077 12812 -32017
rect 12872 -32077 13132 -32017
rect 13192 -32077 13202 -32017
rect 12802 -32180 13202 -32077
rect 13260 -32017 13660 -32007
rect 13260 -32077 13270 -32017
rect 13330 -32077 13590 -32017
rect 13650 -32077 13660 -32017
rect 13260 -32180 13660 -32077
rect 13716 -32017 14116 -32007
rect 13716 -32077 13726 -32017
rect 13786 -32077 14046 -32017
rect 14106 -32077 14116 -32017
rect 13716 -32180 14116 -32077
rect 14172 -32017 14572 -32007
rect 14172 -32077 14182 -32017
rect 14242 -32077 14502 -32017
rect 14562 -32077 14572 -32017
rect 14172 -32180 14572 -32077
rect 14630 -32017 15030 -32007
rect 14630 -32077 14640 -32017
rect 14700 -32077 14960 -32017
rect 15020 -32077 15030 -32017
rect 14630 -32180 15030 -32077
rect 15086 -32017 15486 -32007
rect 15086 -32077 15096 -32017
rect 15156 -32077 15416 -32017
rect 15476 -32077 15486 -32017
rect 15086 -32180 15486 -32077
rect 0 -32193 15486 -32180
rect 0 -32257 150 -32193
rect 15300 -32257 15486 -32193
rect 0 -32270 15486 -32257
rect 0 -32367 400 -32270
rect 0 -32427 10 -32367
rect 70 -32427 330 -32367
rect 390 -32427 400 -32367
rect 0 -32437 400 -32427
rect 456 -32367 856 -32270
rect 456 -32427 466 -32367
rect 526 -32427 786 -32367
rect 846 -32427 856 -32367
rect 456 -32437 856 -32427
rect 912 -32367 1312 -32270
rect 912 -32427 922 -32367
rect 982 -32427 1242 -32367
rect 1302 -32427 1312 -32367
rect 912 -32437 1312 -32427
rect 1370 -32367 1770 -32270
rect 1370 -32427 1380 -32367
rect 1440 -32427 1700 -32367
rect 1760 -32427 1770 -32367
rect 1370 -32437 1770 -32427
rect 1826 -32367 2226 -32270
rect 1826 -32427 1836 -32367
rect 1896 -32427 2156 -32367
rect 2216 -32427 2226 -32367
rect 1826 -32437 2226 -32427
rect 2282 -32367 2682 -32270
rect 2282 -32427 2292 -32367
rect 2352 -32427 2612 -32367
rect 2672 -32427 2682 -32367
rect 2282 -32437 2682 -32427
rect 2740 -32367 3140 -32270
rect 2740 -32427 2750 -32367
rect 2810 -32427 3070 -32367
rect 3130 -32427 3140 -32367
rect 2740 -32437 3140 -32427
rect 3196 -32367 3596 -32270
rect 3196 -32427 3206 -32367
rect 3266 -32427 3526 -32367
rect 3586 -32427 3596 -32367
rect 3196 -32437 3596 -32427
rect 3652 -32367 4052 -32270
rect 3652 -32427 3662 -32367
rect 3722 -32427 3982 -32367
rect 4042 -32427 4052 -32367
rect 3652 -32437 4052 -32427
rect 4110 -32367 4510 -32270
rect 4110 -32427 4120 -32367
rect 4180 -32427 4440 -32367
rect 4500 -32427 4510 -32367
rect 4110 -32437 4510 -32427
rect 4566 -32367 4966 -32270
rect 4566 -32427 4576 -32367
rect 4636 -32427 4896 -32367
rect 4956 -32427 4966 -32367
rect 4566 -32437 4966 -32427
rect 5022 -32367 5422 -32270
rect 5022 -32427 5032 -32367
rect 5092 -32427 5352 -32367
rect 5412 -32427 5422 -32367
rect 5022 -32437 5422 -32427
rect 5480 -32367 5880 -32270
rect 5480 -32427 5490 -32367
rect 5550 -32427 5810 -32367
rect 5870 -32427 5880 -32367
rect 5480 -32437 5880 -32427
rect 5936 -32367 6336 -32270
rect 5936 -32427 5946 -32367
rect 6006 -32427 6266 -32367
rect 6326 -32427 6336 -32367
rect 5936 -32437 6336 -32427
rect 6392 -32367 6792 -32270
rect 6392 -32427 6402 -32367
rect 6462 -32427 6722 -32367
rect 6782 -32427 6792 -32367
rect 6392 -32437 6792 -32427
rect 6850 -32367 7250 -32270
rect 6850 -32427 6860 -32367
rect 6920 -32427 7180 -32367
rect 7240 -32427 7250 -32367
rect 6850 -32437 7250 -32427
rect 7306 -32367 7706 -32270
rect 7306 -32427 7316 -32367
rect 7376 -32427 7636 -32367
rect 7696 -32427 7706 -32367
rect 7306 -32437 7706 -32427
rect 7762 -32367 8162 -32270
rect 7762 -32427 7772 -32367
rect 7832 -32427 8092 -32367
rect 8152 -32427 8162 -32367
rect 7762 -32437 8162 -32427
rect 8236 -32367 8636 -32270
rect 8236 -32427 8246 -32367
rect 8306 -32427 8566 -32367
rect 8626 -32427 8636 -32367
rect 8236 -32437 8636 -32427
rect 8692 -32367 9092 -32270
rect 8692 -32427 8702 -32367
rect 8762 -32427 9022 -32367
rect 9082 -32427 9092 -32367
rect 8692 -32437 9092 -32427
rect 9150 -32367 9550 -32270
rect 9150 -32427 9160 -32367
rect 9220 -32427 9480 -32367
rect 9540 -32427 9550 -32367
rect 9150 -32437 9550 -32427
rect 9606 -32367 10006 -32270
rect 9606 -32427 9616 -32367
rect 9676 -32427 9936 -32367
rect 9996 -32427 10006 -32367
rect 9606 -32437 10006 -32427
rect 10062 -32367 10462 -32270
rect 10062 -32427 10072 -32367
rect 10132 -32427 10392 -32367
rect 10452 -32427 10462 -32367
rect 10062 -32437 10462 -32427
rect 10520 -32367 10920 -32270
rect 10520 -32427 10530 -32367
rect 10590 -32427 10850 -32367
rect 10910 -32427 10920 -32367
rect 10520 -32437 10920 -32427
rect 10976 -32367 11376 -32270
rect 10976 -32427 10986 -32367
rect 11046 -32427 11306 -32367
rect 11366 -32427 11376 -32367
rect 10976 -32437 11376 -32427
rect 11432 -32367 11832 -32270
rect 11432 -32427 11442 -32367
rect 11502 -32427 11762 -32367
rect 11822 -32427 11832 -32367
rect 11432 -32437 11832 -32427
rect 11890 -32367 12290 -32270
rect 11890 -32427 11900 -32367
rect 11960 -32427 12220 -32367
rect 12280 -32427 12290 -32367
rect 11890 -32437 12290 -32427
rect 12346 -32367 12746 -32270
rect 12346 -32427 12356 -32367
rect 12416 -32427 12676 -32367
rect 12736 -32427 12746 -32367
rect 12346 -32437 12746 -32427
rect 12802 -32367 13202 -32270
rect 12802 -32427 12812 -32367
rect 12872 -32427 13132 -32367
rect 13192 -32427 13202 -32367
rect 12802 -32437 13202 -32427
rect 13260 -32367 13660 -32270
rect 13260 -32427 13270 -32367
rect 13330 -32427 13590 -32367
rect 13650 -32427 13660 -32367
rect 13260 -32437 13660 -32427
rect 13716 -32367 14116 -32270
rect 13716 -32427 13726 -32367
rect 13786 -32427 14046 -32367
rect 14106 -32427 14116 -32367
rect 13716 -32437 14116 -32427
rect 14172 -32367 14572 -32270
rect 14172 -32427 14182 -32367
rect 14242 -32427 14502 -32367
rect 14562 -32427 14572 -32367
rect 14172 -32437 14572 -32427
rect 14630 -32367 15030 -32270
rect 14630 -32427 14640 -32367
rect 14700 -32427 14960 -32367
rect 15020 -32427 15030 -32367
rect 14630 -32437 15030 -32427
rect 15086 -32367 15486 -32270
rect 15086 -32427 15096 -32367
rect 15156 -32427 15416 -32367
rect 15476 -32427 15486 -32367
rect 15086 -32437 15486 -32427
<< via2 >>
rect 89 590 150 651
rect 250 590 311 651
rect 15127 609 15201 611
rect 15127 551 15128 609
rect 15128 551 15201 609
rect 15358 609 15432 611
rect 15358 551 15359 609
rect 15359 551 15432 609
rect 1380 380 1440 440
rect 1700 380 1760 440
rect 1836 380 1896 440
rect 2156 380 2216 440
rect 2292 380 2352 440
rect 2612 380 2672 440
rect 2750 380 2810 440
rect 3070 380 3130 440
rect 3206 380 3266 440
rect 3526 380 3586 440
rect 3662 380 3722 440
rect 3982 380 4042 440
rect 4120 380 4180 440
rect 4440 380 4500 440
rect 4576 380 4636 440
rect 4896 380 4956 440
rect 5032 380 5092 440
rect 5352 380 5412 440
rect 5490 380 5550 440
rect 5810 380 5870 440
rect 5946 380 6006 440
rect 6266 380 6326 440
rect 6402 380 6462 440
rect 6722 380 6782 440
rect 6860 380 6920 440
rect 7180 380 7240 440
rect 7316 380 7376 440
rect 7636 380 7696 440
rect 7772 380 7832 440
rect 8092 380 8152 440
rect 8246 380 8306 440
rect 8566 380 8626 440
rect 8702 380 8762 440
rect 9022 380 9082 440
rect 9160 380 9220 440
rect 9480 380 9540 440
rect 9616 380 9676 440
rect 9936 380 9996 440
rect 10072 380 10132 440
rect 10392 380 10452 440
rect 10530 380 10590 440
rect 10850 380 10910 440
rect 10986 380 11046 440
rect 11306 380 11366 440
rect 11442 380 11502 440
rect 11762 380 11822 440
rect 11900 380 11960 440
rect 12220 380 12280 440
rect 12356 380 12416 440
rect 12676 380 12736 440
rect 12812 380 12872 440
rect 13132 380 13192 440
rect 13270 380 13330 440
rect 13590 380 13650 440
rect 13726 380 13786 440
rect 14046 380 14106 440
rect 14182 380 14242 440
rect 14502 380 14562 440
rect 14640 380 14700 440
rect 14960 380 15020 440
rect 15096 380 15156 440
rect 15416 380 15476 440
rect 1380 30 1440 90
rect 1700 30 1760 90
rect 1836 30 1896 90
rect 2156 30 2216 90
rect 2292 30 2352 90
rect 2612 30 2672 90
rect 2750 30 2810 90
rect 3070 30 3130 90
rect 3206 30 3266 90
rect 3526 30 3586 90
rect 3662 30 3722 90
rect 3982 30 4042 90
rect 4120 30 4180 90
rect 4440 30 4500 90
rect 4576 30 4636 90
rect 4896 30 4956 90
rect 5032 30 5092 90
rect 5352 30 5412 90
rect 5490 30 5550 90
rect 5810 30 5870 90
rect 5946 30 6006 90
rect 6266 30 6326 90
rect 6402 30 6462 90
rect 6722 30 6782 90
rect 6860 30 6920 90
rect 7180 30 7240 90
rect 7316 30 7376 90
rect 7636 30 7696 90
rect 7772 30 7832 90
rect 8092 30 8152 90
rect 8246 30 8306 90
rect 8566 30 8626 90
rect 8702 30 8762 90
rect 9022 30 9082 90
rect 9160 30 9220 90
rect 9480 30 9540 90
rect 9616 30 9676 90
rect 9936 30 9996 90
rect 10072 30 10132 90
rect 10392 30 10452 90
rect 10530 30 10590 90
rect 10850 30 10910 90
rect 10986 30 11046 90
rect 11306 30 11366 90
rect 11442 30 11502 90
rect 11762 30 11822 90
rect 11900 30 11960 90
rect 12220 30 12280 90
rect 12356 30 12416 90
rect 12676 30 12736 90
rect 12812 30 12872 90
rect 13132 30 13192 90
rect 13270 30 13330 90
rect 13590 30 13650 90
rect 13726 30 13786 90
rect 14046 30 14106 90
rect 14182 30 14242 90
rect 14502 30 14562 90
rect 14640 30 14700 90
rect 14960 30 15020 90
rect 15096 30 15156 90
rect 15416 30 15476 90
rect 10 -112 14 -52
rect 14 -112 66 -52
rect 66 -112 70 -52
rect 330 -112 390 -52
rect 10 -462 14 -402
rect 14 -462 66 -402
rect 66 -462 70 -402
rect 330 -462 390 -402
rect 466 -112 526 -52
rect 786 -112 846 -52
rect 922 -112 982 -52
rect 1242 -112 1302 -52
rect 1380 -112 1440 -52
rect 1700 -112 1760 -52
rect 1836 -112 1896 -52
rect 2156 -112 2216 -52
rect 2292 -112 2352 -52
rect 2612 -112 2672 -52
rect 2750 -112 2810 -52
rect 3070 -112 3130 -52
rect 3206 -112 3266 -52
rect 3526 -112 3586 -52
rect 3662 -112 3722 -52
rect 3982 -112 4042 -52
rect 4120 -112 4180 -52
rect 4440 -112 4500 -52
rect 4576 -112 4636 -52
rect 4896 -112 4956 -52
rect 5032 -112 5092 -52
rect 5352 -112 5412 -52
rect 5490 -112 5550 -52
rect 5810 -112 5870 -52
rect 5946 -112 6006 -52
rect 6266 -112 6326 -52
rect 6402 -112 6462 -52
rect 6722 -112 6782 -52
rect 6860 -112 6920 -52
rect 7180 -112 7240 -52
rect 7316 -112 7376 -52
rect 7636 -112 7696 -52
rect 7772 -112 7832 -52
rect 8092 -112 8152 -52
rect 8246 -112 8306 -52
rect 8566 -112 8626 -52
rect 8702 -112 8762 -52
rect 9022 -112 9082 -52
rect 9160 -112 9220 -52
rect 9480 -112 9540 -52
rect 9616 -112 9676 -52
rect 9936 -112 9996 -52
rect 10072 -112 10132 -52
rect 10392 -112 10452 -52
rect 10530 -112 10590 -52
rect 10850 -112 10910 -52
rect 10986 -112 11046 -52
rect 11306 -112 11366 -52
rect 11442 -112 11502 -52
rect 11762 -112 11822 -52
rect 11900 -112 11960 -52
rect 12220 -112 12280 -52
rect 12356 -112 12416 -52
rect 12676 -112 12736 -52
rect 12812 -112 12872 -52
rect 13132 -112 13192 -52
rect 13270 -112 13330 -52
rect 13590 -112 13650 -52
rect 13726 -112 13786 -52
rect 14046 -112 14106 -52
rect 14182 -112 14242 -52
rect 14502 -112 14562 -52
rect 14640 -112 14700 -52
rect 14960 -112 15020 -52
rect 15096 -112 15156 -52
rect 15416 -112 15476 -52
rect 466 -462 526 -402
rect 786 -462 846 -402
rect 922 -462 982 -402
rect 1242 -462 1302 -402
rect 1380 -462 1440 -402
rect 1700 -462 1760 -402
rect 1836 -462 1896 -402
rect 2156 -462 2216 -402
rect 2292 -462 2352 -402
rect 2612 -462 2672 -402
rect 2750 -462 2810 -402
rect 3070 -462 3130 -402
rect 3206 -462 3266 -402
rect 3526 -462 3586 -402
rect 3662 -462 3722 -402
rect 3982 -462 4042 -402
rect 4120 -462 4180 -402
rect 4440 -462 4500 -402
rect 4576 -462 4636 -402
rect 4896 -462 4956 -402
rect 5032 -462 5092 -402
rect 5352 -462 5412 -402
rect 5490 -462 5550 -402
rect 5810 -462 5870 -402
rect 5946 -462 6006 -402
rect 6266 -462 6326 -402
rect 6402 -462 6462 -402
rect 6722 -462 6782 -402
rect 6860 -462 6920 -402
rect 7180 -462 7240 -402
rect 7316 -462 7376 -402
rect 7636 -462 7696 -402
rect 7772 -462 7832 -402
rect 8092 -462 8152 -402
rect 8246 -462 8306 -402
rect 8566 -462 8626 -402
rect 8702 -462 8762 -402
rect 9022 -462 9082 -402
rect 9160 -462 9220 -402
rect 9480 -462 9540 -402
rect 9616 -462 9676 -402
rect 9936 -462 9996 -402
rect 10072 -462 10132 -402
rect 10392 -462 10452 -402
rect 10530 -462 10590 -402
rect 10850 -462 10910 -402
rect 10986 -462 11046 -402
rect 11306 -462 11366 -402
rect 11442 -462 11502 -402
rect 11762 -462 11822 -402
rect 11900 -462 11960 -402
rect 12220 -462 12280 -402
rect 12356 -462 12416 -402
rect 12676 -462 12736 -402
rect 12812 -462 12872 -402
rect 13132 -462 13192 -402
rect 13270 -462 13330 -402
rect 13590 -462 13650 -402
rect 13726 -462 13786 -402
rect 14046 -462 14106 -402
rect 14182 -462 14242 -402
rect 14502 -462 14562 -402
rect 14640 -462 14700 -402
rect 14960 -462 15020 -402
rect 15096 -462 15156 -402
rect 15416 -462 15476 -402
rect 10 -614 14 -554
rect 14 -614 66 -554
rect 66 -614 70 -554
rect 330 -614 390 -554
rect 10 -964 14 -904
rect 14 -964 66 -904
rect 66 -964 70 -904
rect 330 -964 390 -904
rect 466 -614 526 -554
rect 786 -614 846 -554
rect 922 -614 982 -554
rect 1242 -614 1302 -554
rect 1380 -614 1440 -554
rect 1700 -614 1760 -554
rect 1836 -614 1896 -554
rect 2156 -614 2216 -554
rect 2292 -614 2352 -554
rect 2612 -614 2672 -554
rect 2750 -614 2810 -554
rect 3070 -614 3130 -554
rect 3206 -614 3266 -554
rect 3526 -614 3586 -554
rect 3662 -614 3722 -554
rect 3982 -614 4042 -554
rect 4120 -614 4180 -554
rect 4440 -614 4500 -554
rect 4576 -614 4636 -554
rect 4896 -614 4956 -554
rect 5032 -614 5092 -554
rect 5352 -614 5412 -554
rect 5490 -614 5550 -554
rect 5810 -614 5870 -554
rect 5946 -614 6006 -554
rect 6266 -614 6326 -554
rect 6402 -614 6462 -554
rect 6722 -614 6782 -554
rect 6860 -614 6920 -554
rect 7180 -614 7240 -554
rect 7316 -614 7376 -554
rect 7636 -614 7696 -554
rect 7772 -614 7832 -554
rect 8092 -614 8152 -554
rect 8246 -614 8306 -554
rect 8566 -614 8626 -554
rect 8702 -614 8762 -554
rect 9022 -614 9082 -554
rect 9160 -614 9220 -554
rect 9480 -614 9540 -554
rect 9616 -614 9676 -554
rect 9936 -614 9996 -554
rect 10072 -614 10132 -554
rect 10392 -614 10452 -554
rect 10530 -614 10590 -554
rect 10850 -614 10910 -554
rect 10986 -614 11046 -554
rect 11306 -614 11366 -554
rect 11442 -614 11502 -554
rect 11762 -614 11822 -554
rect 11900 -614 11960 -554
rect 12220 -614 12280 -554
rect 12356 -614 12416 -554
rect 12676 -614 12736 -554
rect 12812 -614 12872 -554
rect 13132 -614 13192 -554
rect 13270 -614 13330 -554
rect 13590 -614 13650 -554
rect 13726 -614 13786 -554
rect 14046 -614 14106 -554
rect 14182 -614 14242 -554
rect 14502 -614 14562 -554
rect 14640 -614 14700 -554
rect 14960 -614 15020 -554
rect 15096 -614 15156 -554
rect 15416 -614 15476 -554
rect 466 -964 526 -904
rect 786 -964 846 -904
rect 922 -964 982 -904
rect 1242 -964 1302 -904
rect 1380 -964 1440 -904
rect 1700 -964 1760 -904
rect 1836 -964 1896 -904
rect 2156 -964 2216 -904
rect 2292 -964 2352 -904
rect 2612 -964 2672 -904
rect 2750 -964 2810 -904
rect 3070 -964 3130 -904
rect 3206 -964 3266 -904
rect 3526 -964 3586 -904
rect 3662 -964 3722 -904
rect 3982 -964 4042 -904
rect 4120 -964 4180 -904
rect 4440 -964 4500 -904
rect 4576 -964 4636 -904
rect 4896 -964 4956 -904
rect 5032 -964 5092 -904
rect 5352 -964 5412 -904
rect 5490 -964 5550 -904
rect 5810 -964 5870 -904
rect 5946 -964 6006 -904
rect 6266 -964 6326 -904
rect 6402 -964 6462 -904
rect 6722 -964 6782 -904
rect 6860 -964 6920 -904
rect 7180 -964 7240 -904
rect 7316 -964 7376 -904
rect 7636 -964 7696 -904
rect 7772 -964 7832 -904
rect 8092 -964 8152 -904
rect 8246 -964 8306 -904
rect 8566 -964 8626 -904
rect 8702 -964 8762 -904
rect 9022 -964 9082 -904
rect 9160 -964 9220 -904
rect 9480 -964 9540 -904
rect 9616 -964 9676 -904
rect 9936 -964 9996 -904
rect 10072 -964 10132 -904
rect 10392 -964 10452 -904
rect 10530 -964 10590 -904
rect 10850 -964 10910 -904
rect 10986 -964 11046 -904
rect 11306 -964 11366 -904
rect 11442 -964 11502 -904
rect 11762 -964 11822 -904
rect 11900 -964 11960 -904
rect 12220 -964 12280 -904
rect 12356 -964 12416 -904
rect 12676 -964 12736 -904
rect 12812 -964 12872 -904
rect 13132 -964 13192 -904
rect 13270 -964 13330 -904
rect 13590 -964 13650 -904
rect 13726 -964 13786 -904
rect 14046 -964 14106 -904
rect 14182 -964 14242 -904
rect 14502 -964 14562 -904
rect 14640 -964 14700 -904
rect 14960 -964 15020 -904
rect 15096 -964 15156 -904
rect 15416 -964 15476 -904
rect 10 -1106 14 -1046
rect 14 -1106 66 -1046
rect 66 -1106 70 -1046
rect 330 -1106 390 -1046
rect 10 -1456 14 -1396
rect 14 -1456 66 -1396
rect 66 -1456 70 -1396
rect 330 -1456 390 -1396
rect 466 -1106 526 -1046
rect 786 -1106 846 -1046
rect 922 -1106 982 -1046
rect 1242 -1106 1302 -1046
rect 1380 -1106 1440 -1046
rect 1700 -1106 1760 -1046
rect 1836 -1106 1896 -1046
rect 2156 -1106 2216 -1046
rect 2292 -1106 2352 -1046
rect 2612 -1106 2672 -1046
rect 2750 -1106 2810 -1046
rect 3070 -1106 3130 -1046
rect 3206 -1106 3266 -1046
rect 3526 -1106 3586 -1046
rect 3662 -1106 3722 -1046
rect 3982 -1106 4042 -1046
rect 4120 -1106 4180 -1046
rect 4440 -1106 4500 -1046
rect 4576 -1106 4636 -1046
rect 4896 -1106 4956 -1046
rect 5032 -1106 5092 -1046
rect 5352 -1106 5412 -1046
rect 5490 -1106 5550 -1046
rect 5810 -1106 5870 -1046
rect 5946 -1106 6006 -1046
rect 6266 -1106 6326 -1046
rect 6402 -1106 6462 -1046
rect 6722 -1106 6782 -1046
rect 6860 -1106 6920 -1046
rect 7180 -1106 7240 -1046
rect 7316 -1106 7376 -1046
rect 7636 -1106 7696 -1046
rect 7772 -1106 7832 -1046
rect 8092 -1106 8152 -1046
rect 8246 -1106 8306 -1046
rect 8566 -1106 8626 -1046
rect 8702 -1106 8762 -1046
rect 9022 -1106 9082 -1046
rect 9160 -1106 9220 -1046
rect 9480 -1106 9540 -1046
rect 9616 -1106 9676 -1046
rect 9936 -1106 9996 -1046
rect 10072 -1106 10132 -1046
rect 10392 -1106 10452 -1046
rect 10530 -1106 10590 -1046
rect 10850 -1106 10910 -1046
rect 10986 -1106 11046 -1046
rect 11306 -1106 11366 -1046
rect 11442 -1106 11502 -1046
rect 11762 -1106 11822 -1046
rect 11900 -1106 11960 -1046
rect 12220 -1106 12280 -1046
rect 12356 -1106 12416 -1046
rect 12676 -1106 12736 -1046
rect 12812 -1106 12872 -1046
rect 13132 -1106 13192 -1046
rect 13270 -1106 13330 -1046
rect 13590 -1106 13650 -1046
rect 13726 -1106 13786 -1046
rect 14046 -1106 14106 -1046
rect 14182 -1106 14242 -1046
rect 14502 -1106 14562 -1046
rect 14640 -1106 14700 -1046
rect 14960 -1106 15020 -1046
rect 15096 -1106 15156 -1046
rect 15416 -1106 15476 -1046
rect 466 -1456 526 -1396
rect 786 -1456 846 -1396
rect 922 -1456 982 -1396
rect 1242 -1456 1302 -1396
rect 1380 -1456 1440 -1396
rect 1700 -1456 1760 -1396
rect 1836 -1456 1896 -1396
rect 2156 -1456 2216 -1396
rect 2292 -1456 2352 -1396
rect 2612 -1456 2672 -1396
rect 2750 -1456 2810 -1396
rect 3070 -1456 3130 -1396
rect 3206 -1456 3266 -1396
rect 3526 -1456 3586 -1396
rect 3662 -1456 3722 -1396
rect 3982 -1456 4042 -1396
rect 4120 -1456 4180 -1396
rect 4440 -1456 4500 -1396
rect 4576 -1456 4636 -1396
rect 4896 -1456 4956 -1396
rect 5032 -1456 5092 -1396
rect 5352 -1456 5412 -1396
rect 5490 -1456 5550 -1396
rect 5810 -1456 5870 -1396
rect 5946 -1456 6006 -1396
rect 6266 -1456 6326 -1396
rect 6402 -1456 6462 -1396
rect 6722 -1456 6782 -1396
rect 6860 -1456 6920 -1396
rect 7180 -1456 7240 -1396
rect 7316 -1456 7376 -1396
rect 7636 -1456 7696 -1396
rect 7772 -1456 7832 -1396
rect 8092 -1456 8152 -1396
rect 8246 -1456 8306 -1396
rect 8566 -1456 8626 -1396
rect 8702 -1456 8762 -1396
rect 9022 -1456 9082 -1396
rect 9160 -1456 9220 -1396
rect 9480 -1456 9540 -1396
rect 9616 -1456 9676 -1396
rect 9936 -1456 9996 -1396
rect 10072 -1456 10132 -1396
rect 10392 -1456 10452 -1396
rect 10530 -1456 10590 -1396
rect 10850 -1456 10910 -1396
rect 10986 -1456 11046 -1396
rect 11306 -1456 11366 -1396
rect 11442 -1456 11502 -1396
rect 11762 -1456 11822 -1396
rect 11900 -1456 11960 -1396
rect 12220 -1456 12280 -1396
rect 12356 -1456 12416 -1396
rect 12676 -1456 12736 -1396
rect 12812 -1456 12872 -1396
rect 13132 -1456 13192 -1396
rect 13270 -1456 13330 -1396
rect 13590 -1456 13650 -1396
rect 13726 -1456 13786 -1396
rect 14046 -1456 14106 -1396
rect 14182 -1456 14242 -1396
rect 14502 -1456 14562 -1396
rect 14640 -1456 14700 -1396
rect 14960 -1456 15020 -1396
rect 15096 -1456 15156 -1396
rect 15416 -1456 15476 -1396
rect 10 -1622 14 -1562
rect 14 -1622 66 -1562
rect 66 -1622 70 -1562
rect 330 -1622 390 -1562
rect 10 -1972 14 -1912
rect 14 -1972 66 -1912
rect 66 -1972 70 -1912
rect 330 -1972 390 -1912
rect 466 -1622 526 -1562
rect 786 -1622 846 -1562
rect 922 -1622 982 -1562
rect 1242 -1622 1302 -1562
rect 1380 -1622 1440 -1562
rect 1700 -1622 1760 -1562
rect 1836 -1622 1896 -1562
rect 2156 -1622 2216 -1562
rect 2292 -1622 2352 -1562
rect 2612 -1622 2672 -1562
rect 2750 -1622 2810 -1562
rect 3070 -1622 3130 -1562
rect 3206 -1622 3266 -1562
rect 3526 -1622 3586 -1562
rect 3662 -1622 3722 -1562
rect 3982 -1622 4042 -1562
rect 4120 -1622 4180 -1562
rect 4440 -1622 4500 -1562
rect 4576 -1622 4636 -1562
rect 4896 -1622 4956 -1562
rect 5032 -1622 5092 -1562
rect 5352 -1622 5412 -1562
rect 5490 -1622 5550 -1562
rect 5810 -1622 5870 -1562
rect 5946 -1622 6006 -1562
rect 6266 -1622 6326 -1562
rect 6402 -1622 6462 -1562
rect 6722 -1622 6782 -1562
rect 6860 -1622 6920 -1562
rect 7180 -1622 7240 -1562
rect 7316 -1622 7376 -1562
rect 7636 -1622 7696 -1562
rect 7772 -1622 7832 -1562
rect 8092 -1622 8152 -1562
rect 8246 -1622 8306 -1562
rect 8566 -1622 8626 -1562
rect 8702 -1622 8762 -1562
rect 9022 -1622 9082 -1562
rect 9160 -1622 9220 -1562
rect 9480 -1622 9540 -1562
rect 9616 -1622 9676 -1562
rect 9936 -1622 9996 -1562
rect 10072 -1622 10132 -1562
rect 10392 -1622 10452 -1562
rect 10530 -1622 10590 -1562
rect 10850 -1622 10910 -1562
rect 10986 -1622 11046 -1562
rect 11306 -1622 11366 -1562
rect 11442 -1622 11502 -1562
rect 11762 -1622 11822 -1562
rect 11900 -1622 11960 -1562
rect 12220 -1622 12280 -1562
rect 12356 -1622 12416 -1562
rect 12676 -1622 12736 -1562
rect 12812 -1622 12872 -1562
rect 13132 -1622 13192 -1562
rect 13270 -1622 13330 -1562
rect 13590 -1622 13650 -1562
rect 13726 -1622 13786 -1562
rect 14046 -1622 14106 -1562
rect 14182 -1622 14242 -1562
rect 14502 -1622 14562 -1562
rect 14640 -1622 14700 -1562
rect 14960 -1622 15020 -1562
rect 15096 -1622 15156 -1562
rect 15416 -1622 15476 -1562
rect 466 -1972 526 -1912
rect 786 -1972 846 -1912
rect 922 -1972 982 -1912
rect 1242 -1972 1302 -1912
rect 1380 -1972 1440 -1912
rect 1700 -1972 1760 -1912
rect 1836 -1972 1896 -1912
rect 2156 -1972 2216 -1912
rect 2292 -1972 2352 -1912
rect 2612 -1972 2672 -1912
rect 2750 -1972 2810 -1912
rect 3070 -1972 3130 -1912
rect 3206 -1972 3266 -1912
rect 3526 -1972 3586 -1912
rect 3662 -1972 3722 -1912
rect 3982 -1972 4042 -1912
rect 4120 -1972 4180 -1912
rect 4440 -1972 4500 -1912
rect 4576 -1972 4636 -1912
rect 4896 -1972 4956 -1912
rect 5032 -1972 5092 -1912
rect 5352 -1972 5412 -1912
rect 5490 -1972 5550 -1912
rect 5810 -1972 5870 -1912
rect 5946 -1972 6006 -1912
rect 6266 -1972 6326 -1912
rect 6402 -1972 6462 -1912
rect 6722 -1972 6782 -1912
rect 6860 -1972 6920 -1912
rect 7180 -1972 7240 -1912
rect 7316 -1972 7376 -1912
rect 7636 -1972 7696 -1912
rect 7772 -1972 7832 -1912
rect 8092 -1972 8152 -1912
rect 8246 -1972 8306 -1912
rect 8566 -1972 8626 -1912
rect 8702 -1972 8762 -1912
rect 9022 -1972 9082 -1912
rect 9160 -1972 9220 -1912
rect 9480 -1972 9540 -1912
rect 9616 -1972 9676 -1912
rect 9936 -1972 9996 -1912
rect 10072 -1972 10132 -1912
rect 10392 -1972 10452 -1912
rect 10530 -1972 10590 -1912
rect 10850 -1972 10910 -1912
rect 10986 -1972 11046 -1912
rect 11306 -1972 11366 -1912
rect 11442 -1972 11502 -1912
rect 11762 -1972 11822 -1912
rect 11900 -1972 11960 -1912
rect 12220 -1972 12280 -1912
rect 12356 -1972 12416 -1912
rect 12676 -1972 12736 -1912
rect 12812 -1972 12872 -1912
rect 13132 -1972 13192 -1912
rect 13270 -1972 13330 -1912
rect 13590 -1972 13650 -1912
rect 13726 -1972 13786 -1912
rect 14046 -1972 14106 -1912
rect 14182 -1972 14242 -1912
rect 14502 -1972 14562 -1912
rect 14640 -1972 14700 -1912
rect 14960 -1972 15020 -1912
rect 15096 -1972 15156 -1912
rect 15416 -1972 15476 -1912
rect 10 -2124 14 -2064
rect 14 -2124 66 -2064
rect 66 -2124 70 -2064
rect 330 -2124 390 -2064
rect 10 -2474 14 -2414
rect 14 -2474 66 -2414
rect 66 -2474 70 -2414
rect 330 -2474 390 -2414
rect 466 -2124 526 -2064
rect 786 -2124 846 -2064
rect 922 -2124 982 -2064
rect 1242 -2124 1302 -2064
rect 1380 -2124 1440 -2064
rect 1700 -2124 1760 -2064
rect 1836 -2124 1896 -2064
rect 2156 -2124 2216 -2064
rect 2292 -2124 2352 -2064
rect 2612 -2124 2672 -2064
rect 2750 -2124 2810 -2064
rect 3070 -2124 3130 -2064
rect 3206 -2124 3266 -2064
rect 3526 -2124 3586 -2064
rect 3662 -2124 3722 -2064
rect 3982 -2124 4042 -2064
rect 4120 -2124 4180 -2064
rect 4440 -2124 4500 -2064
rect 4576 -2124 4636 -2064
rect 4896 -2124 4956 -2064
rect 5032 -2124 5092 -2064
rect 5352 -2124 5412 -2064
rect 5490 -2124 5550 -2064
rect 5810 -2124 5870 -2064
rect 5946 -2124 6006 -2064
rect 6266 -2124 6326 -2064
rect 6402 -2124 6462 -2064
rect 6722 -2124 6782 -2064
rect 6860 -2124 6920 -2064
rect 7180 -2124 7240 -2064
rect 7316 -2124 7376 -2064
rect 7636 -2124 7696 -2064
rect 7772 -2124 7832 -2064
rect 8092 -2124 8152 -2064
rect 8246 -2124 8306 -2064
rect 8566 -2124 8626 -2064
rect 8702 -2124 8762 -2064
rect 9022 -2124 9082 -2064
rect 9160 -2124 9220 -2064
rect 9480 -2124 9540 -2064
rect 9616 -2124 9676 -2064
rect 9936 -2124 9996 -2064
rect 10072 -2124 10132 -2064
rect 10392 -2124 10452 -2064
rect 10530 -2124 10590 -2064
rect 10850 -2124 10910 -2064
rect 10986 -2124 11046 -2064
rect 11306 -2124 11366 -2064
rect 11442 -2124 11502 -2064
rect 11762 -2124 11822 -2064
rect 11900 -2124 11960 -2064
rect 12220 -2124 12280 -2064
rect 12356 -2124 12416 -2064
rect 12676 -2124 12736 -2064
rect 12812 -2124 12872 -2064
rect 13132 -2124 13192 -2064
rect 13270 -2124 13330 -2064
rect 13590 -2124 13650 -2064
rect 13726 -2124 13786 -2064
rect 14046 -2124 14106 -2064
rect 14182 -2124 14242 -2064
rect 14502 -2124 14562 -2064
rect 14640 -2124 14700 -2064
rect 14960 -2124 15020 -2064
rect 15096 -2124 15156 -2064
rect 15416 -2124 15476 -2064
rect 466 -2474 526 -2414
rect 786 -2474 846 -2414
rect 922 -2474 982 -2414
rect 1242 -2474 1302 -2414
rect 1380 -2474 1440 -2414
rect 1700 -2474 1760 -2414
rect 1836 -2474 1896 -2414
rect 2156 -2474 2216 -2414
rect 2292 -2474 2352 -2414
rect 2612 -2474 2672 -2414
rect 2750 -2474 2810 -2414
rect 3070 -2474 3130 -2414
rect 3206 -2474 3266 -2414
rect 3526 -2474 3586 -2414
rect 3662 -2474 3722 -2414
rect 3982 -2474 4042 -2414
rect 4120 -2474 4180 -2414
rect 4440 -2474 4500 -2414
rect 4576 -2474 4636 -2414
rect 4896 -2474 4956 -2414
rect 5032 -2474 5092 -2414
rect 5352 -2474 5412 -2414
rect 5490 -2474 5550 -2414
rect 5810 -2474 5870 -2414
rect 5946 -2474 6006 -2414
rect 6266 -2474 6326 -2414
rect 6402 -2474 6462 -2414
rect 6722 -2474 6782 -2414
rect 6860 -2474 6920 -2414
rect 7180 -2474 7240 -2414
rect 7316 -2474 7376 -2414
rect 7636 -2474 7696 -2414
rect 7772 -2474 7832 -2414
rect 8092 -2474 8152 -2414
rect 8246 -2474 8306 -2414
rect 8566 -2474 8626 -2414
rect 8702 -2474 8762 -2414
rect 9022 -2474 9082 -2414
rect 9160 -2474 9220 -2414
rect 9480 -2474 9540 -2414
rect 9616 -2474 9676 -2414
rect 9936 -2474 9996 -2414
rect 10072 -2474 10132 -2414
rect 10392 -2474 10452 -2414
rect 10530 -2474 10590 -2414
rect 10850 -2474 10910 -2414
rect 10986 -2474 11046 -2414
rect 11306 -2474 11366 -2414
rect 11442 -2474 11502 -2414
rect 11762 -2474 11822 -2414
rect 11900 -2474 11960 -2414
rect 12220 -2474 12280 -2414
rect 12356 -2474 12416 -2414
rect 12676 -2474 12736 -2414
rect 12812 -2474 12872 -2414
rect 13132 -2474 13192 -2414
rect 13270 -2474 13330 -2414
rect 13590 -2474 13650 -2414
rect 13726 -2474 13786 -2414
rect 14046 -2474 14106 -2414
rect 14182 -2474 14242 -2414
rect 14502 -2474 14562 -2414
rect 14640 -2474 14700 -2414
rect 14960 -2474 15020 -2414
rect 15096 -2474 15156 -2414
rect 15416 -2474 15476 -2414
rect 10 -2616 14 -2556
rect 14 -2616 66 -2556
rect 66 -2616 70 -2556
rect 330 -2616 390 -2556
rect 10 -2966 14 -2906
rect 14 -2966 66 -2906
rect 66 -2966 70 -2906
rect 330 -2966 390 -2906
rect 466 -2616 526 -2556
rect 786 -2616 846 -2556
rect 922 -2616 982 -2556
rect 1242 -2616 1302 -2556
rect 1380 -2616 1440 -2556
rect 1700 -2616 1760 -2556
rect 1836 -2616 1896 -2556
rect 2156 -2616 2216 -2556
rect 2292 -2616 2352 -2556
rect 2612 -2616 2672 -2556
rect 2750 -2616 2810 -2556
rect 3070 -2616 3130 -2556
rect 3206 -2616 3266 -2556
rect 3526 -2616 3586 -2556
rect 3662 -2616 3722 -2556
rect 3982 -2616 4042 -2556
rect 4120 -2616 4180 -2556
rect 4440 -2616 4500 -2556
rect 4576 -2616 4636 -2556
rect 4896 -2616 4956 -2556
rect 5032 -2616 5092 -2556
rect 5352 -2616 5412 -2556
rect 5490 -2616 5550 -2556
rect 5810 -2616 5870 -2556
rect 5946 -2616 6006 -2556
rect 6266 -2616 6326 -2556
rect 6402 -2616 6462 -2556
rect 6722 -2616 6782 -2556
rect 6860 -2616 6920 -2556
rect 7180 -2616 7240 -2556
rect 7316 -2616 7376 -2556
rect 7636 -2616 7696 -2556
rect 7772 -2616 7832 -2556
rect 8092 -2616 8152 -2556
rect 8246 -2616 8306 -2556
rect 8566 -2616 8626 -2556
rect 8702 -2616 8762 -2556
rect 9022 -2616 9082 -2556
rect 9160 -2616 9220 -2556
rect 9480 -2616 9540 -2556
rect 9616 -2616 9676 -2556
rect 9936 -2616 9996 -2556
rect 10072 -2616 10132 -2556
rect 10392 -2616 10452 -2556
rect 10530 -2616 10590 -2556
rect 10850 -2616 10910 -2556
rect 10986 -2616 11046 -2556
rect 11306 -2616 11366 -2556
rect 11442 -2616 11502 -2556
rect 11762 -2616 11822 -2556
rect 11900 -2616 11960 -2556
rect 12220 -2616 12280 -2556
rect 12356 -2616 12416 -2556
rect 12676 -2616 12736 -2556
rect 12812 -2616 12872 -2556
rect 13132 -2616 13192 -2556
rect 13270 -2616 13330 -2556
rect 13590 -2616 13650 -2556
rect 13726 -2616 13786 -2556
rect 14046 -2616 14106 -2556
rect 14182 -2616 14242 -2556
rect 14502 -2616 14562 -2556
rect 14640 -2616 14700 -2556
rect 14960 -2616 15020 -2556
rect 15096 -2616 15156 -2556
rect 15416 -2616 15476 -2556
rect 466 -2966 526 -2906
rect 786 -2966 846 -2906
rect 922 -2966 982 -2906
rect 1242 -2966 1302 -2906
rect 1380 -2966 1440 -2906
rect 1700 -2966 1760 -2906
rect 1836 -2966 1896 -2906
rect 2156 -2966 2216 -2906
rect 2292 -2966 2352 -2906
rect 2612 -2966 2672 -2906
rect 2750 -2966 2810 -2906
rect 3070 -2966 3130 -2906
rect 3206 -2966 3266 -2906
rect 3526 -2966 3586 -2906
rect 3662 -2966 3722 -2906
rect 3982 -2966 4042 -2906
rect 4120 -2966 4180 -2906
rect 4440 -2966 4500 -2906
rect 4576 -2966 4636 -2906
rect 4896 -2966 4956 -2906
rect 5032 -2966 5092 -2906
rect 5352 -2966 5412 -2906
rect 5490 -2966 5550 -2906
rect 5810 -2966 5870 -2906
rect 5946 -2966 6006 -2906
rect 6266 -2966 6326 -2906
rect 6402 -2966 6462 -2906
rect 6722 -2966 6782 -2906
rect 6860 -2966 6920 -2906
rect 7180 -2966 7240 -2906
rect 7316 -2966 7376 -2906
rect 7636 -2966 7696 -2906
rect 7772 -2966 7832 -2906
rect 8092 -2966 8152 -2906
rect 8246 -2966 8306 -2906
rect 8566 -2966 8626 -2906
rect 8702 -2966 8762 -2906
rect 9022 -2966 9082 -2906
rect 9160 -2966 9220 -2906
rect 9480 -2966 9540 -2906
rect 9616 -2966 9676 -2906
rect 9936 -2966 9996 -2906
rect 10072 -2966 10132 -2906
rect 10392 -2966 10452 -2906
rect 10530 -2966 10590 -2906
rect 10850 -2966 10910 -2906
rect 10986 -2966 11046 -2906
rect 11306 -2966 11366 -2906
rect 11442 -2966 11502 -2906
rect 11762 -2966 11822 -2906
rect 11900 -2966 11960 -2906
rect 12220 -2966 12280 -2906
rect 12356 -2966 12416 -2906
rect 12676 -2966 12736 -2906
rect 12812 -2966 12872 -2906
rect 13132 -2966 13192 -2906
rect 13270 -2966 13330 -2906
rect 13590 -2966 13650 -2906
rect 13726 -2966 13786 -2906
rect 14046 -2966 14106 -2906
rect 14182 -2966 14242 -2906
rect 14502 -2966 14562 -2906
rect 14640 -2966 14700 -2906
rect 14960 -2966 15020 -2906
rect 15096 -2966 15156 -2906
rect 15416 -2966 15476 -2906
rect 10 -3612 14 -3552
rect 14 -3612 66 -3552
rect 66 -3612 70 -3552
rect 330 -3612 390 -3552
rect 10 -3962 14 -3902
rect 14 -3962 66 -3902
rect 66 -3962 70 -3902
rect 330 -3962 390 -3902
rect 466 -3612 526 -3552
rect 786 -3612 846 -3552
rect 922 -3612 982 -3552
rect 1242 -3612 1302 -3552
rect 1380 -3612 1440 -3552
rect 1700 -3612 1760 -3552
rect 1836 -3612 1896 -3552
rect 2156 -3612 2216 -3552
rect 2292 -3612 2352 -3552
rect 2612 -3612 2672 -3552
rect 2750 -3612 2810 -3552
rect 3070 -3612 3130 -3552
rect 3206 -3612 3266 -3552
rect 3526 -3612 3586 -3552
rect 3662 -3612 3722 -3552
rect 3982 -3612 4042 -3552
rect 4120 -3612 4180 -3552
rect 4440 -3612 4500 -3552
rect 4576 -3612 4636 -3552
rect 4896 -3612 4956 -3552
rect 5032 -3612 5092 -3552
rect 5352 -3612 5412 -3552
rect 5490 -3612 5550 -3552
rect 5810 -3612 5870 -3552
rect 5946 -3612 6006 -3552
rect 6266 -3612 6326 -3552
rect 6402 -3612 6462 -3552
rect 6722 -3612 6782 -3552
rect 6860 -3612 6920 -3552
rect 7180 -3612 7240 -3552
rect 7316 -3612 7376 -3552
rect 7636 -3612 7696 -3552
rect 7772 -3612 7832 -3552
rect 8092 -3612 8152 -3552
rect 8246 -3612 8306 -3552
rect 8566 -3612 8626 -3552
rect 8702 -3612 8762 -3552
rect 9022 -3612 9082 -3552
rect 9160 -3612 9220 -3552
rect 9480 -3612 9540 -3552
rect 9616 -3612 9676 -3552
rect 9936 -3612 9996 -3552
rect 10072 -3612 10132 -3552
rect 10392 -3612 10452 -3552
rect 10530 -3612 10590 -3552
rect 10850 -3612 10910 -3552
rect 10986 -3612 11046 -3552
rect 11306 -3612 11366 -3552
rect 11442 -3612 11502 -3552
rect 11762 -3612 11822 -3552
rect 11900 -3612 11960 -3552
rect 12220 -3612 12280 -3552
rect 12356 -3612 12416 -3552
rect 12676 -3612 12736 -3552
rect 12812 -3612 12872 -3552
rect 13132 -3612 13192 -3552
rect 13270 -3612 13330 -3552
rect 13590 -3612 13650 -3552
rect 13726 -3612 13786 -3552
rect 14046 -3612 14106 -3552
rect 14182 -3612 14242 -3552
rect 14502 -3612 14562 -3552
rect 14640 -3612 14700 -3552
rect 14960 -3612 15020 -3552
rect 15096 -3612 15156 -3552
rect 15416 -3612 15476 -3552
rect 466 -3962 526 -3902
rect 786 -3962 846 -3902
rect 922 -3962 982 -3902
rect 1242 -3962 1302 -3902
rect 1380 -3962 1440 -3902
rect 1700 -3962 1760 -3902
rect 1836 -3962 1896 -3902
rect 2156 -3962 2216 -3902
rect 2292 -3962 2352 -3902
rect 2612 -3962 2672 -3902
rect 2750 -3962 2810 -3902
rect 3070 -3962 3130 -3902
rect 3206 -3962 3266 -3902
rect 3526 -3962 3586 -3902
rect 3662 -3962 3722 -3902
rect 3982 -3962 4042 -3902
rect 4120 -3962 4180 -3902
rect 4440 -3962 4500 -3902
rect 4576 -3962 4636 -3902
rect 4896 -3962 4956 -3902
rect 5032 -3962 5092 -3902
rect 5352 -3962 5412 -3902
rect 5490 -3962 5550 -3902
rect 5810 -3962 5870 -3902
rect 5946 -3962 6006 -3902
rect 6266 -3962 6326 -3902
rect 6402 -3962 6462 -3902
rect 6722 -3962 6782 -3902
rect 6860 -3962 6920 -3902
rect 7180 -3962 7240 -3902
rect 7316 -3962 7376 -3902
rect 7636 -3962 7696 -3902
rect 7772 -3962 7832 -3902
rect 8092 -3962 8152 -3902
rect 8246 -3962 8306 -3902
rect 8566 -3962 8626 -3902
rect 8702 -3962 8762 -3902
rect 9022 -3962 9082 -3902
rect 9160 -3962 9220 -3902
rect 9480 -3962 9540 -3902
rect 9616 -3962 9676 -3902
rect 9936 -3962 9996 -3902
rect 10072 -3962 10132 -3902
rect 10392 -3962 10452 -3902
rect 10530 -3962 10590 -3902
rect 10850 -3962 10910 -3902
rect 10986 -3962 11046 -3902
rect 11306 -3962 11366 -3902
rect 11442 -3962 11502 -3902
rect 11762 -3962 11822 -3902
rect 11900 -3962 11960 -3902
rect 12220 -3962 12280 -3902
rect 12356 -3962 12416 -3902
rect 12676 -3962 12736 -3902
rect 12812 -3962 12872 -3902
rect 13132 -3962 13192 -3902
rect 13270 -3962 13330 -3902
rect 13590 -3962 13650 -3902
rect 13726 -3962 13786 -3902
rect 14046 -3962 14106 -3902
rect 14182 -3962 14242 -3902
rect 14502 -3962 14562 -3902
rect 14640 -3962 14700 -3902
rect 14960 -3962 15020 -3902
rect 15096 -3962 15156 -3902
rect 15416 -3962 15476 -3902
rect 10 -4104 14 -4044
rect 14 -4104 66 -4044
rect 66 -4104 70 -4044
rect 330 -4104 390 -4044
rect 10 -4454 14 -4394
rect 14 -4454 66 -4394
rect 66 -4454 70 -4394
rect 330 -4454 390 -4394
rect 466 -4104 526 -4044
rect 786 -4104 846 -4044
rect 922 -4104 982 -4044
rect 1242 -4104 1302 -4044
rect 1380 -4104 1440 -4044
rect 1700 -4104 1760 -4044
rect 1836 -4104 1896 -4044
rect 2156 -4104 2216 -4044
rect 2292 -4104 2352 -4044
rect 2612 -4104 2672 -4044
rect 2750 -4104 2810 -4044
rect 3070 -4104 3130 -4044
rect 3206 -4104 3266 -4044
rect 3526 -4104 3586 -4044
rect 3662 -4104 3722 -4044
rect 3982 -4104 4042 -4044
rect 4120 -4104 4180 -4044
rect 4440 -4104 4500 -4044
rect 4576 -4104 4636 -4044
rect 4896 -4104 4956 -4044
rect 5032 -4104 5092 -4044
rect 5352 -4104 5412 -4044
rect 5490 -4104 5550 -4044
rect 5810 -4104 5870 -4044
rect 5946 -4104 6006 -4044
rect 6266 -4104 6326 -4044
rect 6402 -4104 6462 -4044
rect 6722 -4104 6782 -4044
rect 6860 -4104 6920 -4044
rect 7180 -4104 7240 -4044
rect 7316 -4104 7376 -4044
rect 7636 -4104 7696 -4044
rect 7772 -4104 7832 -4044
rect 8092 -4104 8152 -4044
rect 8246 -4104 8306 -4044
rect 8566 -4104 8626 -4044
rect 8702 -4104 8762 -4044
rect 9022 -4104 9082 -4044
rect 9160 -4104 9220 -4044
rect 9480 -4104 9540 -4044
rect 9616 -4104 9676 -4044
rect 9936 -4104 9996 -4044
rect 10072 -4104 10132 -4044
rect 10392 -4104 10452 -4044
rect 10530 -4104 10590 -4044
rect 10850 -4104 10910 -4044
rect 10986 -4104 11046 -4044
rect 11306 -4104 11366 -4044
rect 11442 -4104 11502 -4044
rect 11762 -4104 11822 -4044
rect 11900 -4104 11960 -4044
rect 12220 -4104 12280 -4044
rect 12356 -4104 12416 -4044
rect 12676 -4104 12736 -4044
rect 12812 -4104 12872 -4044
rect 13132 -4104 13192 -4044
rect 13270 -4104 13330 -4044
rect 13590 -4104 13650 -4044
rect 13726 -4104 13786 -4044
rect 14046 -4104 14106 -4044
rect 14182 -4104 14242 -4044
rect 14502 -4104 14562 -4044
rect 14640 -4104 14700 -4044
rect 14960 -4104 15020 -4044
rect 15096 -4104 15156 -4044
rect 15416 -4104 15476 -4044
rect 466 -4454 526 -4394
rect 786 -4454 846 -4394
rect 922 -4454 982 -4394
rect 1242 -4454 1302 -4394
rect 1380 -4454 1440 -4394
rect 1700 -4454 1760 -4394
rect 1836 -4454 1896 -4394
rect 2156 -4454 2216 -4394
rect 2292 -4454 2352 -4394
rect 2612 -4454 2672 -4394
rect 2750 -4454 2810 -4394
rect 3070 -4454 3130 -4394
rect 3206 -4454 3266 -4394
rect 3526 -4454 3586 -4394
rect 3662 -4454 3722 -4394
rect 3982 -4454 4042 -4394
rect 4120 -4454 4180 -4394
rect 4440 -4454 4500 -4394
rect 4576 -4454 4636 -4394
rect 4896 -4454 4956 -4394
rect 5032 -4454 5092 -4394
rect 5352 -4454 5412 -4394
rect 5490 -4454 5550 -4394
rect 5810 -4454 5870 -4394
rect 5946 -4454 6006 -4394
rect 6266 -4454 6326 -4394
rect 6402 -4454 6462 -4394
rect 6722 -4454 6782 -4394
rect 6860 -4454 6920 -4394
rect 7180 -4454 7240 -4394
rect 7316 -4454 7376 -4394
rect 7636 -4454 7696 -4394
rect 7772 -4454 7832 -4394
rect 8092 -4454 8152 -4394
rect 8246 -4454 8306 -4394
rect 8566 -4454 8626 -4394
rect 8702 -4454 8762 -4394
rect 9022 -4454 9082 -4394
rect 9160 -4454 9220 -4394
rect 9480 -4454 9540 -4394
rect 9616 -4454 9676 -4394
rect 9936 -4454 9996 -4394
rect 10072 -4454 10132 -4394
rect 10392 -4454 10452 -4394
rect 10530 -4454 10590 -4394
rect 10850 -4454 10910 -4394
rect 10986 -4454 11046 -4394
rect 11306 -4454 11366 -4394
rect 11442 -4454 11502 -4394
rect 11762 -4454 11822 -4394
rect 11900 -4454 11960 -4394
rect 12220 -4454 12280 -4394
rect 12356 -4454 12416 -4394
rect 12676 -4454 12736 -4394
rect 12812 -4454 12872 -4394
rect 13132 -4454 13192 -4394
rect 13270 -4454 13330 -4394
rect 13590 -4454 13650 -4394
rect 13726 -4454 13786 -4394
rect 14046 -4454 14106 -4394
rect 14182 -4454 14242 -4394
rect 14502 -4454 14562 -4394
rect 14640 -4454 14700 -4394
rect 14960 -4454 15020 -4394
rect 15096 -4454 15156 -4394
rect 15416 -4454 15476 -4394
rect 10 -4620 14 -4560
rect 14 -4620 66 -4560
rect 66 -4620 70 -4560
rect 330 -4620 390 -4560
rect 10 -4970 14 -4910
rect 14 -4970 66 -4910
rect 66 -4970 70 -4910
rect 330 -4970 390 -4910
rect 466 -4620 526 -4560
rect 786 -4620 846 -4560
rect 922 -4620 982 -4560
rect 1242 -4620 1302 -4560
rect 1380 -4620 1440 -4560
rect 1700 -4620 1760 -4560
rect 1836 -4620 1896 -4560
rect 2156 -4620 2216 -4560
rect 2292 -4620 2352 -4560
rect 2612 -4620 2672 -4560
rect 2750 -4620 2810 -4560
rect 3070 -4620 3130 -4560
rect 3206 -4620 3266 -4560
rect 3526 -4620 3586 -4560
rect 3662 -4620 3722 -4560
rect 3982 -4620 4042 -4560
rect 4120 -4620 4180 -4560
rect 4440 -4620 4500 -4560
rect 4576 -4620 4636 -4560
rect 4896 -4620 4956 -4560
rect 5032 -4620 5092 -4560
rect 5352 -4620 5412 -4560
rect 5490 -4620 5550 -4560
rect 5810 -4620 5870 -4560
rect 5946 -4620 6006 -4560
rect 6266 -4620 6326 -4560
rect 6402 -4620 6462 -4560
rect 6722 -4620 6782 -4560
rect 6860 -4620 6920 -4560
rect 7180 -4620 7240 -4560
rect 7316 -4620 7376 -4560
rect 7636 -4620 7696 -4560
rect 7772 -4620 7832 -4560
rect 8092 -4620 8152 -4560
rect 8246 -4620 8306 -4560
rect 8566 -4620 8626 -4560
rect 8702 -4620 8762 -4560
rect 9022 -4620 9082 -4560
rect 9160 -4620 9220 -4560
rect 9480 -4620 9540 -4560
rect 9616 -4620 9676 -4560
rect 9936 -4620 9996 -4560
rect 10072 -4620 10132 -4560
rect 10392 -4620 10452 -4560
rect 10530 -4620 10590 -4560
rect 10850 -4620 10910 -4560
rect 10986 -4620 11046 -4560
rect 11306 -4620 11366 -4560
rect 11442 -4620 11502 -4560
rect 11762 -4620 11822 -4560
rect 11900 -4620 11960 -4560
rect 12220 -4620 12280 -4560
rect 12356 -4620 12416 -4560
rect 12676 -4620 12736 -4560
rect 12812 -4620 12872 -4560
rect 13132 -4620 13192 -4560
rect 13270 -4620 13330 -4560
rect 13590 -4620 13650 -4560
rect 13726 -4620 13786 -4560
rect 14046 -4620 14106 -4560
rect 14182 -4620 14242 -4560
rect 14502 -4620 14562 -4560
rect 14640 -4620 14700 -4560
rect 14960 -4620 15020 -4560
rect 15096 -4620 15156 -4560
rect 15416 -4620 15476 -4560
rect 466 -4970 526 -4910
rect 786 -4970 846 -4910
rect 922 -4970 982 -4910
rect 1242 -4970 1302 -4910
rect 1380 -4970 1440 -4910
rect 1700 -4970 1760 -4910
rect 1836 -4970 1896 -4910
rect 2156 -4970 2216 -4910
rect 2292 -4970 2352 -4910
rect 2612 -4970 2672 -4910
rect 2750 -4970 2810 -4910
rect 3070 -4970 3130 -4910
rect 3206 -4970 3266 -4910
rect 3526 -4970 3586 -4910
rect 3662 -4970 3722 -4910
rect 3982 -4970 4042 -4910
rect 4120 -4970 4180 -4910
rect 4440 -4970 4500 -4910
rect 4576 -4970 4636 -4910
rect 4896 -4970 4956 -4910
rect 5032 -4970 5092 -4910
rect 5352 -4970 5412 -4910
rect 5490 -4970 5550 -4910
rect 5810 -4970 5870 -4910
rect 5946 -4970 6006 -4910
rect 6266 -4970 6326 -4910
rect 6402 -4970 6462 -4910
rect 6722 -4970 6782 -4910
rect 6860 -4970 6920 -4910
rect 7180 -4970 7240 -4910
rect 7316 -4970 7376 -4910
rect 7636 -4970 7696 -4910
rect 7772 -4970 7832 -4910
rect 8092 -4970 8152 -4910
rect 8246 -4970 8306 -4910
rect 8566 -4970 8626 -4910
rect 8702 -4970 8762 -4910
rect 9022 -4970 9082 -4910
rect 9160 -4970 9220 -4910
rect 9480 -4970 9540 -4910
rect 9616 -4970 9676 -4910
rect 9936 -4970 9996 -4910
rect 10072 -4970 10132 -4910
rect 10392 -4970 10452 -4910
rect 10530 -4970 10590 -4910
rect 10850 -4970 10910 -4910
rect 10986 -4970 11046 -4910
rect 11306 -4970 11366 -4910
rect 11442 -4970 11502 -4910
rect 11762 -4970 11822 -4910
rect 11900 -4970 11960 -4910
rect 12220 -4970 12280 -4910
rect 12356 -4970 12416 -4910
rect 12676 -4970 12736 -4910
rect 12812 -4970 12872 -4910
rect 13132 -4970 13192 -4910
rect 13270 -4970 13330 -4910
rect 13590 -4970 13650 -4910
rect 13726 -4970 13786 -4910
rect 14046 -4970 14106 -4910
rect 14182 -4970 14242 -4910
rect 14502 -4970 14562 -4910
rect 14640 -4970 14700 -4910
rect 14960 -4970 15020 -4910
rect 15096 -4970 15156 -4910
rect 15416 -4970 15476 -4910
rect 10 -5122 14 -5062
rect 14 -5122 66 -5062
rect 66 -5122 70 -5062
rect 330 -5122 390 -5062
rect 10 -5472 14 -5412
rect 14 -5472 66 -5412
rect 66 -5472 70 -5412
rect 330 -5472 390 -5412
rect 466 -5122 526 -5062
rect 786 -5122 846 -5062
rect 922 -5122 982 -5062
rect 1242 -5122 1302 -5062
rect 1380 -5122 1440 -5062
rect 1700 -5122 1760 -5062
rect 1836 -5122 1896 -5062
rect 2156 -5122 2216 -5062
rect 2292 -5122 2352 -5062
rect 2612 -5122 2672 -5062
rect 2750 -5122 2810 -5062
rect 3070 -5122 3130 -5062
rect 3206 -5122 3266 -5062
rect 3526 -5122 3586 -5062
rect 3662 -5122 3722 -5062
rect 3982 -5122 4042 -5062
rect 4120 -5122 4180 -5062
rect 4440 -5122 4500 -5062
rect 4576 -5122 4636 -5062
rect 4896 -5122 4956 -5062
rect 5032 -5122 5092 -5062
rect 5352 -5122 5412 -5062
rect 5490 -5122 5550 -5062
rect 5810 -5122 5870 -5062
rect 5946 -5122 6006 -5062
rect 6266 -5122 6326 -5062
rect 6402 -5122 6462 -5062
rect 6722 -5122 6782 -5062
rect 6860 -5122 6920 -5062
rect 7180 -5122 7240 -5062
rect 7316 -5122 7376 -5062
rect 7636 -5122 7696 -5062
rect 7772 -5122 7832 -5062
rect 8092 -5122 8152 -5062
rect 8246 -5122 8306 -5062
rect 8566 -5122 8626 -5062
rect 8702 -5122 8762 -5062
rect 9022 -5122 9082 -5062
rect 9160 -5122 9220 -5062
rect 9480 -5122 9540 -5062
rect 9616 -5122 9676 -5062
rect 9936 -5122 9996 -5062
rect 10072 -5122 10132 -5062
rect 10392 -5122 10452 -5062
rect 10530 -5122 10590 -5062
rect 10850 -5122 10910 -5062
rect 10986 -5122 11046 -5062
rect 11306 -5122 11366 -5062
rect 11442 -5122 11502 -5062
rect 11762 -5122 11822 -5062
rect 11900 -5122 11960 -5062
rect 12220 -5122 12280 -5062
rect 12356 -5122 12416 -5062
rect 12676 -5122 12736 -5062
rect 12812 -5122 12872 -5062
rect 13132 -5122 13192 -5062
rect 13270 -5122 13330 -5062
rect 13590 -5122 13650 -5062
rect 13726 -5122 13786 -5062
rect 14046 -5122 14106 -5062
rect 14182 -5122 14242 -5062
rect 14502 -5122 14562 -5062
rect 14640 -5122 14700 -5062
rect 14960 -5122 15020 -5062
rect 15096 -5122 15156 -5062
rect 15416 -5122 15476 -5062
rect 466 -5472 526 -5412
rect 786 -5472 846 -5412
rect 922 -5472 982 -5412
rect 1242 -5472 1302 -5412
rect 1380 -5472 1440 -5412
rect 1700 -5472 1760 -5412
rect 1836 -5472 1896 -5412
rect 2156 -5472 2216 -5412
rect 2292 -5472 2352 -5412
rect 2612 -5472 2672 -5412
rect 2750 -5472 2810 -5412
rect 3070 -5472 3130 -5412
rect 3206 -5472 3266 -5412
rect 3526 -5472 3586 -5412
rect 3662 -5472 3722 -5412
rect 3982 -5472 4042 -5412
rect 4120 -5472 4180 -5412
rect 4440 -5472 4500 -5412
rect 4576 -5472 4636 -5412
rect 4896 -5472 4956 -5412
rect 5032 -5472 5092 -5412
rect 5352 -5472 5412 -5412
rect 5490 -5472 5550 -5412
rect 5810 -5472 5870 -5412
rect 5946 -5472 6006 -5412
rect 6266 -5472 6326 -5412
rect 6402 -5472 6462 -5412
rect 6722 -5472 6782 -5412
rect 6860 -5472 6920 -5412
rect 7180 -5472 7240 -5412
rect 7316 -5472 7376 -5412
rect 7636 -5472 7696 -5412
rect 7772 -5472 7832 -5412
rect 8092 -5472 8152 -5412
rect 8246 -5472 8306 -5412
rect 8566 -5472 8626 -5412
rect 8702 -5472 8762 -5412
rect 9022 -5472 9082 -5412
rect 9160 -5472 9220 -5412
rect 9480 -5472 9540 -5412
rect 9616 -5472 9676 -5412
rect 9936 -5472 9996 -5412
rect 10072 -5472 10132 -5412
rect 10392 -5472 10452 -5412
rect 10530 -5472 10590 -5412
rect 10850 -5472 10910 -5412
rect 10986 -5472 11046 -5412
rect 11306 -5472 11366 -5412
rect 11442 -5472 11502 -5412
rect 11762 -5472 11822 -5412
rect 11900 -5472 11960 -5412
rect 12220 -5472 12280 -5412
rect 12356 -5472 12416 -5412
rect 12676 -5472 12736 -5412
rect 12812 -5472 12872 -5412
rect 13132 -5472 13192 -5412
rect 13270 -5472 13330 -5412
rect 13590 -5472 13650 -5412
rect 13726 -5472 13786 -5412
rect 14046 -5472 14106 -5412
rect 14182 -5472 14242 -5412
rect 14502 -5472 14562 -5412
rect 14640 -5472 14700 -5412
rect 14960 -5472 15020 -5412
rect 15096 -5472 15156 -5412
rect 15416 -5472 15476 -5412
rect 10 -5614 14 -5554
rect 14 -5614 66 -5554
rect 66 -5614 70 -5554
rect 330 -5614 390 -5554
rect 10 -5964 14 -5904
rect 14 -5964 66 -5904
rect 66 -5964 70 -5904
rect 330 -5964 390 -5904
rect 466 -5614 526 -5554
rect 786 -5614 846 -5554
rect 922 -5614 982 -5554
rect 1242 -5614 1302 -5554
rect 1380 -5614 1440 -5554
rect 1700 -5614 1760 -5554
rect 1836 -5614 1896 -5554
rect 2156 -5614 2216 -5554
rect 2292 -5614 2352 -5554
rect 2612 -5614 2672 -5554
rect 2750 -5614 2810 -5554
rect 3070 -5614 3130 -5554
rect 3206 -5614 3266 -5554
rect 3526 -5614 3586 -5554
rect 3662 -5614 3722 -5554
rect 3982 -5614 4042 -5554
rect 4120 -5614 4180 -5554
rect 4440 -5614 4500 -5554
rect 4576 -5614 4636 -5554
rect 4896 -5614 4956 -5554
rect 5032 -5614 5092 -5554
rect 5352 -5614 5412 -5554
rect 5490 -5614 5550 -5554
rect 5810 -5614 5870 -5554
rect 5946 -5614 6006 -5554
rect 6266 -5614 6326 -5554
rect 6402 -5614 6462 -5554
rect 6722 -5614 6782 -5554
rect 6860 -5614 6920 -5554
rect 7180 -5614 7240 -5554
rect 7316 -5614 7376 -5554
rect 7636 -5614 7696 -5554
rect 7772 -5614 7832 -5554
rect 8092 -5614 8152 -5554
rect 8246 -5614 8306 -5554
rect 8566 -5614 8626 -5554
rect 8702 -5614 8762 -5554
rect 9022 -5614 9082 -5554
rect 9160 -5614 9220 -5554
rect 9480 -5614 9540 -5554
rect 9616 -5614 9676 -5554
rect 9936 -5614 9996 -5554
rect 10072 -5614 10132 -5554
rect 10392 -5614 10452 -5554
rect 10530 -5614 10590 -5554
rect 10850 -5614 10910 -5554
rect 10986 -5614 11046 -5554
rect 11306 -5614 11366 -5554
rect 11442 -5614 11502 -5554
rect 11762 -5614 11822 -5554
rect 11900 -5614 11960 -5554
rect 12220 -5614 12280 -5554
rect 12356 -5614 12416 -5554
rect 12676 -5614 12736 -5554
rect 12812 -5614 12872 -5554
rect 13132 -5614 13192 -5554
rect 13270 -5614 13330 -5554
rect 13590 -5614 13650 -5554
rect 13726 -5614 13786 -5554
rect 14046 -5614 14106 -5554
rect 14182 -5614 14242 -5554
rect 14502 -5614 14562 -5554
rect 14640 -5614 14700 -5554
rect 14960 -5614 15020 -5554
rect 15096 -5614 15156 -5554
rect 15416 -5614 15476 -5554
rect 466 -5964 526 -5904
rect 786 -5964 846 -5904
rect 922 -5964 982 -5904
rect 1242 -5964 1302 -5904
rect 1380 -5964 1440 -5904
rect 1700 -5964 1760 -5904
rect 1836 -5964 1896 -5904
rect 2156 -5964 2216 -5904
rect 2292 -5964 2352 -5904
rect 2612 -5964 2672 -5904
rect 2750 -5964 2810 -5904
rect 3070 -5964 3130 -5904
rect 3206 -5964 3266 -5904
rect 3526 -5964 3586 -5904
rect 3662 -5964 3722 -5904
rect 3982 -5964 4042 -5904
rect 4120 -5964 4180 -5904
rect 4440 -5964 4500 -5904
rect 4576 -5964 4636 -5904
rect 4896 -5964 4956 -5904
rect 5032 -5964 5092 -5904
rect 5352 -5964 5412 -5904
rect 5490 -5964 5550 -5904
rect 5810 -5964 5870 -5904
rect 5946 -5964 6006 -5904
rect 6266 -5964 6326 -5904
rect 6402 -5964 6462 -5904
rect 6722 -5964 6782 -5904
rect 6860 -5964 6920 -5904
rect 7180 -5964 7240 -5904
rect 7316 -5964 7376 -5904
rect 7636 -5964 7696 -5904
rect 7772 -5964 7832 -5904
rect 8092 -5964 8152 -5904
rect 8246 -5964 8306 -5904
rect 8566 -5964 8626 -5904
rect 8702 -5964 8762 -5904
rect 9022 -5964 9082 -5904
rect 9160 -5964 9220 -5904
rect 9480 -5964 9540 -5904
rect 9616 -5964 9676 -5904
rect 9936 -5964 9996 -5904
rect 10072 -5964 10132 -5904
rect 10392 -5964 10452 -5904
rect 10530 -5964 10590 -5904
rect 10850 -5964 10910 -5904
rect 10986 -5964 11046 -5904
rect 11306 -5964 11366 -5904
rect 11442 -5964 11502 -5904
rect 11762 -5964 11822 -5904
rect 11900 -5964 11960 -5904
rect 12220 -5964 12280 -5904
rect 12356 -5964 12416 -5904
rect 12676 -5964 12736 -5904
rect 12812 -5964 12872 -5904
rect 13132 -5964 13192 -5904
rect 13270 -5964 13330 -5904
rect 13590 -5964 13650 -5904
rect 13726 -5964 13786 -5904
rect 14046 -5964 14106 -5904
rect 14182 -5964 14242 -5904
rect 14502 -5964 14562 -5904
rect 14640 -5964 14700 -5904
rect 14960 -5964 15020 -5904
rect 15096 -5964 15156 -5904
rect 15416 -5964 15476 -5904
rect 11 -6111 14 -6051
rect 14 -6111 66 -6051
rect 66 -6111 71 -6051
rect 331 -6111 391 -6051
rect 11 -6461 14 -6401
rect 14 -6461 66 -6401
rect 66 -6461 71 -6401
rect 331 -6461 391 -6401
rect 467 -6111 527 -6051
rect 787 -6111 847 -6051
rect 923 -6111 983 -6051
rect 1243 -6111 1303 -6051
rect 1381 -6111 1441 -6051
rect 1701 -6111 1761 -6051
rect 1837 -6111 1897 -6051
rect 2157 -6111 2217 -6051
rect 2293 -6111 2353 -6051
rect 2613 -6111 2673 -6051
rect 2751 -6111 2811 -6051
rect 3071 -6111 3131 -6051
rect 3207 -6111 3267 -6051
rect 3527 -6111 3587 -6051
rect 3663 -6111 3723 -6051
rect 3983 -6111 4043 -6051
rect 4121 -6111 4181 -6051
rect 4441 -6111 4501 -6051
rect 4577 -6111 4637 -6051
rect 4897 -6111 4957 -6051
rect 5033 -6111 5093 -6051
rect 5353 -6111 5413 -6051
rect 5491 -6111 5551 -6051
rect 5811 -6111 5871 -6051
rect 5947 -6111 6007 -6051
rect 6267 -6111 6327 -6051
rect 6403 -6111 6463 -6051
rect 6723 -6111 6783 -6051
rect 6861 -6111 6921 -6051
rect 7181 -6111 7241 -6051
rect 7317 -6111 7377 -6051
rect 7637 -6111 7697 -6051
rect 7773 -6111 7833 -6051
rect 8093 -6111 8153 -6051
rect 8247 -6111 8307 -6051
rect 8567 -6111 8627 -6051
rect 8703 -6111 8763 -6051
rect 9023 -6111 9083 -6051
rect 9161 -6111 9221 -6051
rect 9481 -6111 9541 -6051
rect 9617 -6111 9677 -6051
rect 9937 -6111 9997 -6051
rect 10073 -6111 10133 -6051
rect 10393 -6111 10453 -6051
rect 10531 -6111 10591 -6051
rect 10851 -6111 10911 -6051
rect 10987 -6111 11047 -6051
rect 11307 -6111 11367 -6051
rect 11443 -6111 11503 -6051
rect 11763 -6111 11823 -6051
rect 11901 -6111 11961 -6051
rect 12221 -6111 12281 -6051
rect 12357 -6111 12417 -6051
rect 12677 -6111 12737 -6051
rect 12813 -6111 12873 -6051
rect 13133 -6111 13193 -6051
rect 13271 -6111 13331 -6051
rect 13591 -6111 13651 -6051
rect 13727 -6111 13787 -6051
rect 14047 -6111 14107 -6051
rect 14183 -6111 14243 -6051
rect 14503 -6111 14563 -6051
rect 14641 -6111 14701 -6051
rect 14961 -6111 15021 -6051
rect 15097 -6111 15157 -6051
rect 15417 -6111 15477 -6051
rect 467 -6461 527 -6401
rect 787 -6461 847 -6401
rect 923 -6461 983 -6401
rect 1243 -6461 1303 -6401
rect 1381 -6461 1441 -6401
rect 1701 -6461 1761 -6401
rect 1837 -6461 1897 -6401
rect 2157 -6461 2217 -6401
rect 2293 -6461 2353 -6401
rect 2613 -6461 2673 -6401
rect 2751 -6461 2811 -6401
rect 3071 -6461 3131 -6401
rect 3207 -6461 3267 -6401
rect 3527 -6461 3587 -6401
rect 3663 -6461 3723 -6401
rect 3983 -6461 4043 -6401
rect 4121 -6461 4181 -6401
rect 4441 -6461 4501 -6401
rect 4577 -6461 4637 -6401
rect 4897 -6461 4957 -6401
rect 5033 -6461 5093 -6401
rect 5353 -6461 5413 -6401
rect 5491 -6461 5551 -6401
rect 5811 -6461 5871 -6401
rect 5947 -6461 6007 -6401
rect 6267 -6461 6327 -6401
rect 6403 -6461 6463 -6401
rect 6723 -6461 6783 -6401
rect 6861 -6461 6921 -6401
rect 7181 -6461 7241 -6401
rect 7317 -6461 7377 -6401
rect 7637 -6461 7697 -6401
rect 7773 -6461 7833 -6401
rect 8093 -6461 8153 -6401
rect 8247 -6461 8307 -6401
rect 8567 -6461 8627 -6401
rect 8703 -6461 8763 -6401
rect 9023 -6461 9083 -6401
rect 9161 -6461 9221 -6401
rect 9481 -6461 9541 -6401
rect 9617 -6461 9677 -6401
rect 9937 -6461 9997 -6401
rect 10073 -6461 10133 -6401
rect 10393 -6461 10453 -6401
rect 10531 -6461 10591 -6401
rect 10851 -6461 10911 -6401
rect 10987 -6461 11047 -6401
rect 11307 -6461 11367 -6401
rect 11443 -6461 11503 -6401
rect 11763 -6461 11823 -6401
rect 11901 -6461 11961 -6401
rect 12221 -6461 12281 -6401
rect 12357 -6461 12417 -6401
rect 12677 -6461 12737 -6401
rect 12813 -6461 12873 -6401
rect 13133 -6461 13193 -6401
rect 13271 -6461 13331 -6401
rect 13591 -6461 13651 -6401
rect 13727 -6461 13787 -6401
rect 14047 -6461 14107 -6401
rect 14183 -6461 14243 -6401
rect 14503 -6461 14563 -6401
rect 14641 -6461 14701 -6401
rect 14961 -6461 15021 -6401
rect 15097 -6461 15157 -6401
rect 15417 -6461 15477 -6401
rect 11 -6603 14 -6543
rect 14 -6603 66 -6543
rect 66 -6603 71 -6543
rect 331 -6603 391 -6543
rect 11 -6953 14 -6893
rect 14 -6953 66 -6893
rect 66 -6953 71 -6893
rect 331 -6953 391 -6893
rect 467 -6603 527 -6543
rect 787 -6603 847 -6543
rect 923 -6603 983 -6543
rect 1243 -6603 1303 -6543
rect 1381 -6603 1441 -6543
rect 1701 -6603 1761 -6543
rect 1837 -6603 1897 -6543
rect 2157 -6603 2217 -6543
rect 2293 -6603 2353 -6543
rect 2613 -6603 2673 -6543
rect 2751 -6603 2811 -6543
rect 3071 -6603 3131 -6543
rect 3207 -6603 3267 -6543
rect 3527 -6603 3587 -6543
rect 3663 -6603 3723 -6543
rect 3983 -6603 4043 -6543
rect 4121 -6603 4181 -6543
rect 4441 -6603 4501 -6543
rect 4577 -6603 4637 -6543
rect 4897 -6603 4957 -6543
rect 5033 -6603 5093 -6543
rect 5353 -6603 5413 -6543
rect 5491 -6603 5551 -6543
rect 5811 -6603 5871 -6543
rect 5947 -6603 6007 -6543
rect 6267 -6603 6327 -6543
rect 6403 -6603 6463 -6543
rect 6723 -6603 6783 -6543
rect 6861 -6603 6921 -6543
rect 7181 -6603 7241 -6543
rect 7317 -6603 7377 -6543
rect 7637 -6603 7697 -6543
rect 7773 -6603 7833 -6543
rect 8093 -6603 8153 -6543
rect 8247 -6603 8307 -6543
rect 8567 -6603 8627 -6543
rect 8703 -6603 8763 -6543
rect 9023 -6603 9083 -6543
rect 9161 -6603 9221 -6543
rect 9481 -6603 9541 -6543
rect 9617 -6603 9677 -6543
rect 9937 -6603 9997 -6543
rect 10073 -6603 10133 -6543
rect 10393 -6603 10453 -6543
rect 10531 -6603 10591 -6543
rect 10851 -6603 10911 -6543
rect 10987 -6603 11047 -6543
rect 11307 -6603 11367 -6543
rect 11443 -6603 11503 -6543
rect 11763 -6603 11823 -6543
rect 11901 -6603 11961 -6543
rect 12221 -6603 12281 -6543
rect 12357 -6603 12417 -6543
rect 12677 -6603 12737 -6543
rect 12813 -6603 12873 -6543
rect 13133 -6603 13193 -6543
rect 13271 -6603 13331 -6543
rect 13591 -6603 13651 -6543
rect 13727 -6603 13787 -6543
rect 14047 -6603 14107 -6543
rect 14183 -6603 14243 -6543
rect 14503 -6603 14563 -6543
rect 14641 -6603 14701 -6543
rect 14961 -6603 15021 -6543
rect 15097 -6603 15157 -6543
rect 15417 -6603 15477 -6543
rect 467 -6953 527 -6893
rect 787 -6953 847 -6893
rect 923 -6953 983 -6893
rect 1243 -6953 1303 -6893
rect 1381 -6953 1441 -6893
rect 1701 -6953 1761 -6893
rect 1837 -6953 1897 -6893
rect 2157 -6953 2217 -6893
rect 2293 -6953 2353 -6893
rect 2613 -6953 2673 -6893
rect 2751 -6953 2811 -6893
rect 3071 -6953 3131 -6893
rect 3207 -6953 3267 -6893
rect 3527 -6953 3587 -6893
rect 3663 -6953 3723 -6893
rect 3983 -6953 4043 -6893
rect 4121 -6953 4181 -6893
rect 4441 -6953 4501 -6893
rect 4577 -6953 4637 -6893
rect 4897 -6953 4957 -6893
rect 5033 -6953 5093 -6893
rect 5353 -6953 5413 -6893
rect 5491 -6953 5551 -6893
rect 5811 -6953 5871 -6893
rect 5947 -6953 6007 -6893
rect 6267 -6953 6327 -6893
rect 6403 -6953 6463 -6893
rect 6723 -6953 6783 -6893
rect 6861 -6953 6921 -6893
rect 7181 -6953 7241 -6893
rect 7317 -6953 7377 -6893
rect 7637 -6953 7697 -6893
rect 7773 -6953 7833 -6893
rect 8093 -6953 8153 -6893
rect 8247 -6953 8307 -6893
rect 8567 -6953 8627 -6893
rect 8703 -6953 8763 -6893
rect 9023 -6953 9083 -6893
rect 9161 -6953 9221 -6893
rect 9481 -6953 9541 -6893
rect 9617 -6953 9677 -6893
rect 9937 -6953 9997 -6893
rect 10073 -6953 10133 -6893
rect 10393 -6953 10453 -6893
rect 10531 -6953 10591 -6893
rect 10851 -6953 10911 -6893
rect 10987 -6953 11047 -6893
rect 11307 -6953 11367 -6893
rect 11443 -6953 11503 -6893
rect 11763 -6953 11823 -6893
rect 11901 -6953 11961 -6893
rect 12221 -6953 12281 -6893
rect 12357 -6953 12417 -6893
rect 12677 -6953 12737 -6893
rect 12813 -6953 12873 -6893
rect 13133 -6953 13193 -6893
rect 13271 -6953 13331 -6893
rect 13591 -6953 13651 -6893
rect 13727 -6953 13787 -6893
rect 14047 -6953 14107 -6893
rect 14183 -6953 14243 -6893
rect 14503 -6953 14563 -6893
rect 14641 -6953 14701 -6893
rect 14961 -6953 15021 -6893
rect 15097 -6953 15157 -6893
rect 15417 -6953 15477 -6893
rect 11 -7119 14 -7059
rect 14 -7119 66 -7059
rect 66 -7119 71 -7059
rect 331 -7119 391 -7059
rect 11 -7469 14 -7409
rect 14 -7469 66 -7409
rect 66 -7469 71 -7409
rect 331 -7469 391 -7409
rect 467 -7119 527 -7059
rect 787 -7119 847 -7059
rect 923 -7119 983 -7059
rect 1243 -7119 1303 -7059
rect 1381 -7119 1441 -7059
rect 1701 -7119 1761 -7059
rect 1837 -7119 1897 -7059
rect 2157 -7119 2217 -7059
rect 2293 -7119 2353 -7059
rect 2613 -7119 2673 -7059
rect 2751 -7119 2811 -7059
rect 3071 -7119 3131 -7059
rect 3207 -7119 3267 -7059
rect 3527 -7119 3587 -7059
rect 3663 -7119 3723 -7059
rect 3983 -7119 4043 -7059
rect 467 -7469 527 -7409
rect 787 -7469 847 -7409
rect 923 -7469 983 -7409
rect 1243 -7469 1303 -7409
rect 1381 -7469 1441 -7409
rect 1701 -7469 1761 -7409
rect 1837 -7469 1897 -7409
rect 2157 -7469 2217 -7409
rect 2293 -7469 2353 -7409
rect 2613 -7469 2673 -7409
rect 2751 -7469 2811 -7409
rect 3071 -7469 3131 -7409
rect 3207 -7469 3267 -7409
rect 3527 -7469 3587 -7409
rect 3663 -7469 3723 -7409
rect 3983 -7469 4043 -7409
rect 4121 -7119 4181 -7059
rect 4441 -7119 4501 -7059
rect 4577 -7119 4637 -7059
rect 4897 -7119 4957 -7059
rect 5033 -7119 5093 -7059
rect 5353 -7119 5413 -7059
rect 5491 -7119 5551 -7059
rect 5811 -7119 5871 -7059
rect 5947 -7119 6007 -7059
rect 6267 -7119 6327 -7059
rect 6403 -7119 6463 -7059
rect 6723 -7119 6783 -7059
rect 6861 -7119 6921 -7059
rect 7181 -7119 7241 -7059
rect 7317 -7119 7377 -7059
rect 7637 -7119 7697 -7059
rect 7773 -7119 7833 -7059
rect 8093 -7119 8153 -7059
rect 8247 -7119 8307 -7059
rect 8567 -7119 8627 -7059
rect 8703 -7119 8763 -7059
rect 9023 -7119 9083 -7059
rect 9161 -7119 9221 -7059
rect 9481 -7119 9541 -7059
rect 9617 -7119 9677 -7059
rect 9937 -7119 9997 -7059
rect 10073 -7119 10133 -7059
rect 10393 -7119 10453 -7059
rect 10531 -7119 10591 -7059
rect 10851 -7119 10911 -7059
rect 10987 -7119 11047 -7059
rect 11307 -7119 11367 -7059
rect 11443 -7119 11503 -7059
rect 11763 -7119 11823 -7059
rect 11901 -7119 11961 -7059
rect 12221 -7119 12281 -7059
rect 12357 -7119 12417 -7059
rect 12677 -7119 12737 -7059
rect 12813 -7119 12873 -7059
rect 13133 -7119 13193 -7059
rect 13271 -7119 13331 -7059
rect 13591 -7119 13651 -7059
rect 13727 -7119 13787 -7059
rect 14047 -7119 14107 -7059
rect 14183 -7119 14243 -7059
rect 14503 -7119 14563 -7059
rect 14641 -7119 14701 -7059
rect 14961 -7119 15021 -7059
rect 15097 -7119 15157 -7059
rect 15417 -7119 15477 -7059
rect 4121 -7469 4181 -7409
rect 4441 -7469 4501 -7409
rect 4577 -7469 4637 -7409
rect 4897 -7469 4957 -7409
rect 5033 -7469 5093 -7409
rect 5353 -7469 5413 -7409
rect 5491 -7469 5551 -7409
rect 5811 -7469 5871 -7409
rect 5947 -7469 6007 -7409
rect 6267 -7469 6327 -7409
rect 6403 -7469 6463 -7409
rect 6723 -7469 6783 -7409
rect 6861 -7469 6921 -7409
rect 7181 -7469 7241 -7409
rect 7317 -7469 7377 -7409
rect 7637 -7469 7697 -7409
rect 7773 -7469 7833 -7409
rect 8093 -7469 8153 -7409
rect 8247 -7469 8307 -7409
rect 8567 -7469 8627 -7409
rect 8703 -7469 8763 -7409
rect 9023 -7469 9083 -7409
rect 9161 -7469 9221 -7409
rect 9481 -7469 9541 -7409
rect 9617 -7469 9677 -7409
rect 9937 -7469 9997 -7409
rect 10073 -7469 10133 -7409
rect 10393 -7469 10453 -7409
rect 10531 -7469 10591 -7409
rect 10851 -7469 10911 -7409
rect 10987 -7469 11047 -7409
rect 11307 -7469 11367 -7409
rect 11443 -7469 11503 -7409
rect 11763 -7469 11823 -7409
rect 11901 -7469 11961 -7409
rect 12221 -7469 12281 -7409
rect 12357 -7469 12417 -7409
rect 12677 -7469 12737 -7409
rect 12813 -7469 12873 -7409
rect 13133 -7469 13193 -7409
rect 13271 -7469 13331 -7409
rect 13591 -7469 13651 -7409
rect 13727 -7469 13787 -7409
rect 14047 -7469 14107 -7409
rect 14183 -7469 14243 -7409
rect 14503 -7469 14563 -7409
rect 14641 -7469 14701 -7409
rect 14961 -7469 15021 -7409
rect 15097 -7469 15157 -7409
rect 15417 -7469 15477 -7409
rect 11 -7621 14 -7561
rect 14 -7621 66 -7561
rect 66 -7621 71 -7561
rect 331 -7621 391 -7561
rect 11 -7971 14 -7911
rect 14 -7971 66 -7911
rect 66 -7971 71 -7911
rect 331 -7971 391 -7911
rect 467 -7621 527 -7561
rect 787 -7621 847 -7561
rect 923 -7621 983 -7561
rect 1243 -7621 1303 -7561
rect 1381 -7621 1441 -7561
rect 1701 -7621 1761 -7561
rect 1837 -7621 1897 -7561
rect 2157 -7621 2217 -7561
rect 2293 -7621 2353 -7561
rect 2613 -7621 2673 -7561
rect 2751 -7621 2811 -7561
rect 3071 -7621 3131 -7561
rect 3207 -7621 3267 -7561
rect 3527 -7621 3587 -7561
rect 3663 -7621 3723 -7561
rect 3983 -7621 4043 -7561
rect 467 -7971 527 -7911
rect 787 -7971 847 -7911
rect 923 -7971 983 -7911
rect 1243 -7971 1303 -7911
rect 1381 -7971 1441 -7911
rect 1701 -7971 1761 -7911
rect 1837 -7971 1897 -7911
rect 2157 -7971 2217 -7911
rect 2293 -7971 2353 -7911
rect 2613 -7971 2673 -7911
rect 2751 -7971 2811 -7911
rect 3071 -7971 3131 -7911
rect 3207 -7971 3267 -7911
rect 3527 -7971 3587 -7911
rect 3663 -7971 3723 -7911
rect 3983 -7971 4043 -7911
rect 4121 -7621 4181 -7561
rect 4441 -7621 4501 -7561
rect 4577 -7621 4637 -7561
rect 4897 -7621 4957 -7561
rect 5033 -7621 5093 -7561
rect 5353 -7621 5413 -7561
rect 5491 -7621 5551 -7561
rect 5811 -7621 5871 -7561
rect 5947 -7621 6007 -7561
rect 6267 -7621 6327 -7561
rect 6403 -7621 6463 -7561
rect 6723 -7621 6783 -7561
rect 6861 -7621 6921 -7561
rect 7181 -7621 7241 -7561
rect 7317 -7621 7377 -7561
rect 7637 -7621 7697 -7561
rect 7773 -7621 7833 -7561
rect 8093 -7621 8153 -7561
rect 8247 -7621 8307 -7561
rect 8567 -7621 8627 -7561
rect 8703 -7621 8763 -7561
rect 9023 -7621 9083 -7561
rect 9161 -7621 9221 -7561
rect 9481 -7621 9541 -7561
rect 9617 -7621 9677 -7561
rect 9937 -7621 9997 -7561
rect 10073 -7621 10133 -7561
rect 10393 -7621 10453 -7561
rect 10531 -7621 10591 -7561
rect 10851 -7621 10911 -7561
rect 10987 -7621 11047 -7561
rect 11307 -7621 11367 -7561
rect 11443 -7621 11503 -7561
rect 11763 -7621 11823 -7561
rect 11901 -7621 11961 -7561
rect 12221 -7621 12281 -7561
rect 12357 -7621 12417 -7561
rect 12677 -7621 12737 -7561
rect 12813 -7621 12873 -7561
rect 13133 -7621 13193 -7561
rect 13271 -7621 13331 -7561
rect 13591 -7621 13651 -7561
rect 13727 -7621 13787 -7561
rect 14047 -7621 14107 -7561
rect 14183 -7621 14243 -7561
rect 14503 -7621 14563 -7561
rect 14641 -7621 14701 -7561
rect 14961 -7621 15021 -7561
rect 15097 -7621 15157 -7561
rect 15417 -7621 15477 -7561
rect 4121 -7971 4181 -7911
rect 4441 -7971 4501 -7911
rect 4577 -7971 4637 -7911
rect 4897 -7971 4957 -7911
rect 5033 -7971 5093 -7911
rect 5353 -7971 5413 -7911
rect 5491 -7971 5551 -7911
rect 5811 -7971 5871 -7911
rect 5947 -7971 6007 -7911
rect 6267 -7971 6327 -7911
rect 6403 -7971 6463 -7911
rect 6723 -7971 6783 -7911
rect 6861 -7971 6921 -7911
rect 7181 -7971 7241 -7911
rect 7317 -7971 7377 -7911
rect 7637 -7971 7697 -7911
rect 7773 -7971 7833 -7911
rect 8093 -7971 8153 -7911
rect 8247 -7971 8307 -7911
rect 8567 -7971 8627 -7911
rect 8703 -7971 8763 -7911
rect 9023 -7971 9083 -7911
rect 9161 -7971 9221 -7911
rect 9481 -7971 9541 -7911
rect 9617 -7971 9677 -7911
rect 9937 -7971 9997 -7911
rect 10073 -7971 10133 -7911
rect 10393 -7971 10453 -7911
rect 10531 -7971 10591 -7911
rect 10851 -7971 10911 -7911
rect 10987 -7971 11047 -7911
rect 11307 -7971 11367 -7911
rect 11443 -7971 11503 -7911
rect 11763 -7971 11823 -7911
rect 11901 -7971 11961 -7911
rect 12221 -7971 12281 -7911
rect 12357 -7971 12417 -7911
rect 12677 -7971 12737 -7911
rect 12813 -7971 12873 -7911
rect 13133 -7971 13193 -7911
rect 13271 -7971 13331 -7911
rect 13591 -7971 13651 -7911
rect 13727 -7971 13787 -7911
rect 14047 -7971 14107 -7911
rect 14183 -7971 14243 -7911
rect 14503 -7971 14563 -7911
rect 14641 -7971 14701 -7911
rect 14961 -7971 15021 -7911
rect 15097 -7971 15157 -7911
rect 15417 -7971 15477 -7911
rect 11 -8113 14 -8053
rect 14 -8113 66 -8053
rect 66 -8113 71 -8053
rect 331 -8113 391 -8053
rect 11 -8463 14 -8403
rect 14 -8463 66 -8403
rect 66 -8463 71 -8403
rect 331 -8463 391 -8403
rect 467 -8113 527 -8053
rect 787 -8113 847 -8053
rect 923 -8113 983 -8053
rect 1243 -8113 1303 -8053
rect 1381 -8113 1441 -8053
rect 1701 -8113 1761 -8053
rect 1837 -8113 1897 -8053
rect 2157 -8113 2217 -8053
rect 2293 -8113 2353 -8053
rect 2613 -8113 2673 -8053
rect 2751 -8113 2811 -8053
rect 3071 -8113 3131 -8053
rect 3207 -8113 3267 -8053
rect 3527 -8113 3587 -8053
rect 3663 -8113 3723 -8053
rect 3983 -8113 4043 -8053
rect 467 -8463 527 -8403
rect 787 -8463 847 -8403
rect 923 -8463 983 -8403
rect 1243 -8463 1303 -8403
rect 1381 -8463 1441 -8403
rect 1701 -8463 1761 -8403
rect 1837 -8463 1897 -8403
rect 2157 -8463 2217 -8403
rect 2293 -8463 2353 -8403
rect 2613 -8463 2673 -8403
rect 2751 -8463 2811 -8403
rect 3071 -8463 3131 -8403
rect 3207 -8463 3267 -8403
rect 3527 -8463 3587 -8403
rect 3663 -8463 3723 -8403
rect 3983 -8463 4043 -8403
rect 4121 -8113 4181 -8053
rect 4441 -8113 4501 -8053
rect 4577 -8113 4637 -8053
rect 4897 -8113 4957 -8053
rect 5033 -8113 5093 -8053
rect 5353 -8113 5413 -8053
rect 5491 -8113 5551 -8053
rect 5811 -8113 5871 -8053
rect 5947 -8113 6007 -8053
rect 6267 -8113 6327 -8053
rect 6403 -8113 6463 -8053
rect 6723 -8113 6783 -8053
rect 6861 -8113 6921 -8053
rect 7181 -8113 7241 -8053
rect 7317 -8113 7377 -8053
rect 7637 -8113 7697 -8053
rect 7773 -8113 7833 -8053
rect 8093 -8113 8153 -8053
rect 8247 -8113 8307 -8053
rect 8567 -8113 8627 -8053
rect 8703 -8113 8763 -8053
rect 9023 -8113 9083 -8053
rect 9161 -8113 9221 -8053
rect 9481 -8113 9541 -8053
rect 9617 -8113 9677 -8053
rect 9937 -8113 9997 -8053
rect 10073 -8113 10133 -8053
rect 10393 -8113 10453 -8053
rect 10531 -8113 10591 -8053
rect 10851 -8113 10911 -8053
rect 10987 -8113 11047 -8053
rect 11307 -8113 11367 -8053
rect 11443 -8113 11503 -8053
rect 11763 -8113 11823 -8053
rect 11901 -8113 11961 -8053
rect 12221 -8113 12281 -8053
rect 12357 -8113 12417 -8053
rect 12677 -8113 12737 -8053
rect 12813 -8113 12873 -8053
rect 13133 -8113 13193 -8053
rect 13271 -8113 13331 -8053
rect 13591 -8113 13651 -8053
rect 13727 -8113 13787 -8053
rect 14047 -8113 14107 -8053
rect 14183 -8113 14243 -8053
rect 14503 -8113 14563 -8053
rect 14641 -8113 14701 -8053
rect 14961 -8113 15021 -8053
rect 15097 -8113 15157 -8053
rect 15417 -8113 15477 -8053
rect 4121 -8463 4181 -8403
rect 4441 -8463 4501 -8403
rect 4577 -8463 4637 -8403
rect 4897 -8463 4957 -8403
rect 5033 -8463 5093 -8403
rect 5353 -8463 5413 -8403
rect 5491 -8463 5551 -8403
rect 5811 -8463 5871 -8403
rect 5947 -8463 6007 -8403
rect 6267 -8463 6327 -8403
rect 6403 -8463 6463 -8403
rect 6723 -8463 6783 -8403
rect 6861 -8463 6921 -8403
rect 7181 -8463 7241 -8403
rect 7317 -8463 7377 -8403
rect 7637 -8463 7697 -8403
rect 7773 -8463 7833 -8403
rect 8093 -8463 8153 -8403
rect 8247 -8463 8307 -8403
rect 8567 -8463 8627 -8403
rect 8703 -8463 8763 -8403
rect 9023 -8463 9083 -8403
rect 9161 -8463 9221 -8403
rect 9481 -8463 9541 -8403
rect 9617 -8463 9677 -8403
rect 9937 -8463 9997 -8403
rect 10073 -8463 10133 -8403
rect 10393 -8463 10453 -8403
rect 10531 -8463 10591 -8403
rect 10851 -8463 10911 -8403
rect 10987 -8463 11047 -8403
rect 11307 -8463 11367 -8403
rect 11443 -8463 11503 -8403
rect 11763 -8463 11823 -8403
rect 11901 -8463 11961 -8403
rect 12221 -8463 12281 -8403
rect 12357 -8463 12417 -8403
rect 12677 -8463 12737 -8403
rect 12813 -8463 12873 -8403
rect 13133 -8463 13193 -8403
rect 13271 -8463 13331 -8403
rect 13591 -8463 13651 -8403
rect 13727 -8463 13787 -8403
rect 14047 -8463 14107 -8403
rect 14183 -8463 14243 -8403
rect 14503 -8463 14563 -8403
rect 14641 -8463 14701 -8403
rect 14961 -8463 15021 -8403
rect 15097 -8463 15157 -8403
rect 15417 -8463 15477 -8403
rect 11 -8607 14 -8547
rect 14 -8607 66 -8547
rect 66 -8607 71 -8547
rect 331 -8607 391 -8547
rect 11 -8957 14 -8897
rect 14 -8957 66 -8897
rect 66 -8957 71 -8897
rect 331 -8957 391 -8897
rect 467 -8607 527 -8547
rect 787 -8607 847 -8547
rect 923 -8607 983 -8547
rect 1243 -8607 1303 -8547
rect 1381 -8607 1441 -8547
rect 1701 -8607 1761 -8547
rect 1837 -8607 1897 -8547
rect 2157 -8607 2217 -8547
rect 2293 -8607 2353 -8547
rect 2613 -8607 2673 -8547
rect 2751 -8607 2811 -8547
rect 3071 -8607 3131 -8547
rect 3207 -8607 3267 -8547
rect 3527 -8607 3587 -8547
rect 3663 -8607 3723 -8547
rect 3983 -8607 4043 -8547
rect 467 -8957 527 -8897
rect 787 -8957 847 -8897
rect 923 -8957 983 -8897
rect 1243 -8957 1303 -8897
rect 1381 -8957 1441 -8897
rect 1701 -8957 1761 -8897
rect 1837 -8957 1897 -8897
rect 2157 -8957 2217 -8897
rect 2293 -8957 2353 -8897
rect 2613 -8957 2673 -8897
rect 2751 -8957 2811 -8897
rect 3071 -8957 3131 -8897
rect 3207 -8957 3267 -8897
rect 3527 -8957 3587 -8897
rect 3663 -8957 3723 -8897
rect 3983 -8957 4043 -8897
rect 4121 -8607 4181 -8547
rect 4441 -8607 4501 -8547
rect 4577 -8607 4637 -8547
rect 4897 -8607 4957 -8547
rect 5033 -8607 5093 -8547
rect 5353 -8607 5413 -8547
rect 5491 -8607 5551 -8547
rect 5811 -8607 5871 -8547
rect 5947 -8607 6007 -8547
rect 6267 -8607 6327 -8547
rect 6403 -8607 6463 -8547
rect 6723 -8607 6783 -8547
rect 6861 -8607 6921 -8547
rect 7181 -8607 7241 -8547
rect 4121 -8957 4181 -8897
rect 4441 -8957 4501 -8897
rect 4577 -8957 4637 -8897
rect 4897 -8957 4957 -8897
rect 5033 -8957 5093 -8897
rect 5353 -8957 5413 -8897
rect 5491 -8957 5551 -8897
rect 5811 -8957 5871 -8897
rect 5947 -8957 6007 -8897
rect 6267 -8957 6327 -8897
rect 6403 -8957 6463 -8897
rect 6723 -8957 6783 -8897
rect 6861 -8957 6921 -8897
rect 7181 -8957 7241 -8897
rect 7317 -8607 7377 -8547
rect 7637 -8607 7697 -8547
rect 7773 -8607 7833 -8547
rect 8093 -8607 8153 -8547
rect 8247 -8607 8307 -8547
rect 8567 -8607 8627 -8547
rect 8703 -8607 8763 -8547
rect 9023 -8607 9083 -8547
rect 9161 -8607 9221 -8547
rect 9481 -8607 9541 -8547
rect 9617 -8607 9677 -8547
rect 9937 -8607 9997 -8547
rect 10073 -8607 10133 -8547
rect 10393 -8607 10453 -8547
rect 10531 -8607 10591 -8547
rect 10851 -8607 10911 -8547
rect 10987 -8607 11047 -8547
rect 11307 -8607 11367 -8547
rect 11443 -8607 11503 -8547
rect 11763 -8607 11823 -8547
rect 11901 -8607 11961 -8547
rect 12221 -8607 12281 -8547
rect 12357 -8607 12417 -8547
rect 12677 -8607 12737 -8547
rect 12813 -8607 12873 -8547
rect 13133 -8607 13193 -8547
rect 13271 -8607 13331 -8547
rect 13591 -8607 13651 -8547
rect 13727 -8607 13787 -8547
rect 14047 -8607 14107 -8547
rect 14183 -8607 14243 -8547
rect 14503 -8607 14563 -8547
rect 14641 -8607 14701 -8547
rect 14961 -8607 15021 -8547
rect 15097 -8607 15157 -8547
rect 15417 -8607 15477 -8547
rect 7317 -8957 7377 -8897
rect 7637 -8957 7697 -8897
rect 7773 -8957 7833 -8897
rect 8093 -8957 8153 -8897
rect 8247 -8957 8307 -8897
rect 8567 -8957 8627 -8897
rect 8703 -8957 8763 -8897
rect 9023 -8957 9083 -8897
rect 9161 -8957 9221 -8897
rect 9481 -8957 9541 -8897
rect 9617 -8957 9677 -8897
rect 9937 -8957 9997 -8897
rect 10073 -8957 10133 -8897
rect 10393 -8957 10453 -8897
rect 10531 -8957 10591 -8897
rect 10851 -8957 10911 -8897
rect 10987 -8957 11047 -8897
rect 11307 -8957 11367 -8897
rect 11443 -8957 11503 -8897
rect 11763 -8957 11823 -8897
rect 11901 -8957 11961 -8897
rect 12221 -8957 12281 -8897
rect 12357 -8957 12417 -8897
rect 12677 -8957 12737 -8897
rect 12813 -8957 12873 -8897
rect 13133 -8957 13193 -8897
rect 13271 -8957 13331 -8897
rect 13591 -8957 13651 -8897
rect 13727 -8957 13787 -8897
rect 14047 -8957 14107 -8897
rect 14183 -8957 14243 -8897
rect 14503 -8957 14563 -8897
rect 14641 -8957 14701 -8897
rect 14961 -8957 15021 -8897
rect 15097 -8957 15157 -8897
rect 15417 -8957 15477 -8897
rect 11 -9109 14 -9049
rect 14 -9109 66 -9049
rect 66 -9109 71 -9049
rect 331 -9109 391 -9049
rect 11 -9459 14 -9399
rect 14 -9459 66 -9399
rect 66 -9459 71 -9399
rect 331 -9459 391 -9399
rect 467 -9109 527 -9049
rect 787 -9109 847 -9049
rect 923 -9109 983 -9049
rect 1243 -9109 1303 -9049
rect 1381 -9109 1441 -9049
rect 1701 -9109 1761 -9049
rect 1837 -9109 1897 -9049
rect 2157 -9109 2217 -9049
rect 2293 -9109 2353 -9049
rect 2613 -9109 2673 -9049
rect 2751 -9109 2811 -9049
rect 3071 -9109 3131 -9049
rect 3207 -9109 3267 -9049
rect 3527 -9109 3587 -9049
rect 3663 -9109 3723 -9049
rect 3983 -9109 4043 -9049
rect 467 -9459 527 -9399
rect 787 -9459 847 -9399
rect 923 -9459 983 -9399
rect 1243 -9459 1303 -9399
rect 1381 -9459 1441 -9399
rect 1701 -9459 1761 -9399
rect 1837 -9459 1897 -9399
rect 2157 -9459 2217 -9399
rect 2293 -9459 2353 -9399
rect 2613 -9459 2673 -9399
rect 2751 -9459 2811 -9399
rect 3071 -9459 3131 -9399
rect 3207 -9459 3267 -9399
rect 3527 -9459 3587 -9399
rect 3663 -9459 3723 -9399
rect 3983 -9459 4043 -9399
rect 4121 -9109 4181 -9049
rect 4441 -9109 4501 -9049
rect 4577 -9109 4637 -9049
rect 4897 -9109 4957 -9049
rect 5033 -9109 5093 -9049
rect 5353 -9109 5413 -9049
rect 5491 -9109 5551 -9049
rect 5811 -9109 5871 -9049
rect 5947 -9109 6007 -9049
rect 6267 -9109 6327 -9049
rect 6403 -9109 6463 -9049
rect 6723 -9109 6783 -9049
rect 6861 -9109 6921 -9049
rect 7181 -9109 7241 -9049
rect 4121 -9459 4181 -9399
rect 4441 -9459 4501 -9399
rect 4577 -9459 4637 -9399
rect 4897 -9459 4957 -9399
rect 5033 -9459 5093 -9399
rect 5353 -9459 5413 -9399
rect 5491 -9459 5551 -9399
rect 5811 -9459 5871 -9399
rect 5947 -9459 6007 -9399
rect 6267 -9459 6327 -9399
rect 6403 -9459 6463 -9399
rect 6723 -9459 6783 -9399
rect 6861 -9459 6921 -9399
rect 7181 -9459 7241 -9399
rect 7317 -9109 7377 -9049
rect 7637 -9109 7697 -9049
rect 7773 -9109 7833 -9049
rect 8093 -9109 8153 -9049
rect 8247 -9109 8307 -9049
rect 8567 -9109 8627 -9049
rect 8703 -9109 8763 -9049
rect 9023 -9109 9083 -9049
rect 9161 -9109 9221 -9049
rect 9481 -9109 9541 -9049
rect 9617 -9109 9677 -9049
rect 9937 -9109 9997 -9049
rect 10073 -9109 10133 -9049
rect 10393 -9109 10453 -9049
rect 10531 -9109 10591 -9049
rect 10851 -9109 10911 -9049
rect 10987 -9109 11047 -9049
rect 11307 -9109 11367 -9049
rect 11443 -9109 11503 -9049
rect 11763 -9109 11823 -9049
rect 11901 -9109 11961 -9049
rect 12221 -9109 12281 -9049
rect 12357 -9109 12417 -9049
rect 12677 -9109 12737 -9049
rect 12813 -9109 12873 -9049
rect 13133 -9109 13193 -9049
rect 13271 -9109 13331 -9049
rect 13591 -9109 13651 -9049
rect 13727 -9109 13787 -9049
rect 14047 -9109 14107 -9049
rect 14183 -9109 14243 -9049
rect 14503 -9109 14563 -9049
rect 14641 -9109 14701 -9049
rect 14961 -9109 15021 -9049
rect 15097 -9109 15157 -9049
rect 15417 -9109 15477 -9049
rect 7317 -9459 7377 -9399
rect 7637 -9459 7697 -9399
rect 7773 -9459 7833 -9399
rect 8093 -9459 8153 -9399
rect 8247 -9459 8307 -9399
rect 8567 -9459 8627 -9399
rect 8703 -9459 8763 -9399
rect 9023 -9459 9083 -9399
rect 9161 -9459 9221 -9399
rect 9481 -9459 9541 -9399
rect 9617 -9459 9677 -9399
rect 9937 -9459 9997 -9399
rect 10073 -9459 10133 -9399
rect 10393 -9459 10453 -9399
rect 10531 -9459 10591 -9399
rect 10851 -9459 10911 -9399
rect 10987 -9459 11047 -9399
rect 11307 -9459 11367 -9399
rect 11443 -9459 11503 -9399
rect 11763 -9459 11823 -9399
rect 11901 -9459 11961 -9399
rect 12221 -9459 12281 -9399
rect 12357 -9459 12417 -9399
rect 12677 -9459 12737 -9399
rect 12813 -9459 12873 -9399
rect 13133 -9459 13193 -9399
rect 13271 -9459 13331 -9399
rect 13591 -9459 13651 -9399
rect 13727 -9459 13787 -9399
rect 14047 -9459 14107 -9399
rect 14183 -9459 14243 -9399
rect 14503 -9459 14563 -9399
rect 14641 -9459 14701 -9399
rect 14961 -9459 15021 -9399
rect 15097 -9459 15157 -9399
rect 15417 -9459 15477 -9399
rect 11 -9601 14 -9541
rect 14 -9601 66 -9541
rect 66 -9601 71 -9541
rect 331 -9601 391 -9541
rect 11 -9951 14 -9891
rect 14 -9951 66 -9891
rect 66 -9951 71 -9891
rect 331 -9951 391 -9891
rect 467 -9601 527 -9541
rect 787 -9601 847 -9541
rect 923 -9601 983 -9541
rect 1243 -9601 1303 -9541
rect 1381 -9601 1441 -9541
rect 1701 -9601 1761 -9541
rect 1837 -9601 1897 -9541
rect 2157 -9601 2217 -9541
rect 2293 -9601 2353 -9541
rect 2613 -9601 2673 -9541
rect 2751 -9601 2811 -9541
rect 3071 -9601 3131 -9541
rect 3207 -9601 3267 -9541
rect 3527 -9601 3587 -9541
rect 3663 -9601 3723 -9541
rect 3983 -9601 4043 -9541
rect 467 -9951 527 -9891
rect 787 -9951 847 -9891
rect 923 -9951 983 -9891
rect 1243 -9951 1303 -9891
rect 1381 -9951 1441 -9891
rect 1701 -9951 1761 -9891
rect 1837 -9951 1897 -9891
rect 2157 -9951 2217 -9891
rect 2293 -9951 2353 -9891
rect 2613 -9951 2673 -9891
rect 2751 -9951 2811 -9891
rect 3071 -9951 3131 -9891
rect 3207 -9951 3267 -9891
rect 3527 -9951 3587 -9891
rect 3663 -9951 3723 -9891
rect 3983 -9951 4043 -9891
rect 4121 -9601 4181 -9541
rect 4441 -9601 4501 -9541
rect 4577 -9601 4637 -9541
rect 4897 -9601 4957 -9541
rect 5033 -9601 5093 -9541
rect 5353 -9601 5413 -9541
rect 5491 -9601 5551 -9541
rect 5811 -9601 5871 -9541
rect 5947 -9601 6007 -9541
rect 6267 -9601 6327 -9541
rect 6403 -9601 6463 -9541
rect 6723 -9601 6783 -9541
rect 6861 -9601 6921 -9541
rect 7181 -9601 7241 -9541
rect 4121 -9951 4181 -9891
rect 4441 -9951 4501 -9891
rect 4577 -9951 4637 -9891
rect 4897 -9951 4957 -9891
rect 5033 -9951 5093 -9891
rect 5353 -9951 5413 -9891
rect 5491 -9951 5551 -9891
rect 5811 -9951 5871 -9891
rect 5947 -9951 6007 -9891
rect 6267 -9951 6327 -9891
rect 6403 -9951 6463 -9891
rect 6723 -9951 6783 -9891
rect 6861 -9951 6921 -9891
rect 7181 -9951 7241 -9891
rect 7317 -9601 7377 -9541
rect 7637 -9601 7697 -9541
rect 7773 -9601 7833 -9541
rect 8093 -9601 8153 -9541
rect 8247 -9601 8307 -9541
rect 8567 -9601 8627 -9541
rect 8703 -9601 8763 -9541
rect 9023 -9601 9083 -9541
rect 9161 -9601 9221 -9541
rect 9481 -9601 9541 -9541
rect 9617 -9601 9677 -9541
rect 9937 -9601 9997 -9541
rect 10073 -9601 10133 -9541
rect 10393 -9601 10453 -9541
rect 10531 -9601 10591 -9541
rect 10851 -9601 10911 -9541
rect 10987 -9601 11047 -9541
rect 11307 -9601 11367 -9541
rect 11443 -9601 11503 -9541
rect 11763 -9601 11823 -9541
rect 11901 -9601 11961 -9541
rect 12221 -9601 12281 -9541
rect 12357 -9601 12417 -9541
rect 12677 -9601 12737 -9541
rect 12813 -9601 12873 -9541
rect 13133 -9601 13193 -9541
rect 13271 -9601 13331 -9541
rect 13591 -9601 13651 -9541
rect 13727 -9601 13787 -9541
rect 14047 -9601 14107 -9541
rect 14183 -9601 14243 -9541
rect 14503 -9601 14563 -9541
rect 14641 -9601 14701 -9541
rect 14961 -9601 15021 -9541
rect 15097 -9601 15157 -9541
rect 15417 -9601 15477 -9541
rect 7317 -9951 7377 -9891
rect 7637 -9951 7697 -9891
rect 7773 -9951 7833 -9891
rect 8093 -9951 8153 -9891
rect 8247 -9951 8307 -9891
rect 8567 -9951 8627 -9891
rect 8703 -9951 8763 -9891
rect 9023 -9951 9083 -9891
rect 9161 -9951 9221 -9891
rect 9481 -9951 9541 -9891
rect 9617 -9951 9677 -9891
rect 9937 -9951 9997 -9891
rect 10073 -9951 10133 -9891
rect 10393 -9951 10453 -9891
rect 10531 -9951 10591 -9891
rect 10851 -9951 10911 -9891
rect 10987 -9951 11047 -9891
rect 11307 -9951 11367 -9891
rect 11443 -9951 11503 -9891
rect 11763 -9951 11823 -9891
rect 11901 -9951 11961 -9891
rect 12221 -9951 12281 -9891
rect 12357 -9951 12417 -9891
rect 12677 -9951 12737 -9891
rect 12813 -9951 12873 -9891
rect 13133 -9951 13193 -9891
rect 13271 -9951 13331 -9891
rect 13591 -9951 13651 -9891
rect 13727 -9951 13787 -9891
rect 14047 -9951 14107 -9891
rect 14183 -9951 14243 -9891
rect 14503 -9951 14563 -9891
rect 14641 -9951 14701 -9891
rect 14961 -9951 15021 -9891
rect 15097 -9951 15157 -9891
rect 15417 -9951 15477 -9891
rect 11 -10117 14 -10057
rect 14 -10117 66 -10057
rect 66 -10117 71 -10057
rect 331 -10117 391 -10057
rect 11 -10467 14 -10407
rect 14 -10467 66 -10407
rect 66 -10467 71 -10407
rect 331 -10467 391 -10407
rect 467 -10117 527 -10057
rect 787 -10117 847 -10057
rect 923 -10117 983 -10057
rect 1243 -10117 1303 -10057
rect 1381 -10117 1441 -10057
rect 1701 -10117 1761 -10057
rect 1837 -10117 1897 -10057
rect 2157 -10117 2217 -10057
rect 2293 -10117 2353 -10057
rect 2613 -10117 2673 -10057
rect 2751 -10117 2811 -10057
rect 3071 -10117 3131 -10057
rect 3207 -10117 3267 -10057
rect 3527 -10117 3587 -10057
rect 3663 -10117 3723 -10057
rect 3983 -10117 4043 -10057
rect 467 -10467 527 -10407
rect 787 -10467 847 -10407
rect 923 -10467 983 -10407
rect 1243 -10467 1303 -10407
rect 1381 -10467 1441 -10407
rect 1701 -10467 1761 -10407
rect 1837 -10467 1897 -10407
rect 2157 -10467 2217 -10407
rect 2293 -10467 2353 -10407
rect 2613 -10467 2673 -10407
rect 2751 -10467 2811 -10407
rect 3071 -10467 3131 -10407
rect 3207 -10467 3267 -10407
rect 3527 -10467 3587 -10407
rect 3663 -10467 3723 -10407
rect 3983 -10467 4043 -10407
rect 4121 -10117 4181 -10057
rect 4441 -10117 4501 -10057
rect 4577 -10117 4637 -10057
rect 4897 -10117 4957 -10057
rect 5033 -10117 5093 -10057
rect 5353 -10117 5413 -10057
rect 5491 -10117 5551 -10057
rect 5811 -10117 5871 -10057
rect 5947 -10117 6007 -10057
rect 6267 -10117 6327 -10057
rect 6403 -10117 6463 -10057
rect 6723 -10117 6783 -10057
rect 6861 -10117 6921 -10057
rect 7181 -10117 7241 -10057
rect 4121 -10467 4181 -10407
rect 4441 -10467 4501 -10407
rect 4577 -10467 4637 -10407
rect 4897 -10467 4957 -10407
rect 5033 -10467 5093 -10407
rect 5353 -10467 5413 -10407
rect 5491 -10467 5551 -10407
rect 5811 -10467 5871 -10407
rect 5947 -10467 6007 -10407
rect 6267 -10467 6327 -10407
rect 6403 -10467 6463 -10407
rect 6723 -10467 6783 -10407
rect 6861 -10467 6921 -10407
rect 7181 -10467 7241 -10407
rect 7317 -10117 7377 -10057
rect 7637 -10117 7697 -10057
rect 7773 -10117 7833 -10057
rect 8093 -10117 8153 -10057
rect 8247 -10117 8307 -10057
rect 8567 -10117 8627 -10057
rect 8703 -10117 8763 -10057
rect 9023 -10117 9083 -10057
rect 9161 -10117 9221 -10057
rect 9481 -10117 9541 -10057
rect 9617 -10117 9677 -10057
rect 9937 -10117 9997 -10057
rect 10073 -10117 10133 -10057
rect 10393 -10117 10453 -10057
rect 10531 -10117 10591 -10057
rect 10851 -10117 10911 -10057
rect 10987 -10117 11047 -10057
rect 11307 -10117 11367 -10057
rect 11443 -10117 11503 -10057
rect 11763 -10117 11823 -10057
rect 11901 -10117 11961 -10057
rect 12221 -10117 12281 -10057
rect 12357 -10117 12417 -10057
rect 12677 -10117 12737 -10057
rect 12813 -10117 12873 -10057
rect 13133 -10117 13193 -10057
rect 13271 -10117 13331 -10057
rect 13591 -10117 13651 -10057
rect 13727 -10117 13787 -10057
rect 14047 -10117 14107 -10057
rect 14183 -10117 14243 -10057
rect 14503 -10117 14563 -10057
rect 14641 -10117 14701 -10057
rect 14961 -10117 15021 -10057
rect 15097 -10117 15157 -10057
rect 15417 -10117 15477 -10057
rect 7317 -10467 7377 -10407
rect 7637 -10467 7697 -10407
rect 7773 -10467 7833 -10407
rect 8093 -10467 8153 -10407
rect 8247 -10467 8307 -10407
rect 8567 -10467 8627 -10407
rect 8703 -10467 8763 -10407
rect 9023 -10467 9083 -10407
rect 9161 -10467 9221 -10407
rect 9481 -10467 9541 -10407
rect 9617 -10467 9677 -10407
rect 9937 -10467 9997 -10407
rect 10073 -10467 10133 -10407
rect 10393 -10467 10453 -10407
rect 10531 -10467 10591 -10407
rect 10851 -10467 10911 -10407
rect 10987 -10467 11047 -10407
rect 11307 -10467 11367 -10407
rect 11443 -10467 11503 -10407
rect 11763 -10467 11823 -10407
rect 11901 -10467 11961 -10407
rect 12221 -10467 12281 -10407
rect 12357 -10467 12417 -10407
rect 12677 -10467 12737 -10407
rect 12813 -10467 12873 -10407
rect 13133 -10467 13193 -10407
rect 13271 -10467 13331 -10407
rect 13591 -10467 13651 -10407
rect 13727 -10467 13787 -10407
rect 14047 -10467 14107 -10407
rect 14183 -10467 14243 -10407
rect 14503 -10467 14563 -10407
rect 14641 -10467 14701 -10407
rect 14961 -10467 15021 -10407
rect 15097 -10467 15157 -10407
rect 15417 -10467 15477 -10407
rect 11 -10619 14 -10559
rect 14 -10619 66 -10559
rect 66 -10619 71 -10559
rect 331 -10619 391 -10559
rect 11 -10969 14 -10909
rect 14 -10969 66 -10909
rect 66 -10969 71 -10909
rect 331 -10969 391 -10909
rect 467 -10619 527 -10559
rect 787 -10619 847 -10559
rect 923 -10619 983 -10559
rect 1243 -10619 1303 -10559
rect 1381 -10619 1441 -10559
rect 1701 -10619 1761 -10559
rect 1837 -10619 1897 -10559
rect 2157 -10619 2217 -10559
rect 2293 -10619 2353 -10559
rect 2613 -10619 2673 -10559
rect 2751 -10619 2811 -10559
rect 3071 -10619 3131 -10559
rect 3207 -10619 3267 -10559
rect 3527 -10619 3587 -10559
rect 3663 -10619 3723 -10559
rect 3983 -10619 4043 -10559
rect 467 -10969 527 -10909
rect 787 -10969 847 -10909
rect 923 -10969 983 -10909
rect 1243 -10969 1303 -10909
rect 1381 -10969 1441 -10909
rect 1701 -10969 1761 -10909
rect 1837 -10969 1897 -10909
rect 2157 -10969 2217 -10909
rect 2293 -10969 2353 -10909
rect 2613 -10969 2673 -10909
rect 2751 -10969 2811 -10909
rect 3071 -10969 3131 -10909
rect 3207 -10969 3267 -10909
rect 3527 -10969 3587 -10909
rect 3663 -10969 3723 -10909
rect 3983 -10969 4043 -10909
rect 4121 -10619 4181 -10559
rect 4441 -10619 4501 -10559
rect 4577 -10619 4637 -10559
rect 4897 -10619 4957 -10559
rect 5033 -10619 5093 -10559
rect 5353 -10619 5413 -10559
rect 5491 -10619 5551 -10559
rect 5811 -10619 5871 -10559
rect 5947 -10619 6007 -10559
rect 6267 -10619 6327 -10559
rect 6403 -10619 6463 -10559
rect 6723 -10619 6783 -10559
rect 6861 -10619 6921 -10559
rect 7181 -10619 7241 -10559
rect 4121 -10969 4181 -10909
rect 4441 -10969 4501 -10909
rect 4577 -10969 4637 -10909
rect 4897 -10969 4957 -10909
rect 5033 -10969 5093 -10909
rect 5353 -10969 5413 -10909
rect 5491 -10969 5551 -10909
rect 5811 -10969 5871 -10909
rect 5947 -10969 6007 -10909
rect 6267 -10969 6327 -10909
rect 6403 -10969 6463 -10909
rect 6723 -10969 6783 -10909
rect 6861 -10969 6921 -10909
rect 7181 -10969 7241 -10909
rect 7317 -10619 7377 -10559
rect 7637 -10619 7697 -10559
rect 7773 -10619 7833 -10559
rect 8093 -10619 8153 -10559
rect 8247 -10619 8307 -10559
rect 8567 -10619 8627 -10559
rect 8703 -10619 8763 -10559
rect 9023 -10619 9083 -10559
rect 9161 -10619 9221 -10559
rect 9481 -10619 9541 -10559
rect 9617 -10619 9677 -10559
rect 9937 -10619 9997 -10559
rect 10073 -10619 10133 -10559
rect 10393 -10619 10453 -10559
rect 10531 -10619 10591 -10559
rect 10851 -10619 10911 -10559
rect 10987 -10619 11047 -10559
rect 11307 -10619 11367 -10559
rect 11443 -10619 11503 -10559
rect 11763 -10619 11823 -10559
rect 11901 -10619 11961 -10559
rect 12221 -10619 12281 -10559
rect 12357 -10619 12417 -10559
rect 12677 -10619 12737 -10559
rect 12813 -10619 12873 -10559
rect 13133 -10619 13193 -10559
rect 13271 -10619 13331 -10559
rect 13591 -10619 13651 -10559
rect 13727 -10619 13787 -10559
rect 14047 -10619 14107 -10559
rect 14183 -10619 14243 -10559
rect 14503 -10619 14563 -10559
rect 14641 -10619 14701 -10559
rect 14961 -10619 15021 -10559
rect 15097 -10619 15157 -10559
rect 15417 -10619 15477 -10559
rect 7317 -10969 7377 -10909
rect 7637 -10969 7697 -10909
rect 7773 -10969 7833 -10909
rect 8093 -10969 8153 -10909
rect 8247 -10969 8307 -10909
rect 8567 -10969 8627 -10909
rect 8703 -10969 8763 -10909
rect 9023 -10969 9083 -10909
rect 9161 -10969 9221 -10909
rect 9481 -10969 9541 -10909
rect 9617 -10969 9677 -10909
rect 9937 -10969 9997 -10909
rect 10073 -10969 10133 -10909
rect 10393 -10969 10453 -10909
rect 10531 -10969 10591 -10909
rect 10851 -10969 10911 -10909
rect 10987 -10969 11047 -10909
rect 11307 -10969 11367 -10909
rect 11443 -10969 11503 -10909
rect 11763 -10969 11823 -10909
rect 11901 -10969 11961 -10909
rect 12221 -10969 12281 -10909
rect 12357 -10969 12417 -10909
rect 12677 -10969 12737 -10909
rect 12813 -10969 12873 -10909
rect 13133 -10969 13193 -10909
rect 13271 -10969 13331 -10909
rect 13591 -10969 13651 -10909
rect 13727 -10969 13787 -10909
rect 14047 -10969 14107 -10909
rect 14183 -10969 14243 -10909
rect 14503 -10969 14563 -10909
rect 14641 -10969 14701 -10909
rect 14961 -10969 15021 -10909
rect 15097 -10969 15157 -10909
rect 15417 -10969 15477 -10909
rect 11 -11111 14 -11051
rect 14 -11111 66 -11051
rect 66 -11111 71 -11051
rect 331 -11111 391 -11051
rect 11 -11461 14 -11401
rect 14 -11461 66 -11401
rect 66 -11461 71 -11401
rect 331 -11461 391 -11401
rect 467 -11111 527 -11051
rect 787 -11111 847 -11051
rect 923 -11111 983 -11051
rect 1243 -11111 1303 -11051
rect 1381 -11111 1441 -11051
rect 1701 -11111 1761 -11051
rect 1837 -11111 1897 -11051
rect 2157 -11111 2217 -11051
rect 2293 -11111 2353 -11051
rect 2613 -11111 2673 -11051
rect 2751 -11111 2811 -11051
rect 3071 -11111 3131 -11051
rect 3207 -11111 3267 -11051
rect 3527 -11111 3587 -11051
rect 3663 -11111 3723 -11051
rect 3983 -11111 4043 -11051
rect 467 -11461 527 -11401
rect 787 -11461 847 -11401
rect 923 -11461 983 -11401
rect 1243 -11461 1303 -11401
rect 1381 -11461 1441 -11401
rect 1701 -11461 1761 -11401
rect 1837 -11461 1897 -11401
rect 2157 -11461 2217 -11401
rect 2293 -11461 2353 -11401
rect 2613 -11461 2673 -11401
rect 2751 -11461 2811 -11401
rect 3071 -11461 3131 -11401
rect 3207 -11461 3267 -11401
rect 3527 -11461 3587 -11401
rect 3663 -11461 3723 -11401
rect 3983 -11461 4043 -11401
rect 4121 -11111 4181 -11051
rect 4441 -11111 4501 -11051
rect 4577 -11111 4637 -11051
rect 4897 -11111 4957 -11051
rect 5033 -11111 5093 -11051
rect 5353 -11111 5413 -11051
rect 5491 -11111 5551 -11051
rect 5811 -11111 5871 -11051
rect 5947 -11111 6007 -11051
rect 6267 -11111 6327 -11051
rect 6403 -11111 6463 -11051
rect 6723 -11111 6783 -11051
rect 6861 -11111 6921 -11051
rect 7181 -11111 7241 -11051
rect 4121 -11461 4181 -11401
rect 4441 -11461 4501 -11401
rect 4577 -11461 4637 -11401
rect 4897 -11461 4957 -11401
rect 5033 -11461 5093 -11401
rect 5353 -11461 5413 -11401
rect 5491 -11461 5551 -11401
rect 5811 -11461 5871 -11401
rect 5947 -11461 6007 -11401
rect 6267 -11461 6327 -11401
rect 6403 -11461 6463 -11401
rect 6723 -11461 6783 -11401
rect 6861 -11461 6921 -11401
rect 7181 -11461 7241 -11401
rect 7317 -11111 7377 -11051
rect 7637 -11111 7697 -11051
rect 7773 -11111 7833 -11051
rect 8093 -11111 8153 -11051
rect 8247 -11111 8307 -11051
rect 8567 -11111 8627 -11051
rect 8703 -11111 8763 -11051
rect 9023 -11111 9083 -11051
rect 9161 -11111 9221 -11051
rect 9481 -11111 9541 -11051
rect 9617 -11111 9677 -11051
rect 9937 -11111 9997 -11051
rect 7317 -11461 7377 -11401
rect 7637 -11461 7697 -11401
rect 7773 -11461 7833 -11401
rect 8093 -11461 8153 -11401
rect 8247 -11461 8307 -11401
rect 8567 -11461 8627 -11401
rect 8703 -11461 8763 -11401
rect 9023 -11461 9083 -11401
rect 9161 -11461 9221 -11401
rect 9481 -11461 9541 -11401
rect 10073 -11111 10133 -11051
rect 10393 -11111 10453 -11051
rect 10531 -11111 10591 -11051
rect 10851 -11111 10911 -11051
rect 10987 -11111 11047 -11051
rect 11307 -11111 11367 -11051
rect 11443 -11111 11503 -11051
rect 11763 -11111 11823 -11051
rect 11901 -11111 11961 -11051
rect 12221 -11111 12281 -11051
rect 12357 -11111 12417 -11051
rect 12677 -11111 12737 -11051
rect 12813 -11111 12873 -11051
rect 13133 -11111 13193 -11051
rect 13271 -11111 13331 -11051
rect 13591 -11111 13651 -11051
rect 13727 -11111 13787 -11051
rect 14047 -11111 14107 -11051
rect 14183 -11111 14243 -11051
rect 14503 -11111 14563 -11051
rect 14641 -11111 14701 -11051
rect 14961 -11111 15021 -11051
rect 15097 -11111 15157 -11051
rect 15417 -11111 15477 -11051
rect 9617 -11461 9677 -11401
rect 9937 -11461 9997 -11401
rect 10073 -11461 10133 -11401
rect 10393 -11461 10453 -11401
rect 10531 -11461 10591 -11401
rect 10851 -11461 10911 -11401
rect 10987 -11461 11047 -11401
rect 11307 -11461 11367 -11401
rect 11443 -11461 11503 -11401
rect 11763 -11461 11823 -11401
rect 11901 -11461 11961 -11401
rect 12221 -11461 12281 -11401
rect 12357 -11461 12417 -11401
rect 12677 -11461 12737 -11401
rect 12813 -11461 12873 -11401
rect 13133 -11461 13193 -11401
rect 13271 -11461 13331 -11401
rect 13591 -11461 13651 -11401
rect 13727 -11461 13787 -11401
rect 14047 -11461 14107 -11401
rect 14183 -11461 14243 -11401
rect 14503 -11461 14563 -11401
rect 14641 -11461 14701 -11401
rect 14961 -11461 15021 -11401
rect 15097 -11461 15157 -11401
rect 15417 -11461 15477 -11401
rect 10 -11604 14 -11544
rect 14 -11604 66 -11544
rect 66 -11604 70 -11544
rect 330 -11604 390 -11544
rect 10 -11954 14 -11894
rect 14 -11954 66 -11894
rect 66 -11954 70 -11894
rect 330 -11954 390 -11894
rect 466 -11604 526 -11544
rect 786 -11604 846 -11544
rect 922 -11604 982 -11544
rect 1242 -11604 1302 -11544
rect 1380 -11604 1440 -11544
rect 1700 -11604 1760 -11544
rect 1836 -11604 1896 -11544
rect 2156 -11604 2216 -11544
rect 2292 -11604 2352 -11544
rect 2612 -11604 2672 -11544
rect 2750 -11604 2810 -11544
rect 3070 -11604 3130 -11544
rect 3206 -11604 3266 -11544
rect 3526 -11604 3586 -11544
rect 3662 -11604 3722 -11544
rect 3982 -11604 4042 -11544
rect 466 -11954 526 -11894
rect 786 -11954 846 -11894
rect 922 -11954 982 -11894
rect 1242 -11954 1302 -11894
rect 1380 -11954 1440 -11894
rect 1700 -11954 1760 -11894
rect 1836 -11954 1896 -11894
rect 2156 -11954 2216 -11894
rect 2292 -11954 2352 -11894
rect 2612 -11954 2672 -11894
rect 2750 -11954 2810 -11894
rect 3070 -11954 3130 -11894
rect 3206 -11954 3266 -11894
rect 3526 -11954 3586 -11894
rect 3662 -11954 3722 -11894
rect 3982 -11954 4042 -11894
rect 4120 -11604 4180 -11544
rect 4440 -11604 4500 -11544
rect 4576 -11604 4636 -11544
rect 4896 -11604 4956 -11544
rect 5032 -11604 5092 -11544
rect 5352 -11604 5412 -11544
rect 5490 -11604 5550 -11544
rect 5810 -11604 5870 -11544
rect 5946 -11604 6006 -11544
rect 6266 -11604 6326 -11544
rect 6402 -11604 6462 -11544
rect 6722 -11604 6782 -11544
rect 6860 -11604 6920 -11544
rect 7180 -11604 7240 -11544
rect 4120 -11954 4180 -11894
rect 4440 -11954 4500 -11894
rect 4576 -11954 4636 -11894
rect 4896 -11954 4956 -11894
rect 5032 -11954 5092 -11894
rect 5352 -11954 5412 -11894
rect 5490 -11954 5550 -11894
rect 5810 -11954 5870 -11894
rect 5946 -11954 6006 -11894
rect 6266 -11954 6326 -11894
rect 6402 -11954 6462 -11894
rect 6722 -11954 6782 -11894
rect 6860 -11954 6920 -11894
rect 7180 -11954 7240 -11894
rect 7316 -11604 7376 -11544
rect 7636 -11604 7696 -11544
rect 7772 -11604 7832 -11544
rect 8092 -11604 8152 -11544
rect 8246 -11604 8306 -11544
rect 8566 -11604 8626 -11544
rect 8702 -11604 8762 -11544
rect 9022 -11604 9082 -11544
rect 9160 -11604 9220 -11544
rect 9480 -11604 9540 -11544
rect 7316 -11954 7376 -11894
rect 7636 -11954 7696 -11894
rect 7772 -11954 7832 -11894
rect 8092 -11954 8152 -11894
rect 8246 -11954 8306 -11894
rect 8566 -11954 8626 -11894
rect 8702 -11954 8762 -11894
rect 9022 -11954 9082 -11894
rect 9616 -11604 9676 -11544
rect 9936 -11604 9996 -11544
rect 10072 -11604 10132 -11544
rect 10392 -11604 10452 -11544
rect 10530 -11604 10590 -11544
rect 10850 -11604 10910 -11544
rect 10986 -11604 11046 -11544
rect 11306 -11604 11366 -11544
rect 11442 -11604 11502 -11544
rect 11762 -11604 11822 -11544
rect 11900 -11604 11960 -11544
rect 12220 -11604 12280 -11544
rect 12356 -11604 12416 -11544
rect 12676 -11604 12736 -11544
rect 12812 -11604 12872 -11544
rect 13132 -11604 13192 -11544
rect 13270 -11604 13330 -11544
rect 13590 -11604 13650 -11544
rect 13726 -11604 13786 -11544
rect 14046 -11604 14106 -11544
rect 14182 -11604 14242 -11544
rect 14502 -11604 14562 -11544
rect 14640 -11604 14700 -11544
rect 14960 -11604 15020 -11544
rect 15096 -11604 15156 -11544
rect 15416 -11604 15476 -11544
rect 9160 -11954 9220 -11894
rect 9480 -11954 9540 -11894
rect 9616 -11954 9676 -11894
rect 9936 -11954 9996 -11894
rect 10072 -11954 10132 -11894
rect 10392 -11954 10452 -11894
rect 10530 -11954 10590 -11894
rect 10850 -11954 10910 -11894
rect 10986 -11954 11046 -11894
rect 11306 -11954 11366 -11894
rect 11442 -11954 11502 -11894
rect 11762 -11954 11822 -11894
rect 11900 -11954 11960 -11894
rect 12220 -11954 12280 -11894
rect 12356 -11954 12416 -11894
rect 12676 -11954 12736 -11894
rect 12812 -11954 12872 -11894
rect 13132 -11954 13192 -11894
rect 13270 -11954 13330 -11894
rect 13590 -11954 13650 -11894
rect 13726 -11954 13786 -11894
rect 14046 -11954 14106 -11894
rect 14182 -11954 14242 -11894
rect 14502 -11954 14562 -11894
rect 14640 -11954 14700 -11894
rect 14960 -11954 15020 -11894
rect 15096 -11954 15156 -11894
rect 15416 -11954 15476 -11894
rect 10 -12096 14 -12036
rect 14 -12096 66 -12036
rect 66 -12096 70 -12036
rect 330 -12096 390 -12036
rect 10 -12446 14 -12386
rect 14 -12446 66 -12386
rect 66 -12446 70 -12386
rect 330 -12446 390 -12386
rect 466 -12096 526 -12036
rect 786 -12096 846 -12036
rect 922 -12096 982 -12036
rect 1242 -12096 1302 -12036
rect 1380 -12096 1440 -12036
rect 1700 -12096 1760 -12036
rect 1836 -12096 1896 -12036
rect 2156 -12096 2216 -12036
rect 2292 -12096 2352 -12036
rect 2612 -12096 2672 -12036
rect 2750 -12096 2810 -12036
rect 3070 -12096 3130 -12036
rect 3206 -12096 3266 -12036
rect 3526 -12096 3586 -12036
rect 466 -12446 526 -12386
rect 786 -12446 846 -12386
rect 922 -12446 982 -12386
rect 1242 -12446 1302 -12386
rect 1380 -12446 1440 -12386
rect 1700 -12446 1760 -12386
rect 1836 -12446 1896 -12386
rect 2156 -12446 2216 -12386
rect 2292 -12446 2352 -12386
rect 2612 -12446 2672 -12386
rect 2750 -12446 2810 -12386
rect 3070 -12446 3130 -12386
rect 3206 -12446 3266 -12386
rect 3526 -12446 3586 -12386
rect 3662 -12096 3722 -12036
rect 3982 -12096 4042 -12036
rect 4120 -12096 4180 -12036
rect 4440 -12096 4500 -12036
rect 4576 -12096 4636 -12036
rect 4896 -12096 4956 -12036
rect 5032 -12096 5092 -12036
rect 5352 -12096 5412 -12036
rect 5490 -12096 5550 -12036
rect 5810 -12096 5870 -12036
rect 5946 -12096 6006 -12036
rect 6266 -12096 6326 -12036
rect 6402 -12096 6462 -12036
rect 6722 -12096 6782 -12036
rect 6860 -12096 6920 -12036
rect 7180 -12096 7240 -12036
rect 3662 -12446 3722 -12386
rect 3982 -12446 4042 -12386
rect 4120 -12446 4180 -12386
rect 4440 -12446 4500 -12386
rect 4576 -12446 4636 -12386
rect 4896 -12446 4956 -12386
rect 5032 -12446 5092 -12386
rect 5352 -12446 5412 -12386
rect 5490 -12446 5550 -12386
rect 5810 -12446 5870 -12386
rect 5946 -12446 6006 -12386
rect 6266 -12446 6326 -12386
rect 6402 -12446 6462 -12386
rect 6722 -12446 6782 -12386
rect 6860 -12446 6920 -12386
rect 7180 -12446 7240 -12386
rect 7316 -12096 7376 -12036
rect 7636 -12096 7696 -12036
rect 7772 -12096 7832 -12036
rect 8092 -12096 8152 -12036
rect 8246 -12096 8306 -12036
rect 8566 -12096 8626 -12036
rect 8702 -12096 8762 -12036
rect 9022 -12096 9082 -12036
rect 9160 -12096 9220 -12036
rect 9480 -12096 9540 -12036
rect 9616 -12096 9676 -12036
rect 9936 -12096 9996 -12036
rect 10072 -12096 10132 -12036
rect 10392 -12096 10452 -12036
rect 10530 -12096 10590 -12036
rect 10850 -12096 10910 -12036
rect 10986 -12096 11046 -12036
rect 11306 -12096 11366 -12036
rect 11442 -12096 11502 -12036
rect 11762 -12096 11822 -12036
rect 11900 -12096 11960 -12036
rect 12220 -12096 12280 -12036
rect 12356 -12096 12416 -12036
rect 12676 -12096 12736 -12036
rect 12812 -12096 12872 -12036
rect 13132 -12096 13192 -12036
rect 13270 -12096 13330 -12036
rect 13590 -12096 13650 -12036
rect 13726 -12096 13786 -12036
rect 14046 -12096 14106 -12036
rect 14182 -12096 14242 -12036
rect 14502 -12096 14562 -12036
rect 14640 -12096 14700 -12036
rect 14960 -12096 15020 -12036
rect 15096 -12096 15156 -12036
rect 15416 -12096 15476 -12036
rect 7316 -12446 7376 -12386
rect 7636 -12446 7696 -12386
rect 7772 -12446 7832 -12386
rect 8092 -12446 8152 -12386
rect 8246 -12446 8306 -12386
rect 8566 -12446 8626 -12386
rect 8702 -12446 8762 -12386
rect 9022 -12446 9082 -12386
rect 9160 -12446 9220 -12386
rect 9480 -12446 9540 -12386
rect 9616 -12446 9676 -12386
rect 9936 -12446 9996 -12386
rect 10072 -12446 10132 -12386
rect 10392 -12446 10452 -12386
rect 10530 -12446 10590 -12386
rect 10850 -12446 10910 -12386
rect 10986 -12446 11046 -12386
rect 11306 -12446 11366 -12386
rect 11442 -12446 11502 -12386
rect 11762 -12446 11822 -12386
rect 11900 -12446 11960 -12386
rect 12220 -12446 12280 -12386
rect 12356 -12446 12416 -12386
rect 12676 -12446 12736 -12386
rect 12812 -12446 12872 -12386
rect 13132 -12446 13192 -12386
rect 13270 -12446 13330 -12386
rect 13590 -12446 13650 -12386
rect 13726 -12446 13786 -12386
rect 14046 -12446 14106 -12386
rect 14182 -12446 14242 -12386
rect 14502 -12446 14562 -12386
rect 14640 -12446 14700 -12386
rect 14960 -12446 15020 -12386
rect 15096 -12446 15156 -12386
rect 15416 -12446 15476 -12386
rect 10 -12612 14 -12552
rect 14 -12612 66 -12552
rect 66 -12612 70 -12552
rect 330 -12612 390 -12552
rect 10 -12962 14 -12902
rect 14 -12962 66 -12902
rect 66 -12962 70 -12902
rect 330 -12962 390 -12902
rect 466 -12612 526 -12552
rect 786 -12612 846 -12552
rect 922 -12612 982 -12552
rect 1242 -12612 1302 -12552
rect 1380 -12612 1440 -12552
rect 1700 -12612 1760 -12552
rect 1836 -12612 1896 -12552
rect 2156 -12612 2216 -12552
rect 2292 -12612 2352 -12552
rect 2612 -12612 2672 -12552
rect 2750 -12612 2810 -12552
rect 3070 -12612 3130 -12552
rect 3206 -12612 3266 -12552
rect 3526 -12612 3586 -12552
rect 466 -12962 526 -12902
rect 786 -12962 846 -12902
rect 922 -12962 982 -12902
rect 1242 -12962 1302 -12902
rect 1380 -12962 1440 -12902
rect 1700 -12962 1760 -12902
rect 1836 -12962 1896 -12902
rect 2156 -12962 2216 -12902
rect 2292 -12962 2352 -12902
rect 2612 -12962 2672 -12902
rect 2750 -12962 2810 -12902
rect 3070 -12962 3130 -12902
rect 3206 -12962 3266 -12902
rect 3526 -12962 3586 -12902
rect 3662 -12612 3722 -12552
rect 3982 -12612 4042 -12552
rect 4120 -12612 4180 -12552
rect 4440 -12612 4500 -12552
rect 4576 -12612 4636 -12552
rect 4896 -12612 4956 -12552
rect 5032 -12612 5092 -12552
rect 5352 -12612 5412 -12552
rect 5490 -12612 5550 -12552
rect 5810 -12612 5870 -12552
rect 5946 -12612 6006 -12552
rect 6266 -12612 6326 -12552
rect 6402 -12612 6462 -12552
rect 6722 -12612 6782 -12552
rect 6860 -12612 6920 -12552
rect 7180 -12612 7240 -12552
rect 3662 -12962 3722 -12902
rect 3982 -12962 4042 -12902
rect 4120 -12962 4180 -12902
rect 4440 -12962 4500 -12902
rect 4576 -12962 4636 -12902
rect 4896 -12962 4956 -12902
rect 5032 -12962 5092 -12902
rect 5352 -12962 5412 -12902
rect 5490 -12962 5550 -12902
rect 5810 -12962 5870 -12902
rect 5946 -12962 6006 -12902
rect 6266 -12962 6326 -12902
rect 6402 -12962 6462 -12902
rect 6722 -12962 6782 -12902
rect 6860 -12962 6920 -12902
rect 7180 -12962 7240 -12902
rect 7316 -12612 7376 -12552
rect 7636 -12612 7696 -12552
rect 7772 -12612 7832 -12552
rect 8092 -12612 8152 -12552
rect 8246 -12612 8306 -12552
rect 8566 -12612 8626 -12552
rect 8702 -12612 8762 -12552
rect 9022 -12612 9082 -12552
rect 9160 -12612 9220 -12552
rect 9480 -12612 9540 -12552
rect 9616 -12612 9676 -12552
rect 9936 -12612 9996 -12552
rect 10072 -12612 10132 -12552
rect 10392 -12612 10452 -12552
rect 10530 -12612 10590 -12552
rect 10850 -12612 10910 -12552
rect 7316 -12962 7376 -12902
rect 7636 -12962 7696 -12902
rect 7772 -12962 7832 -12902
rect 8092 -12962 8152 -12902
rect 8246 -12962 8306 -12902
rect 8566 -12962 8626 -12902
rect 8702 -12962 8762 -12902
rect 9022 -12962 9082 -12902
rect 9160 -12962 9220 -12902
rect 9480 -12962 9540 -12902
rect 9616 -12962 9676 -12902
rect 9936 -12962 9996 -12902
rect 10072 -12962 10132 -12902
rect 10392 -12962 10452 -12902
rect 10530 -12962 10590 -12902
rect 10850 -12962 10910 -12902
rect 10986 -12612 11046 -12552
rect 11306 -12612 11366 -12552
rect 11442 -12612 11502 -12552
rect 11762 -12612 11822 -12552
rect 11900 -12612 11960 -12552
rect 12220 -12612 12280 -12552
rect 12356 -12612 12416 -12552
rect 12676 -12612 12736 -12552
rect 12812 -12612 12872 -12552
rect 13132 -12612 13192 -12552
rect 13270 -12612 13330 -12552
rect 13590 -12612 13650 -12552
rect 13726 -12612 13786 -12552
rect 14046 -12612 14106 -12552
rect 14182 -12612 14242 -12552
rect 14502 -12612 14562 -12552
rect 14640 -12612 14700 -12552
rect 14960 -12612 15020 -12552
rect 15096 -12612 15156 -12552
rect 15416 -12612 15476 -12552
rect 10986 -12962 11046 -12902
rect 11306 -12962 11366 -12902
rect 11442 -12962 11502 -12902
rect 11762 -12962 11822 -12902
rect 11900 -12962 11960 -12902
rect 12220 -12962 12280 -12902
rect 12356 -12962 12416 -12902
rect 12676 -12962 12736 -12902
rect 12812 -12962 12872 -12902
rect 13132 -12962 13192 -12902
rect 13270 -12962 13330 -12902
rect 13590 -12962 13650 -12902
rect 13726 -12962 13786 -12902
rect 14046 -12962 14106 -12902
rect 14182 -12962 14242 -12902
rect 14502 -12962 14562 -12902
rect 14640 -12962 14700 -12902
rect 14960 -12962 15020 -12902
rect 15096 -12962 15156 -12902
rect 15416 -12962 15476 -12902
rect 10 -13114 14 -13054
rect 14 -13114 66 -13054
rect 66 -13114 70 -13054
rect 330 -13114 390 -13054
rect 10 -13464 14 -13404
rect 14 -13464 66 -13404
rect 66 -13464 70 -13404
rect 330 -13464 390 -13404
rect 466 -13114 526 -13054
rect 786 -13114 846 -13054
rect 922 -13114 982 -13054
rect 1242 -13114 1302 -13054
rect 1380 -13114 1440 -13054
rect 1700 -13114 1760 -13054
rect 1836 -13114 1896 -13054
rect 2156 -13114 2216 -13054
rect 2292 -13114 2352 -13054
rect 2612 -13114 2672 -13054
rect 2750 -13114 2810 -13054
rect 3070 -13114 3130 -13054
rect 3206 -13114 3266 -13054
rect 3526 -13114 3586 -13054
rect 466 -13464 526 -13404
rect 786 -13464 846 -13404
rect 922 -13464 982 -13404
rect 1242 -13464 1302 -13404
rect 1380 -13464 1440 -13404
rect 1700 -13464 1760 -13404
rect 1836 -13464 1896 -13404
rect 2156 -13464 2216 -13404
rect 2292 -13464 2352 -13404
rect 2612 -13464 2672 -13404
rect 2750 -13464 2810 -13404
rect 3070 -13464 3130 -13404
rect 3206 -13464 3266 -13404
rect 3526 -13464 3586 -13404
rect 3662 -13114 3722 -13054
rect 3982 -13114 4042 -13054
rect 4120 -13114 4180 -13054
rect 4440 -13114 4500 -13054
rect 4576 -13114 4636 -13054
rect 4896 -13114 4956 -13054
rect 5032 -13114 5092 -13054
rect 5352 -13114 5412 -13054
rect 5490 -13114 5550 -13054
rect 5810 -13114 5870 -13054
rect 5946 -13114 6006 -13054
rect 6266 -13114 6326 -13054
rect 6402 -13114 6462 -13054
rect 6722 -13114 6782 -13054
rect 6860 -13114 6920 -13054
rect 7180 -13114 7240 -13054
rect 3662 -13464 3722 -13404
rect 3982 -13464 4042 -13404
rect 4120 -13464 4180 -13404
rect 4440 -13464 4500 -13404
rect 4576 -13464 4636 -13404
rect 4896 -13464 4956 -13404
rect 5032 -13464 5092 -13404
rect 5352 -13464 5412 -13404
rect 5490 -13464 5550 -13404
rect 5810 -13464 5870 -13404
rect 5946 -13464 6006 -13404
rect 6266 -13464 6326 -13404
rect 6402 -13464 6462 -13404
rect 6722 -13464 6782 -13404
rect 6860 -13464 6920 -13404
rect 7180 -13464 7240 -13404
rect 7316 -13114 7376 -13054
rect 7636 -13114 7696 -13054
rect 7772 -13114 7832 -13054
rect 8092 -13114 8152 -13054
rect 8246 -13114 8306 -13054
rect 8566 -13114 8626 -13054
rect 8702 -13114 8762 -13054
rect 9022 -13114 9082 -13054
rect 9160 -13114 9220 -13054
rect 9480 -13114 9540 -13054
rect 9616 -13114 9676 -13054
rect 9936 -13114 9996 -13054
rect 10072 -13114 10132 -13054
rect 10392 -13114 10452 -13054
rect 10530 -13114 10590 -13054
rect 10850 -13114 10910 -13054
rect 7316 -13464 7376 -13404
rect 7636 -13464 7696 -13404
rect 7772 -13464 7832 -13404
rect 8092 -13464 8152 -13404
rect 8246 -13464 8306 -13404
rect 8566 -13464 8626 -13404
rect 8702 -13464 8762 -13404
rect 9022 -13464 9082 -13404
rect 9160 -13464 9220 -13404
rect 9480 -13464 9540 -13404
rect 9616 -13464 9676 -13404
rect 9936 -13464 9996 -13404
rect 10072 -13464 10132 -13404
rect 10392 -13464 10452 -13404
rect 10530 -13464 10590 -13404
rect 10850 -13464 10910 -13404
rect 10986 -13114 11046 -13054
rect 11306 -13114 11366 -13054
rect 11442 -13114 11502 -13054
rect 11762 -13114 11822 -13054
rect 11900 -13114 11960 -13054
rect 12220 -13114 12280 -13054
rect 12356 -13114 12416 -13054
rect 12676 -13114 12736 -13054
rect 12812 -13114 12872 -13054
rect 13132 -13114 13192 -13054
rect 13270 -13114 13330 -13054
rect 13590 -13114 13650 -13054
rect 13726 -13114 13786 -13054
rect 14046 -13114 14106 -13054
rect 14182 -13114 14242 -13054
rect 14502 -13114 14562 -13054
rect 14640 -13114 14700 -13054
rect 14960 -13114 15020 -13054
rect 15096 -13114 15156 -13054
rect 15416 -13114 15476 -13054
rect 10986 -13464 11046 -13404
rect 11306 -13464 11366 -13404
rect 11442 -13464 11502 -13404
rect 11762 -13464 11822 -13404
rect 11900 -13464 11960 -13404
rect 12220 -13464 12280 -13404
rect 12356 -13464 12416 -13404
rect 12676 -13464 12736 -13404
rect 12812 -13464 12872 -13404
rect 13132 -13464 13192 -13404
rect 13270 -13464 13330 -13404
rect 13590 -13464 13650 -13404
rect 13726 -13464 13786 -13404
rect 14046 -13464 14106 -13404
rect 14182 -13464 14242 -13404
rect 14502 -13464 14562 -13404
rect 14640 -13464 14700 -13404
rect 14960 -13464 15020 -13404
rect 15096 -13464 15156 -13404
rect 15416 -13464 15476 -13404
rect 10 -13606 14 -13546
rect 14 -13606 66 -13546
rect 66 -13606 70 -13546
rect 330 -13606 390 -13546
rect 10 -13956 14 -13896
rect 14 -13956 66 -13896
rect 66 -13956 70 -13896
rect 330 -13956 390 -13896
rect 466 -13606 526 -13546
rect 786 -13606 846 -13546
rect 922 -13606 982 -13546
rect 1242 -13606 1302 -13546
rect 1380 -13606 1440 -13546
rect 1700 -13606 1760 -13546
rect 1836 -13606 1896 -13546
rect 2156 -13606 2216 -13546
rect 2292 -13606 2352 -13546
rect 2612 -13606 2672 -13546
rect 2750 -13606 2810 -13546
rect 3070 -13606 3130 -13546
rect 3206 -13606 3266 -13546
rect 3526 -13606 3586 -13546
rect 466 -13956 526 -13896
rect 786 -13956 846 -13896
rect 922 -13956 982 -13896
rect 1242 -13956 1302 -13896
rect 1380 -13956 1440 -13896
rect 1700 -13956 1760 -13896
rect 1836 -13956 1896 -13896
rect 2156 -13956 2216 -13896
rect 2292 -13956 2352 -13896
rect 2612 -13956 2672 -13896
rect 2750 -13956 2810 -13896
rect 3070 -13956 3130 -13896
rect 3206 -13956 3266 -13896
rect 3526 -13956 3586 -13896
rect 3662 -13606 3722 -13546
rect 3982 -13606 4042 -13546
rect 4120 -13606 4180 -13546
rect 4440 -13606 4500 -13546
rect 4576 -13606 4636 -13546
rect 4896 -13606 4956 -13546
rect 5032 -13606 5092 -13546
rect 5352 -13606 5412 -13546
rect 5490 -13606 5550 -13546
rect 5810 -13606 5870 -13546
rect 5946 -13606 6006 -13546
rect 6266 -13606 6326 -13546
rect 6402 -13606 6462 -13546
rect 6722 -13606 6782 -13546
rect 6860 -13606 6920 -13546
rect 7180 -13606 7240 -13546
rect 3662 -13956 3722 -13896
rect 3982 -13956 4042 -13896
rect 4120 -13956 4180 -13896
rect 4440 -13956 4500 -13896
rect 4576 -13956 4636 -13896
rect 4896 -13956 4956 -13896
rect 5032 -13956 5092 -13896
rect 5352 -13956 5412 -13896
rect 5490 -13956 5550 -13896
rect 5810 -13956 5870 -13896
rect 5946 -13956 6006 -13896
rect 6266 -13956 6326 -13896
rect 6402 -13956 6462 -13896
rect 6722 -13956 6782 -13896
rect 6860 -13956 6920 -13896
rect 7180 -13956 7240 -13896
rect 7316 -13606 7376 -13546
rect 7636 -13606 7696 -13546
rect 7772 -13606 7832 -13546
rect 8092 -13606 8152 -13546
rect 8246 -13606 8306 -13546
rect 8566 -13606 8626 -13546
rect 8702 -13606 8762 -13546
rect 9022 -13606 9082 -13546
rect 9160 -13606 9220 -13546
rect 9480 -13606 9540 -13546
rect 9616 -13606 9676 -13546
rect 9936 -13606 9996 -13546
rect 10072 -13606 10132 -13546
rect 10392 -13606 10452 -13546
rect 10530 -13606 10590 -13546
rect 10850 -13606 10910 -13546
rect 7316 -13956 7376 -13896
rect 7636 -13956 7696 -13896
rect 7772 -13956 7832 -13896
rect 8092 -13956 8152 -13896
rect 8246 -13956 8306 -13896
rect 8566 -13956 8626 -13896
rect 8702 -13956 8762 -13896
rect 9022 -13956 9082 -13896
rect 9160 -13956 9220 -13896
rect 9480 -13956 9540 -13896
rect 9616 -13956 9676 -13896
rect 9936 -13956 9996 -13896
rect 10072 -13956 10132 -13896
rect 10392 -13956 10452 -13896
rect 10530 -13956 10590 -13896
rect 10850 -13956 10910 -13896
rect 10986 -13606 11046 -13546
rect 11306 -13606 11366 -13546
rect 11442 -13606 11502 -13546
rect 11762 -13606 11822 -13546
rect 11900 -13606 11960 -13546
rect 12220 -13606 12280 -13546
rect 10986 -13956 11046 -13896
rect 11306 -13956 11366 -13896
rect 11442 -13956 11502 -13896
rect 11762 -13956 11822 -13896
rect 11900 -13956 11960 -13896
rect 12220 -13956 12280 -13896
rect 12356 -13606 12416 -13546
rect 12676 -13606 12736 -13546
rect 12812 -13606 12872 -13546
rect 13132 -13606 13192 -13546
rect 13270 -13606 13330 -13546
rect 13590 -13606 13650 -13546
rect 13726 -13606 13786 -13546
rect 14046 -13606 14106 -13546
rect 14182 -13606 14242 -13546
rect 14502 -13606 14562 -13546
rect 14640 -13606 14700 -13546
rect 14960 -13606 15020 -13546
rect 15096 -13606 15156 -13546
rect 15416 -13606 15476 -13546
rect 12356 -13956 12416 -13896
rect 12676 -13956 12736 -13896
rect 12812 -13956 12872 -13896
rect 13132 -13956 13192 -13896
rect 13270 -13956 13330 -13896
rect 13590 -13956 13650 -13896
rect 13726 -13956 13786 -13896
rect 14046 -13956 14106 -13896
rect 14182 -13956 14242 -13896
rect 14502 -13956 14562 -13896
rect 14640 -13956 14700 -13896
rect 14960 -13956 15020 -13896
rect 15096 -13956 15156 -13896
rect 15416 -13956 15476 -13896
rect 10 -14100 14 -14040
rect 14 -14100 66 -14040
rect 66 -14100 70 -14040
rect 330 -14100 390 -14040
rect 10 -14450 14 -14390
rect 14 -14450 66 -14390
rect 66 -14450 70 -14390
rect 330 -14450 390 -14390
rect 466 -14100 526 -14040
rect 786 -14100 846 -14040
rect 922 -14100 982 -14040
rect 1242 -14100 1302 -14040
rect 1380 -14100 1440 -14040
rect 1700 -14100 1760 -14040
rect 1836 -14100 1896 -14040
rect 2156 -14100 2216 -14040
rect 2292 -14100 2352 -14040
rect 2612 -14100 2672 -14040
rect 2750 -14100 2810 -14040
rect 3070 -14100 3130 -14040
rect 3206 -14100 3266 -14040
rect 3526 -14100 3586 -14040
rect 466 -14450 526 -14390
rect 786 -14450 846 -14390
rect 922 -14450 982 -14390
rect 1242 -14450 1302 -14390
rect 1380 -14450 1440 -14390
rect 1700 -14450 1760 -14390
rect 1836 -14450 1896 -14390
rect 2156 -14450 2216 -14390
rect 2292 -14450 2352 -14390
rect 2612 -14450 2672 -14390
rect 2750 -14450 2810 -14390
rect 3070 -14450 3130 -14390
rect 3206 -14450 3266 -14390
rect 3526 -14450 3586 -14390
rect 3662 -14100 3722 -14040
rect 3982 -14100 4042 -14040
rect 4120 -14100 4180 -14040
rect 4440 -14100 4500 -14040
rect 4576 -14100 4636 -14040
rect 4896 -14100 4956 -14040
rect 5032 -14100 5092 -14040
rect 5352 -14100 5412 -14040
rect 5490 -14100 5550 -14040
rect 5810 -14100 5870 -14040
rect 5946 -14100 6006 -14040
rect 6266 -14100 6326 -14040
rect 6402 -14100 6462 -14040
rect 6722 -14100 6782 -14040
rect 6860 -14100 6920 -14040
rect 7180 -14100 7240 -14040
rect 3662 -14450 3722 -14390
rect 3982 -14450 4042 -14390
rect 4120 -14450 4180 -14390
rect 4440 -14450 4500 -14390
rect 4576 -14450 4636 -14390
rect 4896 -14450 4956 -14390
rect 5032 -14450 5092 -14390
rect 5352 -14450 5412 -14390
rect 5490 -14450 5550 -14390
rect 5810 -14450 5870 -14390
rect 5946 -14450 6006 -14390
rect 6266 -14450 6326 -14390
rect 6402 -14450 6462 -14390
rect 6722 -14450 6782 -14390
rect 6860 -14450 6920 -14390
rect 7180 -14450 7240 -14390
rect 7316 -14100 7376 -14040
rect 7636 -14100 7696 -14040
rect 7772 -14100 7832 -14040
rect 8092 -14100 8152 -14040
rect 8246 -14100 8306 -14040
rect 8566 -14100 8626 -14040
rect 8702 -14100 8762 -14040
rect 9022 -14100 9082 -14040
rect 9160 -14100 9220 -14040
rect 9480 -14100 9540 -14040
rect 9616 -14100 9676 -14040
rect 9936 -14100 9996 -14040
rect 10072 -14100 10132 -14040
rect 10392 -14100 10452 -14040
rect 10530 -14100 10590 -14040
rect 10850 -14100 10910 -14040
rect 7316 -14450 7376 -14390
rect 7636 -14450 7696 -14390
rect 7772 -14450 7832 -14390
rect 8092 -14450 8152 -14390
rect 8246 -14450 8306 -14390
rect 8566 -14450 8626 -14390
rect 8702 -14450 8762 -14390
rect 9022 -14450 9082 -14390
rect 9160 -14450 9220 -14390
rect 9480 -14450 9540 -14390
rect 9616 -14450 9676 -14390
rect 9936 -14450 9996 -14390
rect 10072 -14450 10132 -14390
rect 10392 -14450 10452 -14390
rect 10530 -14450 10590 -14390
rect 10850 -14450 10910 -14390
rect 10986 -14100 11046 -14040
rect 11306 -14100 11366 -14040
rect 11442 -14100 11502 -14040
rect 11762 -14100 11822 -14040
rect 11900 -14100 11960 -14040
rect 12220 -14100 12280 -14040
rect 10986 -14450 11046 -14390
rect 11306 -14450 11366 -14390
rect 11442 -14450 11502 -14390
rect 11762 -14450 11822 -14390
rect 11900 -14450 11960 -14390
rect 12220 -14450 12280 -14390
rect 12356 -14100 12416 -14040
rect 12676 -14100 12736 -14040
rect 12812 -14100 12872 -14040
rect 13132 -14100 13192 -14040
rect 12356 -14450 12416 -14390
rect 12676 -14450 12736 -14390
rect 12812 -14450 12872 -14390
rect 13132 -14450 13192 -14390
rect 13270 -14100 13330 -14040
rect 13590 -14100 13650 -14040
rect 13726 -14100 13786 -14040
rect 14046 -14100 14106 -14040
rect 14182 -14100 14242 -14040
rect 14502 -14100 14562 -14040
rect 14640 -14100 14700 -14040
rect 14960 -14100 15020 -14040
rect 15096 -14100 15156 -14040
rect 15416 -14100 15476 -14040
rect 13270 -14450 13330 -14390
rect 13590 -14450 13650 -14390
rect 13726 -14450 13786 -14390
rect 14046 -14450 14106 -14390
rect 14182 -14450 14242 -14390
rect 14502 -14450 14562 -14390
rect 14640 -14450 14700 -14390
rect 14960 -14450 15020 -14390
rect 15096 -14450 15156 -14390
rect 15416 -14450 15476 -14390
rect 10 -14602 14 -14542
rect 14 -14602 66 -14542
rect 66 -14602 70 -14542
rect 330 -14602 390 -14542
rect 10 -14952 14 -14892
rect 14 -14952 66 -14892
rect 66 -14952 70 -14892
rect 330 -14952 390 -14892
rect 466 -14602 526 -14542
rect 786 -14602 846 -14542
rect 922 -14602 982 -14542
rect 1242 -14602 1302 -14542
rect 1380 -14602 1440 -14542
rect 1700 -14602 1760 -14542
rect 1836 -14602 1896 -14542
rect 2156 -14602 2216 -14542
rect 2292 -14602 2352 -14542
rect 2612 -14602 2672 -14542
rect 2750 -14602 2810 -14542
rect 3070 -14602 3130 -14542
rect 3206 -14602 3266 -14542
rect 3526 -14602 3586 -14542
rect 466 -14952 526 -14892
rect 786 -14952 846 -14892
rect 922 -14952 982 -14892
rect 1242 -14952 1302 -14892
rect 1380 -14952 1440 -14892
rect 1700 -14952 1760 -14892
rect 1836 -14952 1896 -14892
rect 2156 -14952 2216 -14892
rect 2292 -14952 2352 -14892
rect 2612 -14952 2672 -14892
rect 2750 -14952 2810 -14892
rect 3070 -14952 3130 -14892
rect 3206 -14952 3266 -14892
rect 3526 -14952 3586 -14892
rect 3662 -14602 3722 -14542
rect 3982 -14602 4042 -14542
rect 4120 -14602 4180 -14542
rect 4440 -14602 4500 -14542
rect 4576 -14602 4636 -14542
rect 4896 -14602 4956 -14542
rect 5032 -14602 5092 -14542
rect 5352 -14602 5412 -14542
rect 5490 -14602 5550 -14542
rect 5810 -14602 5870 -14542
rect 5946 -14602 6006 -14542
rect 6266 -14602 6326 -14542
rect 6402 -14602 6462 -14542
rect 6722 -14602 6782 -14542
rect 6860 -14602 6920 -14542
rect 7180 -14602 7240 -14542
rect 3662 -14952 3722 -14892
rect 3982 -14952 4042 -14892
rect 4120 -14952 4180 -14892
rect 4440 -14952 4500 -14892
rect 4576 -14952 4636 -14892
rect 4896 -14952 4956 -14892
rect 5032 -14952 5092 -14892
rect 5352 -14952 5412 -14892
rect 5490 -14952 5550 -14892
rect 5810 -14952 5870 -14892
rect 5946 -14952 6006 -14892
rect 6266 -14952 6326 -14892
rect 6402 -14952 6462 -14892
rect 6722 -14952 6782 -14892
rect 6860 -14952 6920 -14892
rect 7180 -14952 7240 -14892
rect 7316 -14602 7376 -14542
rect 7636 -14602 7696 -14542
rect 7772 -14602 7832 -14542
rect 8092 -14602 8152 -14542
rect 8246 -14602 8306 -14542
rect 8566 -14602 8626 -14542
rect 8702 -14602 8762 -14542
rect 9022 -14602 9082 -14542
rect 9160 -14602 9220 -14542
rect 9480 -14602 9540 -14542
rect 9616 -14602 9676 -14542
rect 9936 -14602 9996 -14542
rect 10072 -14602 10132 -14542
rect 10392 -14602 10452 -14542
rect 10530 -14602 10590 -14542
rect 10850 -14602 10910 -14542
rect 7316 -14952 7376 -14892
rect 7636 -14952 7696 -14892
rect 7772 -14952 7832 -14892
rect 8092 -14952 8152 -14892
rect 8246 -14952 8306 -14892
rect 8566 -14952 8626 -14892
rect 8702 -14952 8762 -14892
rect 9022 -14952 9082 -14892
rect 9160 -14952 9220 -14892
rect 9480 -14952 9540 -14892
rect 9616 -14952 9676 -14892
rect 9936 -14952 9996 -14892
rect 10072 -14952 10132 -14892
rect 10392 -14952 10452 -14892
rect 10530 -14952 10590 -14892
rect 10850 -14952 10910 -14892
rect 10986 -14602 11046 -14542
rect 11306 -14602 11366 -14542
rect 11442 -14602 11502 -14542
rect 11762 -14602 11822 -14542
rect 11900 -14602 11960 -14542
rect 12220 -14602 12280 -14542
rect 10986 -14952 11046 -14892
rect 11306 -14952 11366 -14892
rect 11442 -14952 11502 -14892
rect 11762 -14952 11822 -14892
rect 11900 -14952 11960 -14892
rect 12220 -14952 12280 -14892
rect 12356 -14602 12416 -14542
rect 12676 -14602 12736 -14542
rect 12812 -14602 12872 -14542
rect 13132 -14602 13192 -14542
rect 12356 -14952 12416 -14892
rect 12676 -14952 12736 -14892
rect 12812 -14952 12872 -14892
rect 13132 -14952 13192 -14892
rect 13270 -14602 13330 -14542
rect 13590 -14602 13650 -14542
rect 13270 -14952 13330 -14892
rect 13590 -14952 13650 -14892
rect 13726 -14602 13786 -14542
rect 14046 -14602 14106 -14542
rect 14182 -14602 14242 -14542
rect 14502 -14602 14562 -14542
rect 14640 -14602 14700 -14542
rect 14960 -14602 15020 -14542
rect 15096 -14602 15156 -14542
rect 15416 -14602 15476 -14542
rect 13726 -14952 13786 -14892
rect 14046 -14952 14106 -14892
rect 14182 -14952 14242 -14892
rect 14502 -14952 14562 -14892
rect 14640 -14952 14700 -14892
rect 14960 -14952 15020 -14892
rect 15096 -14952 15156 -14892
rect 15416 -14952 15476 -14892
rect 10 -15094 14 -15034
rect 14 -15094 66 -15034
rect 66 -15094 70 -15034
rect 330 -15094 390 -15034
rect 10 -15444 14 -15384
rect 14 -15444 66 -15384
rect 66 -15444 70 -15384
rect 330 -15444 390 -15384
rect 466 -15094 526 -15034
rect 786 -15094 846 -15034
rect 922 -15094 982 -15034
rect 1242 -15094 1302 -15034
rect 1380 -15094 1440 -15034
rect 1700 -15094 1760 -15034
rect 1836 -15094 1896 -15034
rect 2156 -15094 2216 -15034
rect 2292 -15094 2352 -15034
rect 2612 -15094 2672 -15034
rect 2750 -15094 2810 -15034
rect 3070 -15094 3130 -15034
rect 3206 -15094 3266 -15034
rect 3526 -15094 3586 -15034
rect 466 -15444 526 -15384
rect 786 -15444 846 -15384
rect 922 -15444 982 -15384
rect 1242 -15444 1302 -15384
rect 1380 -15444 1440 -15384
rect 1700 -15444 1760 -15384
rect 1836 -15444 1896 -15384
rect 2156 -15444 2216 -15384
rect 2292 -15444 2352 -15384
rect 2612 -15444 2672 -15384
rect 2750 -15444 2810 -15384
rect 3070 -15444 3130 -15384
rect 3206 -15444 3266 -15384
rect 3526 -15444 3586 -15384
rect 3662 -15094 3722 -15034
rect 3982 -15094 4042 -15034
rect 4120 -15094 4180 -15034
rect 4440 -15094 4500 -15034
rect 4576 -15094 4636 -15034
rect 4896 -15094 4956 -15034
rect 5032 -15094 5092 -15034
rect 5352 -15094 5412 -15034
rect 5490 -15094 5550 -15034
rect 5810 -15094 5870 -15034
rect 5946 -15094 6006 -15034
rect 6266 -15094 6326 -15034
rect 6402 -15094 6462 -15034
rect 6722 -15094 6782 -15034
rect 6860 -15094 6920 -15034
rect 7180 -15094 7240 -15034
rect 3662 -15444 3722 -15384
rect 3982 -15444 4042 -15384
rect 4120 -15444 4180 -15384
rect 4440 -15444 4500 -15384
rect 4576 -15444 4636 -15384
rect 4896 -15444 4956 -15384
rect 5032 -15444 5092 -15384
rect 5352 -15444 5412 -15384
rect 5490 -15444 5550 -15384
rect 5810 -15444 5870 -15384
rect 5946 -15444 6006 -15384
rect 6266 -15444 6326 -15384
rect 6402 -15444 6462 -15384
rect 6722 -15444 6782 -15384
rect 6860 -15444 6920 -15384
rect 7180 -15444 7240 -15384
rect 7316 -15094 7376 -15034
rect 7636 -15094 7696 -15034
rect 7772 -15094 7832 -15034
rect 8092 -15094 8152 -15034
rect 8246 -15094 8306 -15034
rect 8566 -15094 8626 -15034
rect 8702 -15094 8762 -15034
rect 9022 -15094 9082 -15034
rect 9160 -15094 9220 -15034
rect 9480 -15094 9540 -15034
rect 9616 -15094 9676 -15034
rect 9936 -15094 9996 -15034
rect 10072 -15094 10132 -15034
rect 10392 -15094 10452 -15034
rect 10530 -15094 10590 -15034
rect 10850 -15094 10910 -15034
rect 7316 -15444 7376 -15384
rect 7636 -15444 7696 -15384
rect 7772 -15444 7832 -15384
rect 8092 -15444 8152 -15384
rect 8246 -15444 8306 -15384
rect 8566 -15444 8626 -15384
rect 8702 -15444 8762 -15384
rect 9022 -15444 9082 -15384
rect 9160 -15444 9220 -15384
rect 9480 -15444 9540 -15384
rect 9616 -15444 9676 -15384
rect 9936 -15444 9996 -15384
rect 10072 -15444 10132 -15384
rect 10392 -15444 10452 -15384
rect 10530 -15444 10590 -15384
rect 10850 -15444 10910 -15384
rect 10986 -15094 11046 -15034
rect 11306 -15094 11366 -15034
rect 11442 -15094 11502 -15034
rect 11762 -15094 11822 -15034
rect 10986 -15444 11046 -15384
rect 11306 -15444 11366 -15384
rect 11442 -15444 11502 -15384
rect 11762 -15444 11822 -15384
rect 11900 -15094 11960 -15034
rect 12220 -15094 12280 -15034
rect 12356 -15094 12416 -15034
rect 12676 -15094 12736 -15034
rect 12812 -15094 12872 -15034
rect 13132 -15094 13192 -15034
rect 11900 -15444 11960 -15384
rect 12220 -15444 12280 -15384
rect 12356 -15444 12416 -15384
rect 12676 -15444 12736 -15384
rect 12812 -15444 12872 -15384
rect 13132 -15444 13192 -15384
rect 13270 -15094 13330 -15034
rect 13590 -15094 13650 -15034
rect 13270 -15444 13330 -15384
rect 13590 -15444 13650 -15384
rect 13726 -15094 13786 -15034
rect 14046 -15094 14106 -15034
rect 13726 -15444 13786 -15384
rect 14046 -15444 14106 -15384
rect 14182 -15094 14242 -15034
rect 14502 -15094 14562 -15034
rect 14640 -15094 14700 -15034
rect 14960 -15094 15020 -15034
rect 15096 -15094 15156 -15034
rect 15416 -15094 15476 -15034
rect 14182 -15444 14242 -15384
rect 14502 -15444 14562 -15384
rect 14640 -15444 14700 -15384
rect 14960 -15444 15020 -15384
rect 15096 -15444 15156 -15384
rect 15416 -15444 15476 -15384
rect 10 -15610 14 -15550
rect 14 -15610 66 -15550
rect 66 -15610 70 -15550
rect 330 -15610 390 -15550
rect 10 -15960 14 -15900
rect 14 -15960 66 -15900
rect 66 -15960 70 -15900
rect 330 -15960 390 -15900
rect 466 -15610 526 -15550
rect 786 -15610 846 -15550
rect 922 -15610 982 -15550
rect 1242 -15610 1302 -15550
rect 1380 -15610 1440 -15550
rect 1700 -15610 1760 -15550
rect 1836 -15610 1896 -15550
rect 2156 -15610 2216 -15550
rect 2292 -15610 2352 -15550
rect 2612 -15610 2672 -15550
rect 2750 -15610 2810 -15550
rect 3070 -15610 3130 -15550
rect 3206 -15610 3266 -15550
rect 3526 -15610 3586 -15550
rect 466 -15960 526 -15900
rect 786 -15960 846 -15900
rect 922 -15960 982 -15900
rect 1242 -15960 1302 -15900
rect 1380 -15960 1440 -15900
rect 1700 -15960 1760 -15900
rect 1836 -15960 1896 -15900
rect 2156 -15960 2216 -15900
rect 2292 -15960 2352 -15900
rect 2612 -15960 2672 -15900
rect 2750 -15960 2810 -15900
rect 3070 -15960 3130 -15900
rect 3206 -15960 3266 -15900
rect 3526 -15960 3586 -15900
rect 3662 -15610 3722 -15550
rect 3982 -15610 4042 -15550
rect 4120 -15610 4180 -15550
rect 4440 -15610 4500 -15550
rect 4576 -15610 4636 -15550
rect 4896 -15610 4956 -15550
rect 5032 -15610 5092 -15550
rect 5352 -15610 5412 -15550
rect 5490 -15610 5550 -15550
rect 5810 -15610 5870 -15550
rect 5946 -15610 6006 -15550
rect 6266 -15610 6326 -15550
rect 6402 -15610 6462 -15550
rect 6722 -15610 6782 -15550
rect 3662 -15960 3722 -15900
rect 3982 -15960 4042 -15900
rect 4120 -15960 4180 -15900
rect 4440 -15960 4500 -15900
rect 4576 -15960 4636 -15900
rect 4896 -15960 4956 -15900
rect 5032 -15960 5092 -15900
rect 5352 -15960 5412 -15900
rect 5490 -15960 5550 -15900
rect 5810 -15960 5870 -15900
rect 5946 -15960 6006 -15900
rect 6266 -15960 6326 -15900
rect 6402 -15960 6462 -15900
rect 6722 -15960 6782 -15900
rect 6860 -15610 6920 -15550
rect 7180 -15610 7240 -15550
rect 7316 -15610 7376 -15550
rect 7636 -15610 7696 -15550
rect 7772 -15610 7832 -15550
rect 8092 -15610 8152 -15550
rect 8246 -15610 8306 -15550
rect 8566 -15610 8626 -15550
rect 8702 -15610 8762 -15550
rect 9022 -15610 9082 -15550
rect 9160 -15610 9220 -15550
rect 9480 -15610 9540 -15550
rect 9616 -15610 9676 -15550
rect 9936 -15610 9996 -15550
rect 10072 -15610 10132 -15550
rect 10392 -15610 10452 -15550
rect 6860 -15960 6920 -15900
rect 7180 -15960 7240 -15900
rect 7316 -15960 7376 -15900
rect 7636 -15960 7696 -15900
rect 7772 -15960 7832 -15900
rect 8092 -15960 8152 -15900
rect 8246 -15960 8306 -15900
rect 8566 -15960 8626 -15900
rect 8702 -15960 8762 -15900
rect 9022 -15960 9082 -15900
rect 9160 -15960 9220 -15900
rect 9480 -15960 9540 -15900
rect 9616 -15960 9676 -15900
rect 9936 -15960 9996 -15900
rect 10072 -15960 10132 -15900
rect 10392 -15960 10452 -15900
rect 10530 -15610 10590 -15550
rect 10850 -15610 10910 -15550
rect 10986 -15610 11046 -15550
rect 11306 -15610 11366 -15550
rect 11442 -15610 11502 -15550
rect 11762 -15610 11822 -15550
rect 10530 -15960 10590 -15900
rect 10850 -15960 10910 -15900
rect 10986 -15960 11046 -15900
rect 11306 -15960 11366 -15900
rect 11442 -15960 11502 -15900
rect 11762 -15960 11822 -15900
rect 11900 -15610 11960 -15550
rect 12220 -15610 12280 -15550
rect 12356 -15610 12416 -15550
rect 12676 -15610 12736 -15550
rect 12812 -15610 12872 -15550
rect 13132 -15610 13192 -15550
rect 11900 -15960 11960 -15900
rect 12220 -15960 12280 -15900
rect 12356 -15960 12416 -15900
rect 12676 -15960 12736 -15900
rect 12812 -15960 12872 -15900
rect 13132 -15960 13192 -15900
rect 13270 -15610 13330 -15550
rect 13590 -15610 13650 -15550
rect 13270 -15960 13330 -15900
rect 13590 -15960 13650 -15900
rect 13726 -15610 13786 -15550
rect 14046 -15610 14106 -15550
rect 13726 -15960 13786 -15900
rect 14046 -15960 14106 -15900
rect 14182 -15610 14242 -15550
rect 14502 -15610 14562 -15550
rect 14182 -15960 14242 -15900
rect 14502 -15960 14562 -15900
rect 14640 -15610 14700 -15550
rect 14960 -15610 15020 -15550
rect 15096 -15610 15156 -15550
rect 15416 -15610 15476 -15550
rect 14640 -15960 14700 -15900
rect 14960 -15960 15020 -15900
rect 15096 -15960 15156 -15900
rect 15416 -15960 15476 -15900
rect 10 -16112 14 -16052
rect 14 -16112 66 -16052
rect 66 -16112 70 -16052
rect 330 -16112 390 -16052
rect 10 -16462 14 -16402
rect 14 -16462 66 -16402
rect 66 -16462 70 -16402
rect 330 -16462 390 -16402
rect 466 -16112 526 -16052
rect 786 -16112 846 -16052
rect 922 -16112 982 -16052
rect 1242 -16112 1302 -16052
rect 1380 -16112 1440 -16052
rect 1700 -16112 1760 -16052
rect 1836 -16112 1896 -16052
rect 2156 -16112 2216 -16052
rect 2292 -16112 2352 -16052
rect 2612 -16112 2672 -16052
rect 2750 -16112 2810 -16052
rect 3070 -16112 3130 -16052
rect 3206 -16112 3266 -16052
rect 3526 -16112 3586 -16052
rect 466 -16462 526 -16402
rect 786 -16462 846 -16402
rect 922 -16462 982 -16402
rect 1242 -16462 1302 -16402
rect 1380 -16462 1440 -16402
rect 1700 -16462 1760 -16402
rect 1836 -16462 1896 -16402
rect 2156 -16462 2216 -16402
rect 2292 -16462 2352 -16402
rect 2612 -16462 2672 -16402
rect 2750 -16462 2810 -16402
rect 3070 -16462 3130 -16402
rect 3206 -16462 3266 -16402
rect 3526 -16462 3586 -16402
rect 3662 -16112 3722 -16052
rect 3982 -16112 4042 -16052
rect 4120 -16112 4180 -16052
rect 4440 -16112 4500 -16052
rect 4576 -16112 4636 -16052
rect 4896 -16112 4956 -16052
rect 5032 -16112 5092 -16052
rect 5352 -16112 5412 -16052
rect 5490 -16112 5550 -16052
rect 5810 -16112 5870 -16052
rect 5946 -16112 6006 -16052
rect 6266 -16112 6326 -16052
rect 6402 -16112 6462 -16052
rect 6722 -16112 6782 -16052
rect 3662 -16462 3722 -16402
rect 3982 -16462 4042 -16402
rect 4120 -16462 4180 -16402
rect 4440 -16462 4500 -16402
rect 4576 -16462 4636 -16402
rect 4896 -16462 4956 -16402
rect 5032 -16462 5092 -16402
rect 5352 -16462 5412 -16402
rect 5490 -16462 5550 -16402
rect 5810 -16462 5870 -16402
rect 5946 -16462 6006 -16402
rect 6266 -16462 6326 -16402
rect 6402 -16462 6462 -16402
rect 6722 -16462 6782 -16402
rect 6860 -16112 6920 -16052
rect 7180 -16112 7240 -16052
rect 7316 -16112 7376 -16052
rect 7636 -16112 7696 -16052
rect 7772 -16112 7832 -16052
rect 8092 -16112 8152 -16052
rect 8246 -16112 8306 -16052
rect 8566 -16112 8626 -16052
rect 8702 -16112 8762 -16052
rect 9022 -16112 9082 -16052
rect 9160 -16112 9220 -16052
rect 9480 -16112 9540 -16052
rect 9616 -16112 9676 -16052
rect 9936 -16112 9996 -16052
rect 10072 -16112 10132 -16052
rect 10392 -16112 10452 -16052
rect 6860 -16462 6920 -16402
rect 7180 -16462 7240 -16402
rect 7316 -16462 7376 -16402
rect 7636 -16462 7696 -16402
rect 7772 -16462 7832 -16402
rect 8092 -16462 8152 -16402
rect 8246 -16462 8306 -16402
rect 8566 -16462 8626 -16402
rect 8702 -16462 8762 -16402
rect 9022 -16462 9082 -16402
rect 9160 -16462 9220 -16402
rect 9480 -16462 9540 -16402
rect 9616 -16462 9676 -16402
rect 9936 -16462 9996 -16402
rect 10072 -16462 10132 -16402
rect 10392 -16462 10452 -16402
rect 10530 -16112 10590 -16052
rect 10850 -16112 10910 -16052
rect 10986 -16112 11046 -16052
rect 11306 -16112 11366 -16052
rect 11442 -16112 11502 -16052
rect 11762 -16112 11822 -16052
rect 10530 -16462 10590 -16402
rect 10850 -16462 10910 -16402
rect 10986 -16462 11046 -16402
rect 11306 -16462 11366 -16402
rect 11442 -16462 11502 -16402
rect 11762 -16462 11822 -16402
rect 11900 -16112 11960 -16052
rect 12220 -16112 12280 -16052
rect 12356 -16112 12416 -16052
rect 12676 -16112 12736 -16052
rect 12812 -16112 12872 -16052
rect 13132 -16112 13192 -16052
rect 11900 -16462 11960 -16402
rect 12220 -16462 12280 -16402
rect 12356 -16462 12416 -16402
rect 12676 -16462 12736 -16402
rect 12812 -16462 12872 -16402
rect 13132 -16462 13192 -16402
rect 13270 -16112 13330 -16052
rect 13590 -16112 13650 -16052
rect 13270 -16462 13330 -16402
rect 13590 -16462 13650 -16402
rect 13726 -16112 13786 -16052
rect 14046 -16112 14106 -16052
rect 13726 -16462 13786 -16402
rect 14046 -16462 14106 -16402
rect 14182 -16112 14242 -16052
rect 14502 -16112 14562 -16052
rect 14182 -16462 14242 -16402
rect 14502 -16462 14562 -16402
rect 14640 -16112 14700 -16052
rect 14960 -16112 15020 -16052
rect 15096 -16112 15156 -16052
rect 15416 -16112 15476 -16052
rect 14640 -16462 14700 -16402
rect 14960 -16462 15020 -16402
rect 15096 -16462 15156 -16402
rect 15416 -16462 15476 -16402
rect 10 -16604 14 -16544
rect 14 -16604 66 -16544
rect 66 -16604 70 -16544
rect 330 -16604 390 -16544
rect 10 -16954 14 -16894
rect 14 -16954 66 -16894
rect 66 -16954 70 -16894
rect 330 -16954 390 -16894
rect 466 -16604 526 -16544
rect 786 -16604 846 -16544
rect 922 -16604 982 -16544
rect 1242 -16604 1302 -16544
rect 1380 -16604 1440 -16544
rect 1700 -16604 1760 -16544
rect 1836 -16604 1896 -16544
rect 2156 -16604 2216 -16544
rect 2292 -16604 2352 -16544
rect 2612 -16604 2672 -16544
rect 2750 -16604 2810 -16544
rect 3070 -16604 3130 -16544
rect 3206 -16604 3266 -16544
rect 3526 -16604 3586 -16544
rect 466 -16954 526 -16894
rect 786 -16954 846 -16894
rect 922 -16954 982 -16894
rect 1242 -16954 1302 -16894
rect 1380 -16954 1440 -16894
rect 1700 -16954 1760 -16894
rect 1836 -16954 1896 -16894
rect 2156 -16954 2216 -16894
rect 2292 -16954 2352 -16894
rect 2612 -16954 2672 -16894
rect 2750 -16954 2810 -16894
rect 3070 -16954 3130 -16894
rect 3206 -16954 3266 -16894
rect 3526 -16954 3586 -16894
rect 3662 -16604 3722 -16544
rect 3982 -16604 4042 -16544
rect 4120 -16604 4180 -16544
rect 4440 -16604 4500 -16544
rect 4576 -16604 4636 -16544
rect 4896 -16604 4956 -16544
rect 5032 -16604 5092 -16544
rect 5352 -16604 5412 -16544
rect 5490 -16604 5550 -16544
rect 5810 -16604 5870 -16544
rect 5946 -16604 6006 -16544
rect 6266 -16604 6326 -16544
rect 6402 -16604 6462 -16544
rect 6722 -16604 6782 -16544
rect 6860 -16604 6920 -16544
rect 7180 -16604 7240 -16544
rect 3662 -16954 3722 -16894
rect 3982 -16954 4042 -16894
rect 4120 -16954 4180 -16894
rect 4440 -16954 4500 -16894
rect 4576 -16954 4636 -16894
rect 4896 -16954 4956 -16894
rect 5032 -16954 5092 -16894
rect 5352 -16954 5412 -16894
rect 5490 -16954 5550 -16894
rect 5810 -16954 5870 -16894
rect 5946 -16954 6006 -16894
rect 6266 -16954 6326 -16894
rect 6402 -16954 6462 -16894
rect 6722 -16954 6782 -16894
rect 6860 -16954 6920 -16894
rect 7180 -16954 7240 -16894
rect 7316 -16604 7376 -16544
rect 7636 -16604 7696 -16544
rect 7772 -16604 7832 -16544
rect 8092 -16604 8152 -16544
rect 8246 -16604 8306 -16544
rect 8566 -16604 8626 -16544
rect 8702 -16604 8762 -16544
rect 9022 -16604 9082 -16544
rect 9160 -16604 9220 -16544
rect 9480 -16604 9540 -16544
rect 9616 -16604 9676 -16544
rect 9936 -16604 9996 -16544
rect 10072 -16604 10132 -16544
rect 10392 -16604 10452 -16544
rect 10530 -16604 10590 -16544
rect 10850 -16604 10910 -16544
rect 7316 -16954 7376 -16894
rect 7636 -16954 7696 -16894
rect 7772 -16954 7832 -16894
rect 8092 -16954 8152 -16894
rect 8246 -16954 8306 -16894
rect 8566 -16954 8626 -16894
rect 8702 -16954 8762 -16894
rect 9022 -16954 9082 -16894
rect 9160 -16954 9220 -16894
rect 9480 -16954 9540 -16894
rect 9616 -16954 9676 -16894
rect 9936 -16954 9996 -16894
rect 10072 -16954 10132 -16894
rect 10392 -16954 10452 -16894
rect 10530 -16954 10590 -16894
rect 10850 -16954 10910 -16894
rect 10986 -16604 11046 -16544
rect 11306 -16604 11366 -16544
rect 11442 -16604 11502 -16544
rect 11762 -16604 11822 -16544
rect 10986 -16954 11046 -16894
rect 11306 -16954 11366 -16894
rect 11442 -16954 11502 -16894
rect 11762 -16954 11822 -16894
rect 11900 -16604 11960 -16544
rect 12220 -16604 12280 -16544
rect 12356 -16604 12416 -16544
rect 12676 -16604 12736 -16544
rect 12812 -16604 12872 -16544
rect 13132 -16604 13192 -16544
rect 11900 -16954 11960 -16894
rect 12220 -16954 12280 -16894
rect 12356 -16954 12416 -16894
rect 12676 -16954 12736 -16894
rect 12812 -16954 12872 -16894
rect 13132 -16954 13192 -16894
rect 13270 -16604 13330 -16544
rect 13590 -16604 13650 -16544
rect 13270 -16954 13330 -16894
rect 13590 -16954 13650 -16894
rect 13726 -16604 13786 -16544
rect 14046 -16604 14106 -16544
rect 13726 -16954 13786 -16894
rect 14046 -16954 14106 -16894
rect 14182 -16604 14242 -16544
rect 14502 -16604 14562 -16544
rect 14640 -16604 14700 -16544
rect 14960 -16604 15020 -16544
rect 15096 -16604 15156 -16544
rect 15416 -16604 15476 -16544
rect 14182 -16954 14242 -16894
rect 14502 -16954 14562 -16894
rect 14640 -16954 14700 -16894
rect 14960 -16954 15020 -16894
rect 15096 -16954 15156 -16894
rect 15416 -16954 15476 -16894
rect 11 -17101 14 -17041
rect 14 -17101 66 -17041
rect 66 -17101 71 -17041
rect 331 -17101 391 -17041
rect 11 -17451 14 -17391
rect 14 -17451 66 -17391
rect 66 -17451 71 -17391
rect 331 -17451 391 -17391
rect 467 -17101 527 -17041
rect 787 -17101 847 -17041
rect 923 -17101 983 -17041
rect 1243 -17101 1303 -17041
rect 1381 -17101 1441 -17041
rect 1701 -17101 1761 -17041
rect 1837 -17101 1897 -17041
rect 2157 -17101 2217 -17041
rect 2293 -17101 2353 -17041
rect 2613 -17101 2673 -17041
rect 2751 -17101 2811 -17041
rect 3071 -17101 3131 -17041
rect 3207 -17101 3267 -17041
rect 3527 -17101 3587 -17041
rect 467 -17451 527 -17391
rect 787 -17451 847 -17391
rect 923 -17451 983 -17391
rect 1243 -17451 1303 -17391
rect 1381 -17451 1441 -17391
rect 1701 -17451 1761 -17391
rect 1837 -17451 1897 -17391
rect 2157 -17451 2217 -17391
rect 2293 -17451 2353 -17391
rect 2613 -17451 2673 -17391
rect 2751 -17451 2811 -17391
rect 3071 -17451 3131 -17391
rect 3207 -17451 3267 -17391
rect 3527 -17451 3587 -17391
rect 3663 -17101 3723 -17041
rect 3983 -17101 4043 -17041
rect 4121 -17101 4181 -17041
rect 4441 -17101 4501 -17041
rect 4577 -17101 4637 -17041
rect 4897 -17101 4957 -17041
rect 5033 -17101 5093 -17041
rect 5353 -17101 5413 -17041
rect 5491 -17101 5551 -17041
rect 5811 -17101 5871 -17041
rect 5947 -17101 6007 -17041
rect 6267 -17101 6327 -17041
rect 6403 -17101 6463 -17041
rect 6723 -17101 6783 -17041
rect 6861 -17101 6921 -17041
rect 7181 -17101 7241 -17041
rect 3663 -17451 3723 -17391
rect 3983 -17451 4043 -17391
rect 4121 -17451 4181 -17391
rect 4441 -17451 4501 -17391
rect 4577 -17451 4637 -17391
rect 4897 -17451 4957 -17391
rect 5033 -17451 5093 -17391
rect 5353 -17451 5413 -17391
rect 5491 -17451 5551 -17391
rect 5811 -17451 5871 -17391
rect 5947 -17451 6007 -17391
rect 6267 -17451 6327 -17391
rect 6403 -17451 6463 -17391
rect 6723 -17451 6783 -17391
rect 6861 -17451 6921 -17391
rect 7181 -17451 7241 -17391
rect 7317 -17101 7377 -17041
rect 7637 -17101 7697 -17041
rect 7773 -17101 7833 -17041
rect 8093 -17101 8153 -17041
rect 8247 -17101 8307 -17041
rect 8567 -17101 8627 -17041
rect 8703 -17101 8763 -17041
rect 9023 -17101 9083 -17041
rect 9161 -17101 9221 -17041
rect 9481 -17101 9541 -17041
rect 9617 -17101 9677 -17041
rect 9937 -17101 9997 -17041
rect 10073 -17101 10133 -17041
rect 10393 -17101 10453 -17041
rect 10531 -17101 10591 -17041
rect 10851 -17101 10911 -17041
rect 7317 -17451 7377 -17391
rect 7637 -17451 7697 -17391
rect 7773 -17451 7833 -17391
rect 8093 -17451 8153 -17391
rect 8247 -17451 8307 -17391
rect 8567 -17451 8627 -17391
rect 8703 -17451 8763 -17391
rect 9023 -17451 9083 -17391
rect 9161 -17451 9221 -17391
rect 9481 -17451 9541 -17391
rect 9617 -17451 9677 -17391
rect 9937 -17451 9997 -17391
rect 10073 -17451 10133 -17391
rect 10393 -17451 10453 -17391
rect 10531 -17451 10591 -17391
rect 10851 -17451 10911 -17391
rect 10987 -17101 11047 -17041
rect 11307 -17101 11367 -17041
rect 11443 -17101 11503 -17041
rect 11763 -17101 11823 -17041
rect 11901 -17101 11961 -17041
rect 12221 -17101 12281 -17041
rect 10987 -17451 11047 -17391
rect 11307 -17451 11367 -17391
rect 11443 -17451 11503 -17391
rect 11763 -17451 11823 -17391
rect 11901 -17451 11961 -17391
rect 12221 -17451 12281 -17391
rect 12357 -17101 12417 -17041
rect 12677 -17101 12737 -17041
rect 12813 -17101 12873 -17041
rect 13133 -17101 13193 -17041
rect 12357 -17451 12417 -17391
rect 12677 -17451 12737 -17391
rect 12813 -17451 12873 -17391
rect 13133 -17451 13193 -17391
rect 13271 -17101 13331 -17041
rect 13591 -17101 13651 -17041
rect 13271 -17451 13331 -17391
rect 13591 -17451 13651 -17391
rect 13727 -17101 13787 -17041
rect 14047 -17101 14107 -17041
rect 13727 -17451 13787 -17391
rect 14047 -17451 14107 -17391
rect 14183 -17101 14243 -17041
rect 14503 -17101 14563 -17041
rect 14641 -17101 14701 -17041
rect 14961 -17101 15021 -17041
rect 15097 -17101 15157 -17041
rect 15417 -17101 15477 -17041
rect 14183 -17451 14243 -17391
rect 14503 -17451 14563 -17391
rect 14641 -17451 14701 -17391
rect 14961 -17451 15021 -17391
rect 15097 -17451 15157 -17391
rect 15417 -17451 15477 -17391
rect 11 -17593 14 -17533
rect 14 -17593 66 -17533
rect 66 -17593 71 -17533
rect 331 -17593 391 -17533
rect 11 -17943 14 -17883
rect 14 -17943 66 -17883
rect 66 -17943 71 -17883
rect 331 -17943 391 -17883
rect 467 -17593 527 -17533
rect 787 -17593 847 -17533
rect 923 -17593 983 -17533
rect 1243 -17593 1303 -17533
rect 1381 -17593 1441 -17533
rect 1701 -17593 1761 -17533
rect 1837 -17593 1897 -17533
rect 2157 -17593 2217 -17533
rect 2293 -17593 2353 -17533
rect 2613 -17593 2673 -17533
rect 2751 -17593 2811 -17533
rect 3071 -17593 3131 -17533
rect 3207 -17593 3267 -17533
rect 3527 -17593 3587 -17533
rect 467 -17943 527 -17883
rect 787 -17943 847 -17883
rect 923 -17943 983 -17883
rect 1243 -17943 1303 -17883
rect 1381 -17943 1441 -17883
rect 1701 -17943 1761 -17883
rect 1837 -17943 1897 -17883
rect 2157 -17943 2217 -17883
rect 2293 -17943 2353 -17883
rect 2613 -17943 2673 -17883
rect 2751 -17943 2811 -17883
rect 3071 -17943 3131 -17883
rect 3207 -17943 3267 -17883
rect 3527 -17943 3587 -17883
rect 3663 -17593 3723 -17533
rect 3983 -17593 4043 -17533
rect 4121 -17593 4181 -17533
rect 4441 -17593 4501 -17533
rect 4577 -17593 4637 -17533
rect 4897 -17593 4957 -17533
rect 5033 -17593 5093 -17533
rect 5353 -17593 5413 -17533
rect 5491 -17593 5551 -17533
rect 5811 -17593 5871 -17533
rect 5947 -17593 6007 -17533
rect 6267 -17593 6327 -17533
rect 6403 -17593 6463 -17533
rect 6723 -17593 6783 -17533
rect 6861 -17593 6921 -17533
rect 7181 -17593 7241 -17533
rect 3663 -17943 3723 -17883
rect 3983 -17943 4043 -17883
rect 4121 -17943 4181 -17883
rect 4441 -17943 4501 -17883
rect 4577 -17943 4637 -17883
rect 4897 -17943 4957 -17883
rect 5033 -17943 5093 -17883
rect 5353 -17943 5413 -17883
rect 5491 -17943 5551 -17883
rect 5811 -17943 5871 -17883
rect 5947 -17943 6007 -17883
rect 6267 -17943 6327 -17883
rect 6403 -17943 6463 -17883
rect 6723 -17943 6783 -17883
rect 6861 -17943 6921 -17883
rect 7181 -17943 7241 -17883
rect 7317 -17593 7377 -17533
rect 7637 -17593 7697 -17533
rect 7773 -17593 7833 -17533
rect 8093 -17593 8153 -17533
rect 8247 -17593 8307 -17533
rect 8567 -17593 8627 -17533
rect 8703 -17593 8763 -17533
rect 9023 -17593 9083 -17533
rect 9161 -17593 9221 -17533
rect 9481 -17593 9541 -17533
rect 9617 -17593 9677 -17533
rect 9937 -17593 9997 -17533
rect 10073 -17593 10133 -17533
rect 10393 -17593 10453 -17533
rect 10531 -17593 10591 -17533
rect 10851 -17593 10911 -17533
rect 7317 -17943 7377 -17883
rect 7637 -17943 7697 -17883
rect 7773 -17943 7833 -17883
rect 8093 -17943 8153 -17883
rect 8247 -17943 8307 -17883
rect 8567 -17943 8627 -17883
rect 8703 -17943 8763 -17883
rect 9023 -17943 9083 -17883
rect 9161 -17943 9221 -17883
rect 9481 -17943 9541 -17883
rect 9617 -17943 9677 -17883
rect 9937 -17943 9997 -17883
rect 10073 -17943 10133 -17883
rect 10393 -17943 10453 -17883
rect 10531 -17943 10591 -17883
rect 10851 -17943 10911 -17883
rect 10987 -17593 11047 -17533
rect 11307 -17593 11367 -17533
rect 11443 -17593 11503 -17533
rect 11763 -17593 11823 -17533
rect 11901 -17593 11961 -17533
rect 12221 -17593 12281 -17533
rect 10987 -17943 11047 -17883
rect 11307 -17943 11367 -17883
rect 11443 -17943 11503 -17883
rect 11763 -17943 11823 -17883
rect 11901 -17943 11961 -17883
rect 12221 -17943 12281 -17883
rect 12357 -17593 12417 -17533
rect 12677 -17593 12737 -17533
rect 12813 -17593 12873 -17533
rect 13133 -17593 13193 -17533
rect 12357 -17943 12417 -17883
rect 12677 -17943 12737 -17883
rect 12813 -17943 12873 -17883
rect 13133 -17943 13193 -17883
rect 13271 -17593 13331 -17533
rect 13591 -17593 13651 -17533
rect 13727 -17593 13787 -17533
rect 14047 -17593 14107 -17533
rect 14183 -17593 14243 -17533
rect 14503 -17593 14563 -17533
rect 14641 -17593 14701 -17533
rect 14961 -17593 15021 -17533
rect 15097 -17593 15157 -17533
rect 15417 -17593 15477 -17533
rect 13271 -17943 13331 -17883
rect 13591 -17943 13651 -17883
rect 13727 -17943 13787 -17883
rect 14047 -17943 14107 -17883
rect 14183 -17943 14243 -17883
rect 14503 -17943 14563 -17883
rect 14641 -17943 14701 -17883
rect 14961 -17943 15021 -17883
rect 15097 -17943 15157 -17883
rect 15417 -17943 15477 -17883
rect 11 -18109 14 -18049
rect 14 -18109 66 -18049
rect 66 -18109 71 -18049
rect 331 -18109 391 -18049
rect 11 -18459 14 -18399
rect 14 -18459 66 -18399
rect 66 -18459 71 -18399
rect 331 -18459 391 -18399
rect 467 -18109 527 -18049
rect 787 -18109 847 -18049
rect 923 -18109 983 -18049
rect 1243 -18109 1303 -18049
rect 1381 -18109 1441 -18049
rect 1701 -18109 1761 -18049
rect 1837 -18109 1897 -18049
rect 2157 -18109 2217 -18049
rect 2293 -18109 2353 -18049
rect 2613 -18109 2673 -18049
rect 2751 -18109 2811 -18049
rect 3071 -18109 3131 -18049
rect 3207 -18109 3267 -18049
rect 3527 -18109 3587 -18049
rect 467 -18459 527 -18399
rect 787 -18459 847 -18399
rect 923 -18459 983 -18399
rect 1243 -18459 1303 -18399
rect 1381 -18459 1441 -18399
rect 1701 -18459 1761 -18399
rect 1837 -18459 1897 -18399
rect 2157 -18459 2217 -18399
rect 2293 -18459 2353 -18399
rect 2613 -18459 2673 -18399
rect 2751 -18459 2811 -18399
rect 3071 -18459 3131 -18399
rect 3207 -18459 3267 -18399
rect 3527 -18459 3587 -18399
rect 3663 -18109 3723 -18049
rect 3983 -18109 4043 -18049
rect 4121 -18109 4181 -18049
rect 4441 -18109 4501 -18049
rect 4577 -18109 4637 -18049
rect 4897 -18109 4957 -18049
rect 5033 -18109 5093 -18049
rect 5353 -18109 5413 -18049
rect 5491 -18109 5551 -18049
rect 5811 -18109 5871 -18049
rect 5947 -18109 6007 -18049
rect 6267 -18109 6327 -18049
rect 6403 -18109 6463 -18049
rect 6723 -18109 6783 -18049
rect 6861 -18109 6921 -18049
rect 7181 -18109 7241 -18049
rect 3663 -18459 3723 -18399
rect 3983 -18459 4043 -18399
rect 4121 -18459 4181 -18399
rect 4441 -18459 4501 -18399
rect 4577 -18459 4637 -18399
rect 4897 -18459 4957 -18399
rect 5033 -18459 5093 -18399
rect 5353 -18459 5413 -18399
rect 5491 -18459 5551 -18399
rect 5811 -18459 5871 -18399
rect 5947 -18459 6007 -18399
rect 6267 -18459 6327 -18399
rect 6403 -18459 6463 -18399
rect 6723 -18459 6783 -18399
rect 6861 -18459 6921 -18399
rect 7181 -18459 7241 -18399
rect 7317 -18109 7377 -18049
rect 7637 -18109 7697 -18049
rect 7773 -18109 7833 -18049
rect 8093 -18109 8153 -18049
rect 8247 -18109 8307 -18049
rect 8567 -18109 8627 -18049
rect 8703 -18109 8763 -18049
rect 9023 -18109 9083 -18049
rect 9161 -18109 9221 -18049
rect 9481 -18109 9541 -18049
rect 9617 -18109 9677 -18049
rect 9937 -18109 9997 -18049
rect 10073 -18109 10133 -18049
rect 10393 -18109 10453 -18049
rect 10531 -18109 10591 -18049
rect 10851 -18109 10911 -18049
rect 7317 -18459 7377 -18399
rect 7637 -18459 7697 -18399
rect 7773 -18459 7833 -18399
rect 8093 -18459 8153 -18399
rect 8247 -18459 8307 -18399
rect 8567 -18459 8627 -18399
rect 8703 -18459 8763 -18399
rect 9023 -18459 9083 -18399
rect 9161 -18459 9221 -18399
rect 9481 -18459 9541 -18399
rect 9617 -18459 9677 -18399
rect 9937 -18459 9997 -18399
rect 10073 -18459 10133 -18399
rect 10393 -18459 10453 -18399
rect 10531 -18459 10591 -18399
rect 10851 -18459 10911 -18399
rect 10987 -18109 11047 -18049
rect 11307 -18109 11367 -18049
rect 11443 -18109 11503 -18049
rect 11763 -18109 11823 -18049
rect 11901 -18109 11961 -18049
rect 12221 -18109 12281 -18049
rect 10987 -18459 11047 -18399
rect 11307 -18459 11367 -18399
rect 11443 -18459 11503 -18399
rect 11763 -18459 11823 -18399
rect 11901 -18459 11961 -18399
rect 12221 -18459 12281 -18399
rect 12357 -18109 12417 -18049
rect 12677 -18109 12737 -18049
rect 12813 -18109 12873 -18049
rect 13133 -18109 13193 -18049
rect 13271 -18109 13331 -18049
rect 13591 -18109 13651 -18049
rect 13727 -18109 13787 -18049
rect 14047 -18109 14107 -18049
rect 14183 -18109 14243 -18049
rect 14503 -18109 14563 -18049
rect 14641 -18109 14701 -18049
rect 14961 -18109 15021 -18049
rect 15097 -18109 15157 -18049
rect 15417 -18109 15477 -18049
rect 12357 -18459 12417 -18399
rect 12677 -18459 12737 -18399
rect 12813 -18459 12873 -18399
rect 13133 -18459 13193 -18399
rect 13271 -18459 13331 -18399
rect 13591 -18459 13651 -18399
rect 13727 -18459 13787 -18399
rect 14047 -18459 14107 -18399
rect 14183 -18459 14243 -18399
rect 14503 -18459 14563 -18399
rect 14641 -18459 14701 -18399
rect 14961 -18459 15021 -18399
rect 15097 -18459 15157 -18399
rect 15417 -18459 15477 -18399
rect 11 -18611 14 -18551
rect 14 -18611 66 -18551
rect 66 -18611 71 -18551
rect 331 -18611 391 -18551
rect 11 -18961 14 -18901
rect 14 -18961 66 -18901
rect 66 -18961 71 -18901
rect 331 -18961 391 -18901
rect 467 -18611 527 -18551
rect 787 -18611 847 -18551
rect 923 -18611 983 -18551
rect 1243 -18611 1303 -18551
rect 1381 -18611 1441 -18551
rect 1701 -18611 1761 -18551
rect 1837 -18611 1897 -18551
rect 2157 -18611 2217 -18551
rect 2293 -18611 2353 -18551
rect 2613 -18611 2673 -18551
rect 2751 -18611 2811 -18551
rect 3071 -18611 3131 -18551
rect 3207 -18611 3267 -18551
rect 3527 -18611 3587 -18551
rect 467 -18961 527 -18901
rect 787 -18961 847 -18901
rect 923 -18961 983 -18901
rect 1243 -18961 1303 -18901
rect 1381 -18961 1441 -18901
rect 1701 -18961 1761 -18901
rect 1837 -18961 1897 -18901
rect 2157 -18961 2217 -18901
rect 2293 -18961 2353 -18901
rect 2613 -18961 2673 -18901
rect 2751 -18961 2811 -18901
rect 3071 -18961 3131 -18901
rect 3207 -18961 3267 -18901
rect 3527 -18961 3587 -18901
rect 3663 -18611 3723 -18551
rect 3983 -18611 4043 -18551
rect 4121 -18611 4181 -18551
rect 4441 -18611 4501 -18551
rect 4577 -18611 4637 -18551
rect 4897 -18611 4957 -18551
rect 5033 -18611 5093 -18551
rect 5353 -18611 5413 -18551
rect 5491 -18611 5551 -18551
rect 5811 -18611 5871 -18551
rect 5947 -18611 6007 -18551
rect 6267 -18611 6327 -18551
rect 6403 -18611 6463 -18551
rect 6723 -18611 6783 -18551
rect 6861 -18611 6921 -18551
rect 7181 -18611 7241 -18551
rect 3663 -18961 3723 -18901
rect 3983 -18961 4043 -18901
rect 4121 -18961 4181 -18901
rect 4441 -18961 4501 -18901
rect 4577 -18961 4637 -18901
rect 4897 -18961 4957 -18901
rect 5033 -18961 5093 -18901
rect 5353 -18961 5413 -18901
rect 5491 -18961 5551 -18901
rect 5811 -18961 5871 -18901
rect 5947 -18961 6007 -18901
rect 6267 -18961 6327 -18901
rect 6403 -18961 6463 -18901
rect 6723 -18961 6783 -18901
rect 6861 -18961 6921 -18901
rect 7181 -18961 7241 -18901
rect 7317 -18611 7377 -18551
rect 7637 -18611 7697 -18551
rect 7773 -18611 7833 -18551
rect 8093 -18611 8153 -18551
rect 8247 -18611 8307 -18551
rect 8567 -18611 8627 -18551
rect 8703 -18611 8763 -18551
rect 9023 -18611 9083 -18551
rect 9161 -18611 9221 -18551
rect 9481 -18611 9541 -18551
rect 9617 -18611 9677 -18551
rect 9937 -18611 9997 -18551
rect 10073 -18611 10133 -18551
rect 10393 -18611 10453 -18551
rect 10531 -18611 10591 -18551
rect 10851 -18611 10911 -18551
rect 7317 -18961 7377 -18901
rect 7637 -18961 7697 -18901
rect 7773 -18961 7833 -18901
rect 8093 -18961 8153 -18901
rect 8247 -18961 8307 -18901
rect 8567 -18961 8627 -18901
rect 8703 -18961 8763 -18901
rect 9023 -18961 9083 -18901
rect 9161 -18961 9221 -18901
rect 9481 -18961 9541 -18901
rect 9617 -18961 9677 -18901
rect 9937 -18961 9997 -18901
rect 10073 -18961 10133 -18901
rect 10393 -18961 10453 -18901
rect 10531 -18961 10591 -18901
rect 10851 -18961 10911 -18901
rect 10987 -18611 11047 -18551
rect 11307 -18611 11367 -18551
rect 11443 -18611 11503 -18551
rect 11763 -18611 11823 -18551
rect 11901 -18611 11961 -18551
rect 12221 -18611 12281 -18551
rect 12357 -18611 12417 -18551
rect 12677 -18611 12737 -18551
rect 12813 -18611 12873 -18551
rect 13133 -18611 13193 -18551
rect 13271 -18611 13331 -18551
rect 13591 -18611 13651 -18551
rect 13727 -18611 13787 -18551
rect 14047 -18611 14107 -18551
rect 14183 -18611 14243 -18551
rect 14503 -18611 14563 -18551
rect 14641 -18611 14701 -18551
rect 14961 -18611 15021 -18551
rect 15097 -18611 15157 -18551
rect 15417 -18611 15477 -18551
rect 10987 -18961 11047 -18901
rect 11307 -18961 11367 -18901
rect 11443 -18961 11503 -18901
rect 11763 -18961 11823 -18901
rect 11901 -18961 11961 -18901
rect 12221 -18961 12281 -18901
rect 12357 -18961 12417 -18901
rect 12677 -18961 12737 -18901
rect 12813 -18961 12873 -18901
rect 13133 -18961 13193 -18901
rect 13271 -18961 13331 -18901
rect 13591 -18961 13651 -18901
rect 13727 -18961 13787 -18901
rect 14047 -18961 14107 -18901
rect 14183 -18961 14243 -18901
rect 14503 -18961 14563 -18901
rect 14641 -18961 14701 -18901
rect 14961 -18961 15021 -18901
rect 15097 -18961 15157 -18901
rect 15417 -18961 15477 -18901
rect 11 -19103 14 -19043
rect 14 -19103 66 -19043
rect 66 -19103 71 -19043
rect 331 -19103 391 -19043
rect 11 -19453 14 -19393
rect 14 -19453 66 -19393
rect 66 -19453 71 -19393
rect 331 -19453 391 -19393
rect 467 -19103 527 -19043
rect 787 -19103 847 -19043
rect 923 -19103 983 -19043
rect 1243 -19103 1303 -19043
rect 1381 -19103 1441 -19043
rect 1701 -19103 1761 -19043
rect 1837 -19103 1897 -19043
rect 2157 -19103 2217 -19043
rect 2293 -19103 2353 -19043
rect 2613 -19103 2673 -19043
rect 2751 -19103 2811 -19043
rect 3071 -19103 3131 -19043
rect 3207 -19103 3267 -19043
rect 3527 -19103 3587 -19043
rect 467 -19453 527 -19393
rect 787 -19453 847 -19393
rect 923 -19453 983 -19393
rect 1243 -19453 1303 -19393
rect 1381 -19453 1441 -19393
rect 1701 -19453 1761 -19393
rect 1837 -19453 1897 -19393
rect 2157 -19453 2217 -19393
rect 2293 -19453 2353 -19393
rect 2613 -19453 2673 -19393
rect 2751 -19453 2811 -19393
rect 3071 -19453 3131 -19393
rect 3207 -19453 3267 -19393
rect 3527 -19453 3587 -19393
rect 3663 -19103 3723 -19043
rect 3983 -19103 4043 -19043
rect 4121 -19103 4181 -19043
rect 4441 -19103 4501 -19043
rect 4577 -19103 4637 -19043
rect 4897 -19103 4957 -19043
rect 5033 -19103 5093 -19043
rect 5353 -19103 5413 -19043
rect 5491 -19103 5551 -19043
rect 5811 -19103 5871 -19043
rect 5947 -19103 6007 -19043
rect 6267 -19103 6327 -19043
rect 6403 -19103 6463 -19043
rect 6723 -19103 6783 -19043
rect 6861 -19103 6921 -19043
rect 7181 -19103 7241 -19043
rect 3663 -19453 3723 -19393
rect 3983 -19453 4043 -19393
rect 4121 -19453 4181 -19393
rect 4441 -19453 4501 -19393
rect 4577 -19453 4637 -19393
rect 4897 -19453 4957 -19393
rect 5033 -19453 5093 -19393
rect 5353 -19453 5413 -19393
rect 5491 -19453 5551 -19393
rect 5811 -19453 5871 -19393
rect 5947 -19453 6007 -19393
rect 6267 -19453 6327 -19393
rect 6403 -19453 6463 -19393
rect 6723 -19453 6783 -19393
rect 6861 -19453 6921 -19393
rect 7181 -19453 7241 -19393
rect 7317 -19103 7377 -19043
rect 7637 -19103 7697 -19043
rect 7773 -19103 7833 -19043
rect 8093 -19103 8153 -19043
rect 8247 -19103 8307 -19043
rect 8567 -19103 8627 -19043
rect 8703 -19103 8763 -19043
rect 9023 -19103 9083 -19043
rect 9161 -19103 9221 -19043
rect 9481 -19103 9541 -19043
rect 9617 -19103 9677 -19043
rect 9937 -19103 9997 -19043
rect 10073 -19103 10133 -19043
rect 10393 -19103 10453 -19043
rect 10531 -19103 10591 -19043
rect 10851 -19103 10911 -19043
rect 7317 -19453 7377 -19393
rect 7637 -19453 7697 -19393
rect 7773 -19453 7833 -19393
rect 8093 -19453 8153 -19393
rect 8247 -19453 8307 -19393
rect 8567 -19453 8627 -19393
rect 8703 -19453 8763 -19393
rect 9023 -19453 9083 -19393
rect 9161 -19453 9221 -19393
rect 9481 -19453 9541 -19393
rect 9617 -19453 9677 -19393
rect 9937 -19453 9997 -19393
rect 10073 -19453 10133 -19393
rect 10393 -19453 10453 -19393
rect 10531 -19453 10591 -19393
rect 10851 -19453 10911 -19393
rect 10987 -19103 11047 -19043
rect 11307 -19103 11367 -19043
rect 11443 -19103 11503 -19043
rect 11763 -19103 11823 -19043
rect 11901 -19103 11961 -19043
rect 12221 -19103 12281 -19043
rect 12357 -19103 12417 -19043
rect 12677 -19103 12737 -19043
rect 12813 -19103 12873 -19043
rect 13133 -19103 13193 -19043
rect 13271 -19103 13331 -19043
rect 13591 -19103 13651 -19043
rect 13727 -19103 13787 -19043
rect 14047 -19103 14107 -19043
rect 14183 -19103 14243 -19043
rect 14503 -19103 14563 -19043
rect 14641 -19103 14701 -19043
rect 14961 -19103 15021 -19043
rect 15097 -19103 15157 -19043
rect 15417 -19103 15477 -19043
rect 10987 -19453 11047 -19393
rect 11307 -19453 11367 -19393
rect 11443 -19453 11503 -19393
rect 11763 -19453 11823 -19393
rect 11901 -19453 11961 -19393
rect 12221 -19453 12281 -19393
rect 12357 -19453 12417 -19393
rect 12677 -19453 12737 -19393
rect 12813 -19453 12873 -19393
rect 13133 -19453 13193 -19393
rect 13271 -19453 13331 -19393
rect 13591 -19453 13651 -19393
rect 13727 -19453 13787 -19393
rect 14047 -19453 14107 -19393
rect 14183 -19453 14243 -19393
rect 14503 -19453 14563 -19393
rect 14641 -19453 14701 -19393
rect 14961 -19453 15021 -19393
rect 15097 -19453 15157 -19393
rect 15417 -19453 15477 -19393
rect 11 -19597 14 -19537
rect 14 -19597 66 -19537
rect 66 -19597 71 -19537
rect 331 -19597 391 -19537
rect 11 -19947 14 -19887
rect 14 -19947 66 -19887
rect 66 -19947 71 -19887
rect 331 -19947 391 -19887
rect 467 -19597 527 -19537
rect 787 -19597 847 -19537
rect 923 -19597 983 -19537
rect 1243 -19597 1303 -19537
rect 1381 -19597 1441 -19537
rect 1701 -19597 1761 -19537
rect 1837 -19597 1897 -19537
rect 2157 -19597 2217 -19537
rect 2293 -19597 2353 -19537
rect 2613 -19597 2673 -19537
rect 2751 -19597 2811 -19537
rect 3071 -19597 3131 -19537
rect 3207 -19597 3267 -19537
rect 3527 -19597 3587 -19537
rect 467 -19947 527 -19887
rect 787 -19947 847 -19887
rect 923 -19947 983 -19887
rect 1243 -19947 1303 -19887
rect 1381 -19947 1441 -19887
rect 1701 -19947 1761 -19887
rect 1837 -19947 1897 -19887
rect 2157 -19947 2217 -19887
rect 2293 -19947 2353 -19887
rect 2613 -19947 2673 -19887
rect 2751 -19947 2811 -19887
rect 3071 -19947 3131 -19887
rect 3207 -19947 3267 -19887
rect 3527 -19947 3587 -19887
rect 3663 -19597 3723 -19537
rect 3983 -19597 4043 -19537
rect 4121 -19597 4181 -19537
rect 4441 -19597 4501 -19537
rect 4577 -19597 4637 -19537
rect 4897 -19597 4957 -19537
rect 5033 -19597 5093 -19537
rect 5353 -19597 5413 -19537
rect 5491 -19597 5551 -19537
rect 5811 -19597 5871 -19537
rect 5947 -19597 6007 -19537
rect 6267 -19597 6327 -19537
rect 6403 -19597 6463 -19537
rect 6723 -19597 6783 -19537
rect 6861 -19597 6921 -19537
rect 7181 -19597 7241 -19537
rect 3663 -19947 3723 -19887
rect 3983 -19947 4043 -19887
rect 4121 -19947 4181 -19887
rect 4441 -19947 4501 -19887
rect 4577 -19947 4637 -19887
rect 4897 -19947 4957 -19887
rect 5033 -19947 5093 -19887
rect 5353 -19947 5413 -19887
rect 5491 -19947 5551 -19887
rect 5811 -19947 5871 -19887
rect 5947 -19947 6007 -19887
rect 6267 -19947 6327 -19887
rect 6403 -19947 6463 -19887
rect 6723 -19947 6783 -19887
rect 6861 -19947 6921 -19887
rect 7181 -19947 7241 -19887
rect 7317 -19597 7377 -19537
rect 7637 -19597 7697 -19537
rect 7773 -19597 7833 -19537
rect 8093 -19597 8153 -19537
rect 8247 -19597 8307 -19537
rect 8567 -19597 8627 -19537
rect 8703 -19597 8763 -19537
rect 9023 -19597 9083 -19537
rect 9161 -19597 9221 -19537
rect 9481 -19597 9541 -19537
rect 9617 -19597 9677 -19537
rect 9937 -19597 9997 -19537
rect 10073 -19597 10133 -19537
rect 10393 -19597 10453 -19537
rect 10531 -19597 10591 -19537
rect 10851 -19597 10911 -19537
rect 10987 -19597 11047 -19537
rect 11307 -19597 11367 -19537
rect 11443 -19597 11503 -19537
rect 11763 -19597 11823 -19537
rect 11901 -19597 11961 -19537
rect 12221 -19597 12281 -19537
rect 12357 -19597 12417 -19537
rect 12677 -19597 12737 -19537
rect 12813 -19597 12873 -19537
rect 13133 -19597 13193 -19537
rect 13271 -19597 13331 -19537
rect 13591 -19597 13651 -19537
rect 13727 -19597 13787 -19537
rect 14047 -19597 14107 -19537
rect 14183 -19597 14243 -19537
rect 14503 -19597 14563 -19537
rect 14641 -19597 14701 -19537
rect 14961 -19597 15021 -19537
rect 15097 -19597 15157 -19537
rect 15417 -19597 15477 -19537
rect 7317 -19947 7377 -19887
rect 7637 -19947 7697 -19887
rect 7773 -19947 7833 -19887
rect 8093 -19947 8153 -19887
rect 8247 -19947 8307 -19887
rect 8567 -19947 8627 -19887
rect 8703 -19947 8763 -19887
rect 9023 -19947 9083 -19887
rect 9161 -19947 9221 -19887
rect 9481 -19947 9541 -19887
rect 9617 -19947 9677 -19887
rect 9937 -19947 9997 -19887
rect 10073 -19947 10133 -19887
rect 10393 -19947 10453 -19887
rect 10531 -19947 10591 -19887
rect 10851 -19947 10911 -19887
rect 10987 -19947 11047 -19887
rect 11307 -19947 11367 -19887
rect 11443 -19947 11503 -19887
rect 11763 -19947 11823 -19887
rect 11901 -19947 11961 -19887
rect 12221 -19947 12281 -19887
rect 12357 -19947 12417 -19887
rect 12677 -19947 12737 -19887
rect 12813 -19947 12873 -19887
rect 13133 -19947 13193 -19887
rect 13271 -19947 13331 -19887
rect 13591 -19947 13651 -19887
rect 13727 -19947 13787 -19887
rect 14047 -19947 14107 -19887
rect 14183 -19947 14243 -19887
rect 14503 -19947 14563 -19887
rect 14641 -19947 14701 -19887
rect 14961 -19947 15021 -19887
rect 15097 -19947 15157 -19887
rect 15417 -19947 15477 -19887
rect 11 -20099 14 -20039
rect 14 -20099 66 -20039
rect 66 -20099 71 -20039
rect 331 -20099 391 -20039
rect 11 -20449 14 -20389
rect 14 -20449 66 -20389
rect 66 -20449 71 -20389
rect 331 -20449 391 -20389
rect 467 -20099 527 -20039
rect 787 -20099 847 -20039
rect 923 -20099 983 -20039
rect 1243 -20099 1303 -20039
rect 1381 -20099 1441 -20039
rect 1701 -20099 1761 -20039
rect 1837 -20099 1897 -20039
rect 2157 -20099 2217 -20039
rect 2293 -20099 2353 -20039
rect 2613 -20099 2673 -20039
rect 2751 -20099 2811 -20039
rect 3071 -20099 3131 -20039
rect 3207 -20099 3267 -20039
rect 3527 -20099 3587 -20039
rect 3663 -20099 3723 -20039
rect 3983 -20099 4043 -20039
rect 467 -20449 527 -20389
rect 787 -20449 847 -20389
rect 923 -20449 983 -20389
rect 1243 -20449 1303 -20389
rect 1381 -20449 1441 -20389
rect 1701 -20449 1761 -20389
rect 1837 -20449 1897 -20389
rect 2157 -20449 2217 -20389
rect 2293 -20449 2353 -20389
rect 2613 -20449 2673 -20389
rect 2751 -20449 2811 -20389
rect 3071 -20449 3131 -20389
rect 3207 -20449 3267 -20389
rect 3527 -20449 3587 -20389
rect 3663 -20449 3723 -20389
rect 3983 -20449 4043 -20389
rect 4121 -20099 4181 -20039
rect 4441 -20099 4501 -20039
rect 4577 -20099 4637 -20039
rect 4897 -20099 4957 -20039
rect 5033 -20099 5093 -20039
rect 5353 -20099 5413 -20039
rect 5491 -20099 5551 -20039
rect 5811 -20099 5871 -20039
rect 5947 -20099 6007 -20039
rect 6267 -20099 6327 -20039
rect 6403 -20099 6463 -20039
rect 6723 -20099 6783 -20039
rect 6861 -20099 6921 -20039
rect 7181 -20099 7241 -20039
rect 4121 -20449 4181 -20389
rect 4441 -20449 4501 -20389
rect 4577 -20449 4637 -20389
rect 4897 -20449 4957 -20389
rect 5033 -20449 5093 -20389
rect 5353 -20449 5413 -20389
rect 5491 -20449 5551 -20389
rect 5811 -20449 5871 -20389
rect 5947 -20449 6007 -20389
rect 6267 -20449 6327 -20389
rect 6403 -20449 6463 -20389
rect 6723 -20449 6783 -20389
rect 6861 -20449 6921 -20389
rect 7181 -20449 7241 -20389
rect 7317 -20099 7377 -20039
rect 7637 -20099 7697 -20039
rect 7773 -20099 7833 -20039
rect 8093 -20099 8153 -20039
rect 8247 -20099 8307 -20039
rect 8567 -20099 8627 -20039
rect 8703 -20099 8763 -20039
rect 9023 -20099 9083 -20039
rect 9161 -20099 9221 -20039
rect 9481 -20099 9541 -20039
rect 7317 -20449 7377 -20389
rect 7637 -20449 7697 -20389
rect 7773 -20449 7833 -20389
rect 8093 -20449 8153 -20389
rect 8247 -20449 8307 -20389
rect 8567 -20449 8627 -20389
rect 8703 -20449 8763 -20389
rect 9023 -20449 9083 -20389
rect 9161 -20449 9221 -20389
rect 9481 -20449 9541 -20389
rect 9617 -20099 9677 -20039
rect 9937 -20099 9997 -20039
rect 10073 -20099 10133 -20039
rect 10393 -20099 10453 -20039
rect 10531 -20099 10591 -20039
rect 10851 -20099 10911 -20039
rect 10987 -20099 11047 -20039
rect 11307 -20099 11367 -20039
rect 11443 -20099 11503 -20039
rect 11763 -20099 11823 -20039
rect 11901 -20099 11961 -20039
rect 12221 -20099 12281 -20039
rect 12357 -20099 12417 -20039
rect 12677 -20099 12737 -20039
rect 12813 -20099 12873 -20039
rect 13133 -20099 13193 -20039
rect 13271 -20099 13331 -20039
rect 13591 -20099 13651 -20039
rect 13727 -20099 13787 -20039
rect 14047 -20099 14107 -20039
rect 14183 -20099 14243 -20039
rect 14503 -20099 14563 -20039
rect 14641 -20099 14701 -20039
rect 14961 -20099 15021 -20039
rect 15097 -20099 15157 -20039
rect 15417 -20099 15477 -20039
rect 9617 -20449 9677 -20389
rect 9937 -20449 9997 -20389
rect 10073 -20449 10133 -20389
rect 10393 -20449 10453 -20389
rect 10531 -20449 10591 -20389
rect 10851 -20449 10911 -20389
rect 10987 -20449 11047 -20389
rect 11307 -20449 11367 -20389
rect 11443 -20449 11503 -20389
rect 11763 -20449 11823 -20389
rect 11901 -20449 11961 -20389
rect 12221 -20449 12281 -20389
rect 12357 -20449 12417 -20389
rect 12677 -20449 12737 -20389
rect 12813 -20449 12873 -20389
rect 13133 -20449 13193 -20389
rect 13271 -20449 13331 -20389
rect 13591 -20449 13651 -20389
rect 13727 -20449 13787 -20389
rect 14047 -20449 14107 -20389
rect 14183 -20449 14243 -20389
rect 14503 -20449 14563 -20389
rect 14641 -20449 14701 -20389
rect 14961 -20449 15021 -20389
rect 15097 -20449 15157 -20389
rect 15417 -20449 15477 -20389
rect 11 -20591 14 -20531
rect 14 -20591 66 -20531
rect 66 -20591 71 -20531
rect 331 -20591 391 -20531
rect 11 -20941 14 -20881
rect 14 -20941 66 -20881
rect 66 -20941 71 -20881
rect 331 -20941 391 -20881
rect 467 -20591 527 -20531
rect 787 -20591 847 -20531
rect 923 -20591 983 -20531
rect 1243 -20591 1303 -20531
rect 1381 -20591 1441 -20531
rect 1701 -20591 1761 -20531
rect 1837 -20591 1897 -20531
rect 2157 -20591 2217 -20531
rect 2293 -20591 2353 -20531
rect 2613 -20591 2673 -20531
rect 2751 -20591 2811 -20531
rect 3071 -20591 3131 -20531
rect 3207 -20591 3267 -20531
rect 3527 -20591 3587 -20531
rect 3663 -20591 3723 -20531
rect 3983 -20591 4043 -20531
rect 467 -20941 527 -20881
rect 787 -20941 847 -20881
rect 923 -20941 983 -20881
rect 1243 -20941 1303 -20881
rect 1381 -20941 1441 -20881
rect 1701 -20941 1761 -20881
rect 1837 -20941 1897 -20881
rect 2157 -20941 2217 -20881
rect 2293 -20941 2353 -20881
rect 2613 -20941 2673 -20881
rect 2751 -20941 2811 -20881
rect 3071 -20941 3131 -20881
rect 3207 -20941 3267 -20881
rect 3527 -20941 3587 -20881
rect 3663 -20941 3723 -20881
rect 3983 -20941 4043 -20881
rect 4121 -20591 4181 -20531
rect 4441 -20591 4501 -20531
rect 4577 -20591 4637 -20531
rect 4897 -20591 4957 -20531
rect 5033 -20591 5093 -20531
rect 5353 -20591 5413 -20531
rect 5491 -20591 5551 -20531
rect 5811 -20591 5871 -20531
rect 5947 -20591 6007 -20531
rect 6267 -20591 6327 -20531
rect 6403 -20591 6463 -20531
rect 6723 -20591 6783 -20531
rect 6861 -20591 6921 -20531
rect 7181 -20591 7241 -20531
rect 4121 -20941 4181 -20881
rect 4441 -20941 4501 -20881
rect 4577 -20941 4637 -20881
rect 4897 -20941 4957 -20881
rect 5033 -20941 5093 -20881
rect 5353 -20941 5413 -20881
rect 5491 -20941 5551 -20881
rect 5811 -20941 5871 -20881
rect 5947 -20941 6007 -20881
rect 6267 -20941 6327 -20881
rect 6403 -20941 6463 -20881
rect 6723 -20941 6783 -20881
rect 6861 -20941 6921 -20881
rect 7181 -20941 7241 -20881
rect 7317 -20591 7377 -20531
rect 7637 -20591 7697 -20531
rect 7773 -20591 7833 -20531
rect 8093 -20591 8153 -20531
rect 8247 -20591 8307 -20531
rect 8567 -20591 8627 -20531
rect 8703 -20591 8763 -20531
rect 9023 -20591 9083 -20531
rect 9161 -20591 9221 -20531
rect 9481 -20591 9541 -20531
rect 7317 -20941 7377 -20881
rect 7637 -20941 7697 -20881
rect 7773 -20941 7833 -20881
rect 8093 -20941 8153 -20881
rect 8247 -20941 8307 -20881
rect 8567 -20941 8627 -20881
rect 8703 -20941 8763 -20881
rect 9023 -20941 9083 -20881
rect 9161 -20941 9221 -20881
rect 9481 -20941 9541 -20881
rect 9617 -20591 9677 -20531
rect 9937 -20591 9997 -20531
rect 10073 -20591 10133 -20531
rect 10393 -20591 10453 -20531
rect 10531 -20591 10591 -20531
rect 10851 -20591 10911 -20531
rect 10987 -20591 11047 -20531
rect 11307 -20591 11367 -20531
rect 11443 -20591 11503 -20531
rect 11763 -20591 11823 -20531
rect 11901 -20591 11961 -20531
rect 12221 -20591 12281 -20531
rect 12357 -20591 12417 -20531
rect 12677 -20591 12737 -20531
rect 12813 -20591 12873 -20531
rect 13133 -20591 13193 -20531
rect 13271 -20591 13331 -20531
rect 13591 -20591 13651 -20531
rect 13727 -20591 13787 -20531
rect 14047 -20591 14107 -20531
rect 14183 -20591 14243 -20531
rect 14503 -20591 14563 -20531
rect 14641 -20591 14701 -20531
rect 14961 -20591 15021 -20531
rect 15097 -20591 15157 -20531
rect 15417 -20591 15477 -20531
rect 9617 -20941 9677 -20881
rect 9937 -20941 9997 -20881
rect 10073 -20941 10133 -20881
rect 10393 -20941 10453 -20881
rect 10531 -20941 10591 -20881
rect 10851 -20941 10911 -20881
rect 10987 -20941 11047 -20881
rect 11307 -20941 11367 -20881
rect 11443 -20941 11503 -20881
rect 11763 -20941 11823 -20881
rect 11901 -20941 11961 -20881
rect 12221 -20941 12281 -20881
rect 12357 -20941 12417 -20881
rect 12677 -20941 12737 -20881
rect 12813 -20941 12873 -20881
rect 13133 -20941 13193 -20881
rect 13271 -20941 13331 -20881
rect 13591 -20941 13651 -20881
rect 13727 -20941 13787 -20881
rect 14047 -20941 14107 -20881
rect 14183 -20941 14243 -20881
rect 14503 -20941 14563 -20881
rect 14641 -20941 14701 -20881
rect 14961 -20941 15021 -20881
rect 15097 -20941 15157 -20881
rect 15417 -20941 15477 -20881
rect 11 -21107 14 -21047
rect 14 -21107 66 -21047
rect 66 -21107 71 -21047
rect 331 -21107 391 -21047
rect 11 -21457 14 -21397
rect 14 -21457 66 -21397
rect 66 -21457 71 -21397
rect 331 -21457 391 -21397
rect 467 -21107 527 -21047
rect 787 -21107 847 -21047
rect 923 -21107 983 -21047
rect 1243 -21107 1303 -21047
rect 1381 -21107 1441 -21047
rect 1701 -21107 1761 -21047
rect 1837 -21107 1897 -21047
rect 2157 -21107 2217 -21047
rect 2293 -21107 2353 -21047
rect 2613 -21107 2673 -21047
rect 2751 -21107 2811 -21047
rect 3071 -21107 3131 -21047
rect 3207 -21107 3267 -21047
rect 3527 -21107 3587 -21047
rect 3663 -21107 3723 -21047
rect 3983 -21107 4043 -21047
rect 467 -21457 527 -21397
rect 787 -21457 847 -21397
rect 923 -21457 983 -21397
rect 1243 -21457 1303 -21397
rect 1381 -21457 1441 -21397
rect 1701 -21457 1761 -21397
rect 1837 -21457 1897 -21397
rect 2157 -21457 2217 -21397
rect 2293 -21457 2353 -21397
rect 2613 -21457 2673 -21397
rect 2751 -21457 2811 -21397
rect 3071 -21457 3131 -21397
rect 3207 -21457 3267 -21397
rect 3527 -21457 3587 -21397
rect 3663 -21457 3723 -21397
rect 3983 -21457 4043 -21397
rect 4121 -21107 4181 -21047
rect 4441 -21107 4501 -21047
rect 4577 -21107 4637 -21047
rect 4897 -21107 4957 -21047
rect 5033 -21107 5093 -21047
rect 5353 -21107 5413 -21047
rect 5491 -21107 5551 -21047
rect 5811 -21107 5871 -21047
rect 5947 -21107 6007 -21047
rect 6267 -21107 6327 -21047
rect 6403 -21107 6463 -21047
rect 6723 -21107 6783 -21047
rect 6861 -21107 6921 -21047
rect 7181 -21107 7241 -21047
rect 4121 -21457 4181 -21397
rect 4441 -21457 4501 -21397
rect 4577 -21457 4637 -21397
rect 4897 -21457 4957 -21397
rect 5033 -21457 5093 -21397
rect 5353 -21457 5413 -21397
rect 5491 -21457 5551 -21397
rect 5811 -21457 5871 -21397
rect 5947 -21457 6007 -21397
rect 6267 -21457 6327 -21397
rect 6403 -21457 6463 -21397
rect 6723 -21457 6783 -21397
rect 6861 -21457 6921 -21397
rect 7181 -21457 7241 -21397
rect 7317 -21107 7377 -21047
rect 7637 -21107 7697 -21047
rect 7773 -21107 7833 -21047
rect 8093 -21107 8153 -21047
rect 8247 -21107 8307 -21047
rect 8567 -21107 8627 -21047
rect 8703 -21107 8763 -21047
rect 9023 -21107 9083 -21047
rect 9161 -21107 9221 -21047
rect 9481 -21107 9541 -21047
rect 9617 -21107 9677 -21047
rect 9937 -21107 9997 -21047
rect 10073 -21107 10133 -21047
rect 10393 -21107 10453 -21047
rect 10531 -21107 10591 -21047
rect 10851 -21107 10911 -21047
rect 10987 -21107 11047 -21047
rect 11307 -21107 11367 -21047
rect 11443 -21107 11503 -21047
rect 11763 -21107 11823 -21047
rect 11901 -21107 11961 -21047
rect 12221 -21107 12281 -21047
rect 12357 -21107 12417 -21047
rect 12677 -21107 12737 -21047
rect 12813 -21107 12873 -21047
rect 13133 -21107 13193 -21047
rect 13271 -21107 13331 -21047
rect 13591 -21107 13651 -21047
rect 13727 -21107 13787 -21047
rect 14047 -21107 14107 -21047
rect 14183 -21107 14243 -21047
rect 14503 -21107 14563 -21047
rect 14641 -21107 14701 -21047
rect 14961 -21107 15021 -21047
rect 15097 -21107 15157 -21047
rect 15417 -21107 15477 -21047
rect 7317 -21457 7377 -21397
rect 7637 -21457 7697 -21397
rect 7773 -21457 7833 -21397
rect 8093 -21457 8153 -21397
rect 8247 -21457 8307 -21397
rect 8567 -21457 8627 -21397
rect 8703 -21457 8763 -21397
rect 9023 -21457 9083 -21397
rect 9161 -21457 9221 -21397
rect 9481 -21457 9541 -21397
rect 9617 -21457 9677 -21397
rect 9937 -21457 9997 -21397
rect 10073 -21457 10133 -21397
rect 10393 -21457 10453 -21397
rect 10531 -21457 10591 -21397
rect 10851 -21457 10911 -21397
rect 10987 -21457 11047 -21397
rect 11307 -21457 11367 -21397
rect 11443 -21457 11503 -21397
rect 11763 -21457 11823 -21397
rect 11901 -21457 11961 -21397
rect 12221 -21457 12281 -21397
rect 12357 -21457 12417 -21397
rect 12677 -21457 12737 -21397
rect 12813 -21457 12873 -21397
rect 13133 -21457 13193 -21397
rect 13271 -21457 13331 -21397
rect 13591 -21457 13651 -21397
rect 13727 -21457 13787 -21397
rect 14047 -21457 14107 -21397
rect 14183 -21457 14243 -21397
rect 14503 -21457 14563 -21397
rect 14641 -21457 14701 -21397
rect 14961 -21457 15021 -21397
rect 15097 -21457 15157 -21397
rect 15417 -21457 15477 -21397
rect 11 -21609 14 -21549
rect 14 -21609 66 -21549
rect 66 -21609 71 -21549
rect 331 -21609 391 -21549
rect 11 -21959 14 -21899
rect 14 -21959 66 -21899
rect 66 -21959 71 -21899
rect 331 -21959 391 -21899
rect 467 -21609 527 -21549
rect 787 -21609 847 -21549
rect 923 -21609 983 -21549
rect 1243 -21609 1303 -21549
rect 1381 -21609 1441 -21549
rect 1701 -21609 1761 -21549
rect 1837 -21609 1897 -21549
rect 2157 -21609 2217 -21549
rect 2293 -21609 2353 -21549
rect 2613 -21609 2673 -21549
rect 2751 -21609 2811 -21549
rect 3071 -21609 3131 -21549
rect 3207 -21609 3267 -21549
rect 3527 -21609 3587 -21549
rect 3663 -21609 3723 -21549
rect 3983 -21609 4043 -21549
rect 467 -21959 527 -21899
rect 787 -21959 847 -21899
rect 923 -21959 983 -21899
rect 1243 -21959 1303 -21899
rect 1381 -21959 1441 -21899
rect 1701 -21959 1761 -21899
rect 1837 -21959 1897 -21899
rect 2157 -21959 2217 -21899
rect 2293 -21959 2353 -21899
rect 2613 -21959 2673 -21899
rect 2751 -21959 2811 -21899
rect 3071 -21959 3131 -21899
rect 3207 -21959 3267 -21899
rect 3527 -21959 3587 -21899
rect 3663 -21959 3723 -21899
rect 3983 -21959 4043 -21899
rect 4121 -21609 4181 -21549
rect 4441 -21609 4501 -21549
rect 4577 -21609 4637 -21549
rect 4897 -21609 4957 -21549
rect 5033 -21609 5093 -21549
rect 5353 -21609 5413 -21549
rect 5491 -21609 5551 -21549
rect 5811 -21609 5871 -21549
rect 5947 -21609 6007 -21549
rect 6267 -21609 6327 -21549
rect 6403 -21609 6463 -21549
rect 6723 -21609 6783 -21549
rect 6861 -21609 6921 -21549
rect 7181 -21609 7241 -21549
rect 4121 -21959 4181 -21899
rect 4441 -21959 4501 -21899
rect 4577 -21959 4637 -21899
rect 4897 -21959 4957 -21899
rect 5033 -21959 5093 -21899
rect 5353 -21959 5413 -21899
rect 5491 -21959 5551 -21899
rect 5811 -21959 5871 -21899
rect 5947 -21959 6007 -21899
rect 6267 -21959 6327 -21899
rect 6403 -21959 6463 -21899
rect 6723 -21959 6783 -21899
rect 6861 -21959 6921 -21899
rect 7181 -21959 7241 -21899
rect 7317 -21609 7377 -21549
rect 7637 -21609 7697 -21549
rect 7773 -21609 7833 -21549
rect 8093 -21609 8153 -21549
rect 8247 -21609 8307 -21549
rect 8567 -21609 8627 -21549
rect 8703 -21609 8763 -21549
rect 9023 -21609 9083 -21549
rect 9161 -21609 9221 -21549
rect 9481 -21609 9541 -21549
rect 9617 -21609 9677 -21549
rect 9937 -21609 9997 -21549
rect 10073 -21609 10133 -21549
rect 10393 -21609 10453 -21549
rect 10531 -21609 10591 -21549
rect 10851 -21609 10911 -21549
rect 10987 -21609 11047 -21549
rect 11307 -21609 11367 -21549
rect 11443 -21609 11503 -21549
rect 11763 -21609 11823 -21549
rect 11901 -21609 11961 -21549
rect 12221 -21609 12281 -21549
rect 12357 -21609 12417 -21549
rect 12677 -21609 12737 -21549
rect 12813 -21609 12873 -21549
rect 13133 -21609 13193 -21549
rect 13271 -21609 13331 -21549
rect 13591 -21609 13651 -21549
rect 13727 -21609 13787 -21549
rect 14047 -21609 14107 -21549
rect 14183 -21609 14243 -21549
rect 14503 -21609 14563 -21549
rect 14641 -21609 14701 -21549
rect 14961 -21609 15021 -21549
rect 15097 -21609 15157 -21549
rect 15417 -21609 15477 -21549
rect 7317 -21959 7377 -21899
rect 7637 -21959 7697 -21899
rect 7773 -21959 7833 -21899
rect 8093 -21959 8153 -21899
rect 8247 -21959 8307 -21899
rect 8567 -21959 8627 -21899
rect 8703 -21959 8763 -21899
rect 9023 -21959 9083 -21899
rect 9161 -21959 9221 -21899
rect 9481 -21959 9541 -21899
rect 9617 -21959 9677 -21899
rect 9937 -21959 9997 -21899
rect 10073 -21959 10133 -21899
rect 10393 -21959 10453 -21899
rect 10531 -21959 10591 -21899
rect 10851 -21959 10911 -21899
rect 10987 -21959 11047 -21899
rect 11307 -21959 11367 -21899
rect 11443 -21959 11503 -21899
rect 11763 -21959 11823 -21899
rect 11901 -21959 11961 -21899
rect 12221 -21959 12281 -21899
rect 12357 -21959 12417 -21899
rect 12677 -21959 12737 -21899
rect 12813 -21959 12873 -21899
rect 13133 -21959 13193 -21899
rect 13271 -21959 13331 -21899
rect 13591 -21959 13651 -21899
rect 13727 -21959 13787 -21899
rect 14047 -21959 14107 -21899
rect 14183 -21959 14243 -21899
rect 14503 -21959 14563 -21899
rect 14641 -21959 14701 -21899
rect 14961 -21959 15021 -21899
rect 15097 -21959 15157 -21899
rect 15417 -21959 15477 -21899
rect 11 -22101 14 -22041
rect 14 -22101 66 -22041
rect 66 -22101 71 -22041
rect 331 -22101 391 -22041
rect 11 -22451 14 -22391
rect 14 -22451 66 -22391
rect 66 -22451 71 -22391
rect 331 -22451 391 -22391
rect 467 -22101 527 -22041
rect 787 -22101 847 -22041
rect 923 -22101 983 -22041
rect 1243 -22101 1303 -22041
rect 1381 -22101 1441 -22041
rect 1701 -22101 1761 -22041
rect 1837 -22101 1897 -22041
rect 2157 -22101 2217 -22041
rect 2293 -22101 2353 -22041
rect 2613 -22101 2673 -22041
rect 2751 -22101 2811 -22041
rect 3071 -22101 3131 -22041
rect 3207 -22101 3267 -22041
rect 3527 -22101 3587 -22041
rect 3663 -22101 3723 -22041
rect 3983 -22101 4043 -22041
rect 467 -22451 527 -22391
rect 787 -22451 847 -22391
rect 923 -22451 983 -22391
rect 1243 -22451 1303 -22391
rect 1381 -22451 1441 -22391
rect 1701 -22451 1761 -22391
rect 1837 -22451 1897 -22391
rect 2157 -22451 2217 -22391
rect 2293 -22451 2353 -22391
rect 2613 -22451 2673 -22391
rect 2751 -22451 2811 -22391
rect 3071 -22451 3131 -22391
rect 3207 -22451 3267 -22391
rect 3527 -22451 3587 -22391
rect 3663 -22451 3723 -22391
rect 3983 -22451 4043 -22391
rect 4121 -22101 4181 -22041
rect 4441 -22101 4501 -22041
rect 4577 -22101 4637 -22041
rect 4897 -22101 4957 -22041
rect 5033 -22101 5093 -22041
rect 5353 -22101 5413 -22041
rect 5491 -22101 5551 -22041
rect 5811 -22101 5871 -22041
rect 5947 -22101 6007 -22041
rect 6267 -22101 6327 -22041
rect 6403 -22101 6463 -22041
rect 6723 -22101 6783 -22041
rect 6861 -22101 6921 -22041
rect 7181 -22101 7241 -22041
rect 4121 -22451 4181 -22391
rect 4441 -22451 4501 -22391
rect 4577 -22451 4637 -22391
rect 4897 -22451 4957 -22391
rect 5033 -22451 5093 -22391
rect 5353 -22451 5413 -22391
rect 5491 -22451 5551 -22391
rect 5811 -22451 5871 -22391
rect 5947 -22451 6007 -22391
rect 6267 -22451 6327 -22391
rect 6403 -22451 6463 -22391
rect 6723 -22451 6783 -22391
rect 6861 -22451 6921 -22391
rect 7181 -22451 7241 -22391
rect 7317 -22101 7377 -22041
rect 7637 -22101 7697 -22041
rect 7773 -22101 7833 -22041
rect 8093 -22101 8153 -22041
rect 8247 -22101 8307 -22041
rect 8567 -22101 8627 -22041
rect 8703 -22101 8763 -22041
rect 9023 -22101 9083 -22041
rect 9161 -22101 9221 -22041
rect 9481 -22101 9541 -22041
rect 9617 -22101 9677 -22041
rect 9937 -22101 9997 -22041
rect 10073 -22101 10133 -22041
rect 10393 -22101 10453 -22041
rect 10531 -22101 10591 -22041
rect 10851 -22101 10911 -22041
rect 10987 -22101 11047 -22041
rect 11307 -22101 11367 -22041
rect 11443 -22101 11503 -22041
rect 11763 -22101 11823 -22041
rect 11901 -22101 11961 -22041
rect 12221 -22101 12281 -22041
rect 12357 -22101 12417 -22041
rect 12677 -22101 12737 -22041
rect 12813 -22101 12873 -22041
rect 13133 -22101 13193 -22041
rect 13271 -22101 13331 -22041
rect 13591 -22101 13651 -22041
rect 13727 -22101 13787 -22041
rect 14047 -22101 14107 -22041
rect 14183 -22101 14243 -22041
rect 14503 -22101 14563 -22041
rect 14641 -22101 14701 -22041
rect 14961 -22101 15021 -22041
rect 15097 -22101 15157 -22041
rect 15417 -22101 15477 -22041
rect 7317 -22451 7377 -22391
rect 7637 -22451 7697 -22391
rect 7773 -22451 7833 -22391
rect 8093 -22451 8153 -22391
rect 8247 -22451 8307 -22391
rect 8567 -22451 8627 -22391
rect 8703 -22451 8763 -22391
rect 9023 -22451 9083 -22391
rect 9161 -22451 9221 -22391
rect 9481 -22451 9541 -22391
rect 9617 -22451 9677 -22391
rect 9937 -22451 9997 -22391
rect 10073 -22451 10133 -22391
rect 10393 -22451 10453 -22391
rect 10531 -22451 10591 -22391
rect 10851 -22451 10911 -22391
rect 10987 -22451 11047 -22391
rect 11307 -22451 11367 -22391
rect 11443 -22451 11503 -22391
rect 11763 -22451 11823 -22391
rect 11901 -22451 11961 -22391
rect 12221 -22451 12281 -22391
rect 12357 -22451 12417 -22391
rect 12677 -22451 12737 -22391
rect 12813 -22451 12873 -22391
rect 13133 -22451 13193 -22391
rect 13271 -22451 13331 -22391
rect 13591 -22451 13651 -22391
rect 13727 -22451 13787 -22391
rect 14047 -22451 14107 -22391
rect 14183 -22451 14243 -22391
rect 14503 -22451 14563 -22391
rect 14641 -22451 14701 -22391
rect 14961 -22451 15021 -22391
rect 15097 -22451 15157 -22391
rect 15417 -22451 15477 -22391
rect 11 -22588 14 -22528
rect 14 -22588 66 -22528
rect 66 -22588 71 -22528
rect 331 -22588 391 -22528
rect 11 -22938 14 -22878
rect 14 -22938 66 -22878
rect 66 -22938 71 -22878
rect 331 -22938 391 -22878
rect 467 -22588 527 -22528
rect 787 -22588 847 -22528
rect 923 -22588 983 -22528
rect 1243 -22588 1303 -22528
rect 1381 -22588 1441 -22528
rect 1701 -22588 1761 -22528
rect 1837 -22588 1897 -22528
rect 2157 -22588 2217 -22528
rect 2293 -22588 2353 -22528
rect 2613 -22588 2673 -22528
rect 2751 -22588 2811 -22528
rect 3071 -22588 3131 -22528
rect 3207 -22588 3267 -22528
rect 3527 -22588 3587 -22528
rect 3663 -22588 3723 -22528
rect 3983 -22588 4043 -22528
rect 467 -22938 527 -22878
rect 787 -22938 847 -22878
rect 923 -22938 983 -22878
rect 1243 -22938 1303 -22878
rect 1381 -22938 1441 -22878
rect 1701 -22938 1761 -22878
rect 1837 -22938 1897 -22878
rect 2157 -22938 2217 -22878
rect 2293 -22938 2353 -22878
rect 2613 -22938 2673 -22878
rect 2751 -22938 2811 -22878
rect 3071 -22938 3131 -22878
rect 3207 -22938 3267 -22878
rect 3527 -22938 3587 -22878
rect 3663 -22938 3723 -22878
rect 3983 -22938 4043 -22878
rect 4121 -22588 4181 -22528
rect 4441 -22588 4501 -22528
rect 4577 -22588 4637 -22528
rect 4897 -22588 4957 -22528
rect 5033 -22588 5093 -22528
rect 5353 -22588 5413 -22528
rect 5491 -22588 5551 -22528
rect 5811 -22588 5871 -22528
rect 5947 -22588 6007 -22528
rect 6267 -22588 6327 -22528
rect 6403 -22588 6463 -22528
rect 6723 -22588 6783 -22528
rect 6861 -22588 6921 -22528
rect 7181 -22588 7241 -22528
rect 4121 -22938 4181 -22878
rect 4441 -22938 4501 -22878
rect 4577 -22938 4637 -22878
rect 4897 -22938 4957 -22878
rect 5033 -22938 5093 -22878
rect 5353 -22938 5413 -22878
rect 5491 -22938 5551 -22878
rect 5811 -22938 5871 -22878
rect 5947 -22938 6007 -22878
rect 6267 -22938 6327 -22878
rect 6403 -22938 6463 -22878
rect 6723 -22938 6783 -22878
rect 6861 -22938 6921 -22878
rect 7181 -22938 7241 -22878
rect 7317 -22588 7377 -22528
rect 7637 -22588 7697 -22528
rect 7773 -22588 7833 -22528
rect 8093 -22588 8153 -22528
rect 8247 -22588 8307 -22528
rect 8567 -22588 8627 -22528
rect 8703 -22588 8763 -22528
rect 9023 -22588 9083 -22528
rect 9161 -22588 9221 -22528
rect 9481 -22588 9541 -22528
rect 9617 -22588 9677 -22528
rect 9937 -22588 9997 -22528
rect 10073 -22588 10133 -22528
rect 10393 -22588 10453 -22528
rect 10531 -22588 10591 -22528
rect 10851 -22588 10911 -22528
rect 10987 -22588 11047 -22528
rect 11307 -22588 11367 -22528
rect 11443 -22588 11503 -22528
rect 11763 -22588 11823 -22528
rect 11901 -22588 11961 -22528
rect 12221 -22588 12281 -22528
rect 12357 -22588 12417 -22528
rect 12677 -22588 12737 -22528
rect 12813 -22588 12873 -22528
rect 13133 -22588 13193 -22528
rect 13271 -22588 13331 -22528
rect 13591 -22588 13651 -22528
rect 13727 -22588 13787 -22528
rect 14047 -22588 14107 -22528
rect 14183 -22588 14243 -22528
rect 14503 -22588 14563 -22528
rect 14641 -22588 14701 -22528
rect 14961 -22588 15021 -22528
rect 15097 -22588 15157 -22528
rect 15417 -22588 15477 -22528
rect 7317 -22938 7377 -22878
rect 7637 -22938 7697 -22878
rect 7773 -22938 7833 -22878
rect 8093 -22938 8153 -22878
rect 8247 -22938 8307 -22878
rect 8567 -22938 8627 -22878
rect 8703 -22938 8763 -22878
rect 9023 -22938 9083 -22878
rect 9161 -22938 9221 -22878
rect 9481 -22938 9541 -22878
rect 9617 -22938 9677 -22878
rect 9937 -22938 9997 -22878
rect 10073 -22938 10133 -22878
rect 10393 -22938 10453 -22878
rect 10531 -22938 10591 -22878
rect 10851 -22938 10911 -22878
rect 10987 -22938 11047 -22878
rect 11307 -22938 11367 -22878
rect 11443 -22938 11503 -22878
rect 11763 -22938 11823 -22878
rect 11901 -22938 11961 -22878
rect 12221 -22938 12281 -22878
rect 12357 -22938 12417 -22878
rect 12677 -22938 12737 -22878
rect 12813 -22938 12873 -22878
rect 13133 -22938 13193 -22878
rect 13271 -22938 13331 -22878
rect 13591 -22938 13651 -22878
rect 13727 -22938 13787 -22878
rect 14047 -22938 14107 -22878
rect 14183 -22938 14243 -22878
rect 14503 -22938 14563 -22878
rect 14641 -22938 14701 -22878
rect 14961 -22938 15021 -22878
rect 15097 -22938 15157 -22878
rect 15417 -22938 15477 -22878
rect 11 -23090 14 -23030
rect 14 -23090 66 -23030
rect 66 -23090 71 -23030
rect 331 -23090 391 -23030
rect 11 -23440 14 -23380
rect 14 -23440 66 -23380
rect 66 -23440 71 -23380
rect 331 -23440 391 -23380
rect 467 -23090 527 -23030
rect 787 -23090 847 -23030
rect 923 -23090 983 -23030
rect 1243 -23090 1303 -23030
rect 1381 -23090 1441 -23030
rect 1701 -23090 1761 -23030
rect 1837 -23090 1897 -23030
rect 2157 -23090 2217 -23030
rect 2293 -23090 2353 -23030
rect 2613 -23090 2673 -23030
rect 2751 -23090 2811 -23030
rect 3071 -23090 3131 -23030
rect 3207 -23090 3267 -23030
rect 3527 -23090 3587 -23030
rect 3663 -23090 3723 -23030
rect 3983 -23090 4043 -23030
rect 467 -23440 527 -23380
rect 787 -23440 847 -23380
rect 923 -23440 983 -23380
rect 1243 -23440 1303 -23380
rect 1381 -23440 1441 -23380
rect 1701 -23440 1761 -23380
rect 1837 -23440 1897 -23380
rect 2157 -23440 2217 -23380
rect 2293 -23440 2353 -23380
rect 2613 -23440 2673 -23380
rect 2751 -23440 2811 -23380
rect 3071 -23440 3131 -23380
rect 3207 -23440 3267 -23380
rect 3527 -23440 3587 -23380
rect 3663 -23440 3723 -23380
rect 3983 -23440 4043 -23380
rect 4121 -23090 4181 -23030
rect 4441 -23090 4501 -23030
rect 4577 -23090 4637 -23030
rect 4897 -23090 4957 -23030
rect 5033 -23090 5093 -23030
rect 5353 -23090 5413 -23030
rect 5491 -23090 5551 -23030
rect 5811 -23090 5871 -23030
rect 5947 -23090 6007 -23030
rect 6267 -23090 6327 -23030
rect 6403 -23090 6463 -23030
rect 6723 -23090 6783 -23030
rect 6861 -23090 6921 -23030
rect 7181 -23090 7241 -23030
rect 4121 -23440 4181 -23380
rect 4441 -23440 4501 -23380
rect 4577 -23440 4637 -23380
rect 4897 -23440 4957 -23380
rect 5033 -23440 5093 -23380
rect 5353 -23440 5413 -23380
rect 5491 -23440 5551 -23380
rect 5811 -23440 5871 -23380
rect 5947 -23440 6007 -23380
rect 6267 -23440 6327 -23380
rect 6403 -23440 6463 -23380
rect 6723 -23440 6783 -23380
rect 6861 -23440 6921 -23380
rect 7181 -23440 7241 -23380
rect 7317 -23090 7377 -23030
rect 7637 -23090 7697 -23030
rect 7773 -23090 7833 -23030
rect 8093 -23090 8153 -23030
rect 8247 -23090 8307 -23030
rect 8567 -23090 8627 -23030
rect 8703 -23090 8763 -23030
rect 9023 -23090 9083 -23030
rect 9161 -23090 9221 -23030
rect 9481 -23090 9541 -23030
rect 9617 -23090 9677 -23030
rect 9937 -23090 9997 -23030
rect 10073 -23090 10133 -23030
rect 10393 -23090 10453 -23030
rect 10531 -23090 10591 -23030
rect 10851 -23090 10911 -23030
rect 10987 -23090 11047 -23030
rect 11307 -23090 11367 -23030
rect 11443 -23090 11503 -23030
rect 11763 -23090 11823 -23030
rect 11901 -23090 11961 -23030
rect 12221 -23090 12281 -23030
rect 12357 -23090 12417 -23030
rect 12677 -23090 12737 -23030
rect 12813 -23090 12873 -23030
rect 13133 -23090 13193 -23030
rect 13271 -23090 13331 -23030
rect 13591 -23090 13651 -23030
rect 13727 -23090 13787 -23030
rect 14047 -23090 14107 -23030
rect 14183 -23090 14243 -23030
rect 14503 -23090 14563 -23030
rect 14641 -23090 14701 -23030
rect 14961 -23090 15021 -23030
rect 15097 -23090 15157 -23030
rect 15417 -23090 15477 -23030
rect 7317 -23440 7377 -23380
rect 7637 -23440 7697 -23380
rect 7773 -23440 7833 -23380
rect 8093 -23440 8153 -23380
rect 8247 -23440 8307 -23380
rect 8567 -23440 8627 -23380
rect 8703 -23440 8763 -23380
rect 9023 -23440 9083 -23380
rect 9161 -23440 9221 -23380
rect 9481 -23440 9541 -23380
rect 9617 -23440 9677 -23380
rect 9937 -23440 9997 -23380
rect 10073 -23440 10133 -23380
rect 10393 -23440 10453 -23380
rect 10531 -23440 10591 -23380
rect 10851 -23440 10911 -23380
rect 10987 -23440 11047 -23380
rect 11307 -23440 11367 -23380
rect 11443 -23440 11503 -23380
rect 11763 -23440 11823 -23380
rect 11901 -23440 11961 -23380
rect 12221 -23440 12281 -23380
rect 12357 -23440 12417 -23380
rect 12677 -23440 12737 -23380
rect 12813 -23440 12873 -23380
rect 13133 -23440 13193 -23380
rect 13271 -23440 13331 -23380
rect 13591 -23440 13651 -23380
rect 13727 -23440 13787 -23380
rect 14047 -23440 14107 -23380
rect 14183 -23440 14243 -23380
rect 14503 -23440 14563 -23380
rect 14641 -23440 14701 -23380
rect 14961 -23440 15021 -23380
rect 15097 -23440 15157 -23380
rect 15417 -23440 15477 -23380
rect 11 -23584 14 -23524
rect 14 -23584 66 -23524
rect 66 -23584 71 -23524
rect 331 -23584 391 -23524
rect 11 -23934 14 -23874
rect 14 -23934 66 -23874
rect 66 -23934 71 -23874
rect 331 -23934 391 -23874
rect 467 -23584 527 -23524
rect 787 -23584 847 -23524
rect 923 -23584 983 -23524
rect 1243 -23584 1303 -23524
rect 1381 -23584 1441 -23524
rect 1701 -23584 1761 -23524
rect 1837 -23584 1897 -23524
rect 2157 -23584 2217 -23524
rect 2293 -23584 2353 -23524
rect 2613 -23584 2673 -23524
rect 2751 -23584 2811 -23524
rect 3071 -23584 3131 -23524
rect 3207 -23584 3267 -23524
rect 3527 -23584 3587 -23524
rect 3663 -23584 3723 -23524
rect 3983 -23584 4043 -23524
rect 467 -23934 527 -23874
rect 787 -23934 847 -23874
rect 923 -23934 983 -23874
rect 1243 -23934 1303 -23874
rect 1381 -23934 1441 -23874
rect 1701 -23934 1761 -23874
rect 1837 -23934 1897 -23874
rect 2157 -23934 2217 -23874
rect 2293 -23934 2353 -23874
rect 2613 -23934 2673 -23874
rect 2751 -23934 2811 -23874
rect 3071 -23934 3131 -23874
rect 3207 -23934 3267 -23874
rect 3527 -23934 3587 -23874
rect 3663 -23934 3723 -23874
rect 3983 -23934 4043 -23874
rect 4121 -23584 4181 -23524
rect 4441 -23584 4501 -23524
rect 4577 -23584 4637 -23524
rect 4897 -23584 4957 -23524
rect 5033 -23584 5093 -23524
rect 5353 -23584 5413 -23524
rect 5491 -23584 5551 -23524
rect 5811 -23584 5871 -23524
rect 5947 -23584 6007 -23524
rect 6267 -23584 6327 -23524
rect 6403 -23584 6463 -23524
rect 6723 -23584 6783 -23524
rect 6861 -23584 6921 -23524
rect 7181 -23584 7241 -23524
rect 7317 -23584 7377 -23524
rect 7637 -23584 7697 -23524
rect 7773 -23584 7833 -23524
rect 8093 -23584 8153 -23524
rect 8247 -23584 8307 -23524
rect 8567 -23584 8627 -23524
rect 8703 -23584 8763 -23524
rect 9023 -23584 9083 -23524
rect 9161 -23584 9221 -23524
rect 9481 -23584 9541 -23524
rect 9617 -23584 9677 -23524
rect 9937 -23584 9997 -23524
rect 10073 -23584 10133 -23524
rect 10393 -23584 10453 -23524
rect 10531 -23584 10591 -23524
rect 10851 -23584 10911 -23524
rect 10987 -23584 11047 -23524
rect 11307 -23584 11367 -23524
rect 11443 -23584 11503 -23524
rect 11763 -23584 11823 -23524
rect 11901 -23584 11961 -23524
rect 12221 -23584 12281 -23524
rect 12357 -23584 12417 -23524
rect 12677 -23584 12737 -23524
rect 12813 -23584 12873 -23524
rect 13133 -23584 13193 -23524
rect 13271 -23584 13331 -23524
rect 13591 -23584 13651 -23524
rect 13727 -23584 13787 -23524
rect 14047 -23584 14107 -23524
rect 14183 -23584 14243 -23524
rect 14503 -23584 14563 -23524
rect 14641 -23584 14701 -23524
rect 14961 -23584 15021 -23524
rect 15097 -23584 15157 -23524
rect 15417 -23584 15477 -23524
rect 4121 -23934 4181 -23874
rect 4441 -23934 4501 -23874
rect 4577 -23934 4637 -23874
rect 4897 -23934 4957 -23874
rect 5033 -23934 5093 -23874
rect 5353 -23934 5413 -23874
rect 5491 -23934 5551 -23874
rect 5811 -23934 5871 -23874
rect 5947 -23934 6007 -23874
rect 6267 -23934 6327 -23874
rect 6403 -23934 6463 -23874
rect 6723 -23934 6783 -23874
rect 6861 -23934 6921 -23874
rect 7181 -23934 7241 -23874
rect 7317 -23934 7377 -23874
rect 7637 -23934 7697 -23874
rect 7773 -23934 7833 -23874
rect 8093 -23934 8153 -23874
rect 8247 -23934 8307 -23874
rect 8567 -23934 8627 -23874
rect 8703 -23934 8763 -23874
rect 9023 -23934 9083 -23874
rect 9161 -23934 9221 -23874
rect 9481 -23934 9541 -23874
rect 9617 -23934 9677 -23874
rect 9937 -23934 9997 -23874
rect 10073 -23934 10133 -23874
rect 10393 -23934 10453 -23874
rect 10531 -23934 10591 -23874
rect 10851 -23934 10911 -23874
rect 10987 -23934 11047 -23874
rect 11307 -23934 11367 -23874
rect 11443 -23934 11503 -23874
rect 11763 -23934 11823 -23874
rect 11901 -23934 11961 -23874
rect 12221 -23934 12281 -23874
rect 12357 -23934 12417 -23874
rect 12677 -23934 12737 -23874
rect 12813 -23934 12873 -23874
rect 13133 -23934 13193 -23874
rect 13271 -23934 13331 -23874
rect 13591 -23934 13651 -23874
rect 13727 -23934 13787 -23874
rect 14047 -23934 14107 -23874
rect 14183 -23934 14243 -23874
rect 14503 -23934 14563 -23874
rect 14641 -23934 14701 -23874
rect 14961 -23934 15021 -23874
rect 15097 -23934 15157 -23874
rect 15417 -23934 15477 -23874
rect 11 -24076 14 -24016
rect 14 -24076 66 -24016
rect 66 -24076 71 -24016
rect 331 -24076 391 -24016
rect 11 -24426 14 -24366
rect 14 -24426 66 -24366
rect 66 -24426 71 -24366
rect 331 -24426 391 -24366
rect 467 -24076 527 -24016
rect 787 -24076 847 -24016
rect 923 -24076 983 -24016
rect 1243 -24076 1303 -24016
rect 1381 -24076 1441 -24016
rect 1701 -24076 1761 -24016
rect 1837 -24076 1897 -24016
rect 2157 -24076 2217 -24016
rect 2293 -24076 2353 -24016
rect 2613 -24076 2673 -24016
rect 2751 -24076 2811 -24016
rect 3071 -24076 3131 -24016
rect 3207 -24076 3267 -24016
rect 3527 -24076 3587 -24016
rect 3663 -24076 3723 -24016
rect 3983 -24076 4043 -24016
rect 467 -24426 527 -24366
rect 787 -24426 847 -24366
rect 923 -24426 983 -24366
rect 1243 -24426 1303 -24366
rect 1381 -24426 1441 -24366
rect 1701 -24426 1761 -24366
rect 1837 -24426 1897 -24366
rect 2157 -24426 2217 -24366
rect 2293 -24426 2353 -24366
rect 2613 -24426 2673 -24366
rect 2751 -24426 2811 -24366
rect 3071 -24426 3131 -24366
rect 3207 -24426 3267 -24366
rect 3527 -24426 3587 -24366
rect 3663 -24426 3723 -24366
rect 3983 -24426 4043 -24366
rect 4121 -24076 4181 -24016
rect 4441 -24076 4501 -24016
rect 4577 -24076 4637 -24016
rect 4897 -24076 4957 -24016
rect 5033 -24076 5093 -24016
rect 5353 -24076 5413 -24016
rect 5491 -24076 5551 -24016
rect 5811 -24076 5871 -24016
rect 5947 -24076 6007 -24016
rect 6267 -24076 6327 -24016
rect 6403 -24076 6463 -24016
rect 6723 -24076 6783 -24016
rect 6861 -24076 6921 -24016
rect 7181 -24076 7241 -24016
rect 7317 -24076 7377 -24016
rect 7637 -24076 7697 -24016
rect 7773 -24076 7833 -24016
rect 8093 -24076 8153 -24016
rect 8247 -24076 8307 -24016
rect 8567 -24076 8627 -24016
rect 8703 -24076 8763 -24016
rect 9023 -24076 9083 -24016
rect 9161 -24076 9221 -24016
rect 9481 -24076 9541 -24016
rect 9617 -24076 9677 -24016
rect 9937 -24076 9997 -24016
rect 10073 -24076 10133 -24016
rect 10393 -24076 10453 -24016
rect 10531 -24076 10591 -24016
rect 10851 -24076 10911 -24016
rect 10987 -24076 11047 -24016
rect 11307 -24076 11367 -24016
rect 11443 -24076 11503 -24016
rect 11763 -24076 11823 -24016
rect 11901 -24076 11961 -24016
rect 12221 -24076 12281 -24016
rect 12357 -24076 12417 -24016
rect 12677 -24076 12737 -24016
rect 12813 -24076 12873 -24016
rect 13133 -24076 13193 -24016
rect 13271 -24076 13331 -24016
rect 13591 -24076 13651 -24016
rect 13727 -24076 13787 -24016
rect 14047 -24076 14107 -24016
rect 14183 -24076 14243 -24016
rect 14503 -24076 14563 -24016
rect 14641 -24076 14701 -24016
rect 14961 -24076 15021 -24016
rect 15097 -24076 15157 -24016
rect 15417 -24076 15477 -24016
rect 4121 -24426 4181 -24366
rect 4441 -24426 4501 -24366
rect 4577 -24426 4637 -24366
rect 4897 -24426 4957 -24366
rect 5033 -24426 5093 -24366
rect 5353 -24426 5413 -24366
rect 5491 -24426 5551 -24366
rect 5811 -24426 5871 -24366
rect 5947 -24426 6007 -24366
rect 6267 -24426 6327 -24366
rect 6403 -24426 6463 -24366
rect 6723 -24426 6783 -24366
rect 6861 -24426 6921 -24366
rect 7181 -24426 7241 -24366
rect 7317 -24426 7377 -24366
rect 7637 -24426 7697 -24366
rect 7773 -24426 7833 -24366
rect 8093 -24426 8153 -24366
rect 8247 -24426 8307 -24366
rect 8567 -24426 8627 -24366
rect 8703 -24426 8763 -24366
rect 9023 -24426 9083 -24366
rect 9161 -24426 9221 -24366
rect 9481 -24426 9541 -24366
rect 9617 -24426 9677 -24366
rect 9937 -24426 9997 -24366
rect 10073 -24426 10133 -24366
rect 10393 -24426 10453 -24366
rect 10531 -24426 10591 -24366
rect 10851 -24426 10911 -24366
rect 10987 -24426 11047 -24366
rect 11307 -24426 11367 -24366
rect 11443 -24426 11503 -24366
rect 11763 -24426 11823 -24366
rect 11901 -24426 11961 -24366
rect 12221 -24426 12281 -24366
rect 12357 -24426 12417 -24366
rect 12677 -24426 12737 -24366
rect 12813 -24426 12873 -24366
rect 13133 -24426 13193 -24366
rect 13271 -24426 13331 -24366
rect 13591 -24426 13651 -24366
rect 13727 -24426 13787 -24366
rect 14047 -24426 14107 -24366
rect 14183 -24426 14243 -24366
rect 14503 -24426 14563 -24366
rect 14641 -24426 14701 -24366
rect 14961 -24426 15021 -24366
rect 15097 -24426 15157 -24366
rect 15417 -24426 15477 -24366
rect 11 -24578 14 -24518
rect 14 -24578 66 -24518
rect 66 -24578 71 -24518
rect 331 -24578 391 -24518
rect 11 -24928 14 -24868
rect 14 -24928 66 -24868
rect 66 -24928 71 -24868
rect 331 -24928 391 -24868
rect 467 -24578 527 -24518
rect 787 -24578 847 -24518
rect 923 -24578 983 -24518
rect 1243 -24578 1303 -24518
rect 1381 -24578 1441 -24518
rect 1701 -24578 1761 -24518
rect 1837 -24578 1897 -24518
rect 2157 -24578 2217 -24518
rect 2293 -24578 2353 -24518
rect 2613 -24578 2673 -24518
rect 2751 -24578 2811 -24518
rect 3071 -24578 3131 -24518
rect 3207 -24578 3267 -24518
rect 3527 -24578 3587 -24518
rect 3663 -24578 3723 -24518
rect 3983 -24578 4043 -24518
rect 467 -24928 527 -24868
rect 787 -24928 847 -24868
rect 923 -24928 983 -24868
rect 1243 -24928 1303 -24868
rect 1381 -24928 1441 -24868
rect 1701 -24928 1761 -24868
rect 1837 -24928 1897 -24868
rect 2157 -24928 2217 -24868
rect 2293 -24928 2353 -24868
rect 2613 -24928 2673 -24868
rect 2751 -24928 2811 -24868
rect 3071 -24928 3131 -24868
rect 3207 -24928 3267 -24868
rect 3527 -24928 3587 -24868
rect 3663 -24928 3723 -24868
rect 3983 -24928 4043 -24868
rect 4121 -24578 4181 -24518
rect 4441 -24578 4501 -24518
rect 4577 -24578 4637 -24518
rect 4897 -24578 4957 -24518
rect 5033 -24578 5093 -24518
rect 5353 -24578 5413 -24518
rect 5491 -24578 5551 -24518
rect 5811 -24578 5871 -24518
rect 5947 -24578 6007 -24518
rect 6267 -24578 6327 -24518
rect 6403 -24578 6463 -24518
rect 6723 -24578 6783 -24518
rect 6861 -24578 6921 -24518
rect 7181 -24578 7241 -24518
rect 7317 -24578 7377 -24518
rect 7637 -24578 7697 -24518
rect 7773 -24578 7833 -24518
rect 8093 -24578 8153 -24518
rect 8247 -24578 8307 -24518
rect 8567 -24578 8627 -24518
rect 8703 -24578 8763 -24518
rect 9023 -24578 9083 -24518
rect 9161 -24578 9221 -24518
rect 9481 -24578 9541 -24518
rect 9617 -24578 9677 -24518
rect 9937 -24578 9997 -24518
rect 10073 -24578 10133 -24518
rect 10393 -24578 10453 -24518
rect 10531 -24578 10591 -24518
rect 10851 -24578 10911 -24518
rect 10987 -24578 11047 -24518
rect 11307 -24578 11367 -24518
rect 11443 -24578 11503 -24518
rect 11763 -24578 11823 -24518
rect 11901 -24578 11961 -24518
rect 12221 -24578 12281 -24518
rect 12357 -24578 12417 -24518
rect 12677 -24578 12737 -24518
rect 12813 -24578 12873 -24518
rect 13133 -24578 13193 -24518
rect 13271 -24578 13331 -24518
rect 13591 -24578 13651 -24518
rect 13727 -24578 13787 -24518
rect 14047 -24578 14107 -24518
rect 14183 -24578 14243 -24518
rect 14503 -24578 14563 -24518
rect 14641 -24578 14701 -24518
rect 14961 -24578 15021 -24518
rect 15097 -24578 15157 -24518
rect 15417 -24578 15477 -24518
rect 4121 -24928 4181 -24868
rect 4441 -24928 4501 -24868
rect 4577 -24928 4637 -24868
rect 4897 -24928 4957 -24868
rect 5033 -24928 5093 -24868
rect 5353 -24928 5413 -24868
rect 5491 -24928 5551 -24868
rect 5811 -24928 5871 -24868
rect 5947 -24928 6007 -24868
rect 6267 -24928 6327 -24868
rect 6403 -24928 6463 -24868
rect 6723 -24928 6783 -24868
rect 6861 -24928 6921 -24868
rect 7181 -24928 7241 -24868
rect 7317 -24928 7377 -24868
rect 7637 -24928 7697 -24868
rect 7773 -24928 7833 -24868
rect 8093 -24928 8153 -24868
rect 8247 -24928 8307 -24868
rect 8567 -24928 8627 -24868
rect 8703 -24928 8763 -24868
rect 9023 -24928 9083 -24868
rect 9161 -24928 9221 -24868
rect 9481 -24928 9541 -24868
rect 9617 -24928 9677 -24868
rect 9937 -24928 9997 -24868
rect 10073 -24928 10133 -24868
rect 10393 -24928 10453 -24868
rect 10531 -24928 10591 -24868
rect 10851 -24928 10911 -24868
rect 10987 -24928 11047 -24868
rect 11307 -24928 11367 -24868
rect 11443 -24928 11503 -24868
rect 11763 -24928 11823 -24868
rect 11901 -24928 11961 -24868
rect 12221 -24928 12281 -24868
rect 12357 -24928 12417 -24868
rect 12677 -24928 12737 -24868
rect 12813 -24928 12873 -24868
rect 13133 -24928 13193 -24868
rect 13271 -24928 13331 -24868
rect 13591 -24928 13651 -24868
rect 13727 -24928 13787 -24868
rect 14047 -24928 14107 -24868
rect 14183 -24928 14243 -24868
rect 14503 -24928 14563 -24868
rect 14641 -24928 14701 -24868
rect 14961 -24928 15021 -24868
rect 15097 -24928 15157 -24868
rect 15417 -24928 15477 -24868
rect 11 -25094 14 -25034
rect 14 -25094 66 -25034
rect 66 -25094 71 -25034
rect 331 -25094 391 -25034
rect 11 -25444 14 -25384
rect 14 -25444 66 -25384
rect 66 -25444 71 -25384
rect 331 -25444 391 -25384
rect 467 -25094 527 -25034
rect 787 -25094 847 -25034
rect 923 -25094 983 -25034
rect 1243 -25094 1303 -25034
rect 1381 -25094 1441 -25034
rect 1701 -25094 1761 -25034
rect 1837 -25094 1897 -25034
rect 2157 -25094 2217 -25034
rect 2293 -25094 2353 -25034
rect 2613 -25094 2673 -25034
rect 2751 -25094 2811 -25034
rect 3071 -25094 3131 -25034
rect 3207 -25094 3267 -25034
rect 3527 -25094 3587 -25034
rect 3663 -25094 3723 -25034
rect 3983 -25094 4043 -25034
rect 467 -25444 527 -25384
rect 787 -25444 847 -25384
rect 923 -25444 983 -25384
rect 1243 -25444 1303 -25384
rect 1381 -25444 1441 -25384
rect 1701 -25444 1761 -25384
rect 1837 -25444 1897 -25384
rect 2157 -25444 2217 -25384
rect 2293 -25444 2353 -25384
rect 2613 -25444 2673 -25384
rect 2751 -25444 2811 -25384
rect 3071 -25444 3131 -25384
rect 3207 -25444 3267 -25384
rect 3527 -25444 3587 -25384
rect 3663 -25444 3723 -25384
rect 3983 -25444 4043 -25384
rect 4121 -25094 4181 -25034
rect 4441 -25094 4501 -25034
rect 4577 -25094 4637 -25034
rect 4897 -25094 4957 -25034
rect 5033 -25094 5093 -25034
rect 5353 -25094 5413 -25034
rect 5491 -25094 5551 -25034
rect 5811 -25094 5871 -25034
rect 5947 -25094 6007 -25034
rect 6267 -25094 6327 -25034
rect 6403 -25094 6463 -25034
rect 6723 -25094 6783 -25034
rect 6861 -25094 6921 -25034
rect 7181 -25094 7241 -25034
rect 7317 -25094 7377 -25034
rect 7637 -25094 7697 -25034
rect 7773 -25094 7833 -25034
rect 8093 -25094 8153 -25034
rect 8247 -25094 8307 -25034
rect 8567 -25094 8627 -25034
rect 8703 -25094 8763 -25034
rect 9023 -25094 9083 -25034
rect 9161 -25094 9221 -25034
rect 9481 -25094 9541 -25034
rect 9617 -25094 9677 -25034
rect 9937 -25094 9997 -25034
rect 10073 -25094 10133 -25034
rect 10393 -25094 10453 -25034
rect 10531 -25094 10591 -25034
rect 10851 -25094 10911 -25034
rect 10987 -25094 11047 -25034
rect 11307 -25094 11367 -25034
rect 11443 -25094 11503 -25034
rect 11763 -25094 11823 -25034
rect 11901 -25094 11961 -25034
rect 12221 -25094 12281 -25034
rect 12357 -25094 12417 -25034
rect 12677 -25094 12737 -25034
rect 12813 -25094 12873 -25034
rect 13133 -25094 13193 -25034
rect 13271 -25094 13331 -25034
rect 13591 -25094 13651 -25034
rect 13727 -25094 13787 -25034
rect 14047 -25094 14107 -25034
rect 14183 -25094 14243 -25034
rect 14503 -25094 14563 -25034
rect 14641 -25094 14701 -25034
rect 14961 -25094 15021 -25034
rect 15097 -25094 15157 -25034
rect 15417 -25094 15477 -25034
rect 4121 -25444 4181 -25384
rect 4441 -25444 4501 -25384
rect 4577 -25444 4637 -25384
rect 4897 -25444 4957 -25384
rect 5033 -25444 5093 -25384
rect 5353 -25444 5413 -25384
rect 5491 -25444 5551 -25384
rect 5811 -25444 5871 -25384
rect 5947 -25444 6007 -25384
rect 6267 -25444 6327 -25384
rect 6403 -25444 6463 -25384
rect 6723 -25444 6783 -25384
rect 6861 -25444 6921 -25384
rect 7181 -25444 7241 -25384
rect 7317 -25444 7377 -25384
rect 7637 -25444 7697 -25384
rect 7773 -25444 7833 -25384
rect 8093 -25444 8153 -25384
rect 8247 -25444 8307 -25384
rect 8567 -25444 8627 -25384
rect 8703 -25444 8763 -25384
rect 9023 -25444 9083 -25384
rect 9161 -25444 9221 -25384
rect 9481 -25444 9541 -25384
rect 9617 -25444 9677 -25384
rect 9937 -25444 9997 -25384
rect 10073 -25444 10133 -25384
rect 10393 -25444 10453 -25384
rect 10531 -25444 10591 -25384
rect 10851 -25444 10911 -25384
rect 10987 -25444 11047 -25384
rect 11307 -25444 11367 -25384
rect 11443 -25444 11503 -25384
rect 11763 -25444 11823 -25384
rect 11901 -25444 11961 -25384
rect 12221 -25444 12281 -25384
rect 12357 -25444 12417 -25384
rect 12677 -25444 12737 -25384
rect 12813 -25444 12873 -25384
rect 13133 -25444 13193 -25384
rect 13271 -25444 13331 -25384
rect 13591 -25444 13651 -25384
rect 13727 -25444 13787 -25384
rect 14047 -25444 14107 -25384
rect 14183 -25444 14243 -25384
rect 14503 -25444 14563 -25384
rect 14641 -25444 14701 -25384
rect 14961 -25444 15021 -25384
rect 15097 -25444 15157 -25384
rect 15417 -25444 15477 -25384
rect 11 -25586 14 -25526
rect 14 -25586 66 -25526
rect 66 -25586 71 -25526
rect 331 -25586 391 -25526
rect 11 -25936 14 -25876
rect 14 -25936 66 -25876
rect 66 -25936 71 -25876
rect 331 -25936 391 -25876
rect 467 -25586 527 -25526
rect 787 -25586 847 -25526
rect 923 -25586 983 -25526
rect 1243 -25586 1303 -25526
rect 1381 -25586 1441 -25526
rect 1701 -25586 1761 -25526
rect 1837 -25586 1897 -25526
rect 2157 -25586 2217 -25526
rect 2293 -25586 2353 -25526
rect 2613 -25586 2673 -25526
rect 2751 -25586 2811 -25526
rect 3071 -25586 3131 -25526
rect 3207 -25586 3267 -25526
rect 3527 -25586 3587 -25526
rect 3663 -25586 3723 -25526
rect 3983 -25586 4043 -25526
rect 467 -25936 527 -25876
rect 787 -25936 847 -25876
rect 923 -25936 983 -25876
rect 1243 -25936 1303 -25876
rect 1381 -25936 1441 -25876
rect 1701 -25936 1761 -25876
rect 1837 -25936 1897 -25876
rect 2157 -25936 2217 -25876
rect 2293 -25936 2353 -25876
rect 2613 -25936 2673 -25876
rect 2751 -25936 2811 -25876
rect 3071 -25936 3131 -25876
rect 3207 -25936 3267 -25876
rect 3527 -25936 3587 -25876
rect 3663 -25936 3723 -25876
rect 3983 -25936 4043 -25876
rect 4121 -25586 4181 -25526
rect 4441 -25586 4501 -25526
rect 4577 -25586 4637 -25526
rect 4897 -25586 4957 -25526
rect 5033 -25586 5093 -25526
rect 5353 -25586 5413 -25526
rect 5491 -25586 5551 -25526
rect 5811 -25586 5871 -25526
rect 5947 -25586 6007 -25526
rect 6267 -25586 6327 -25526
rect 6403 -25586 6463 -25526
rect 6723 -25586 6783 -25526
rect 6861 -25586 6921 -25526
rect 7181 -25586 7241 -25526
rect 7317 -25586 7377 -25526
rect 7637 -25586 7697 -25526
rect 7773 -25586 7833 -25526
rect 8093 -25586 8153 -25526
rect 8247 -25586 8307 -25526
rect 8567 -25586 8627 -25526
rect 8703 -25586 8763 -25526
rect 9023 -25586 9083 -25526
rect 9161 -25586 9221 -25526
rect 9481 -25586 9541 -25526
rect 9617 -25586 9677 -25526
rect 9937 -25586 9997 -25526
rect 10073 -25586 10133 -25526
rect 10393 -25586 10453 -25526
rect 10531 -25586 10591 -25526
rect 10851 -25586 10911 -25526
rect 10987 -25586 11047 -25526
rect 11307 -25586 11367 -25526
rect 11443 -25586 11503 -25526
rect 11763 -25586 11823 -25526
rect 11901 -25586 11961 -25526
rect 12221 -25586 12281 -25526
rect 12357 -25586 12417 -25526
rect 12677 -25586 12737 -25526
rect 12813 -25586 12873 -25526
rect 13133 -25586 13193 -25526
rect 13271 -25586 13331 -25526
rect 13591 -25586 13651 -25526
rect 13727 -25586 13787 -25526
rect 14047 -25586 14107 -25526
rect 14183 -25586 14243 -25526
rect 14503 -25586 14563 -25526
rect 14641 -25586 14701 -25526
rect 14961 -25586 15021 -25526
rect 15097 -25586 15157 -25526
rect 15417 -25586 15477 -25526
rect 4121 -25936 4181 -25876
rect 4441 -25936 4501 -25876
rect 4577 -25936 4637 -25876
rect 4897 -25936 4957 -25876
rect 5033 -25936 5093 -25876
rect 5353 -25936 5413 -25876
rect 5491 -25936 5551 -25876
rect 5811 -25936 5871 -25876
rect 5947 -25936 6007 -25876
rect 6267 -25936 6327 -25876
rect 6403 -25936 6463 -25876
rect 6723 -25936 6783 -25876
rect 6861 -25936 6921 -25876
rect 7181 -25936 7241 -25876
rect 7317 -25936 7377 -25876
rect 7637 -25936 7697 -25876
rect 7773 -25936 7833 -25876
rect 8093 -25936 8153 -25876
rect 8247 -25936 8307 -25876
rect 8567 -25936 8627 -25876
rect 8703 -25936 8763 -25876
rect 9023 -25936 9083 -25876
rect 9161 -25936 9221 -25876
rect 9481 -25936 9541 -25876
rect 9617 -25936 9677 -25876
rect 9937 -25936 9997 -25876
rect 10073 -25936 10133 -25876
rect 10393 -25936 10453 -25876
rect 10531 -25936 10591 -25876
rect 10851 -25936 10911 -25876
rect 10987 -25936 11047 -25876
rect 11307 -25936 11367 -25876
rect 11443 -25936 11503 -25876
rect 11763 -25936 11823 -25876
rect 11901 -25936 11961 -25876
rect 12221 -25936 12281 -25876
rect 12357 -25936 12417 -25876
rect 12677 -25936 12737 -25876
rect 12813 -25936 12873 -25876
rect 13133 -25936 13193 -25876
rect 13271 -25936 13331 -25876
rect 13591 -25936 13651 -25876
rect 13727 -25936 13787 -25876
rect 14047 -25936 14107 -25876
rect 14183 -25936 14243 -25876
rect 14503 -25936 14563 -25876
rect 14641 -25936 14701 -25876
rect 14961 -25936 15021 -25876
rect 15097 -25936 15157 -25876
rect 15417 -25936 15477 -25876
rect 10 -26083 14 -26023
rect 14 -26083 66 -26023
rect 66 -26083 70 -26023
rect 330 -26083 390 -26023
rect 10 -26433 14 -26373
rect 14 -26433 66 -26373
rect 66 -26433 70 -26373
rect 330 -26433 390 -26373
rect 466 -26083 526 -26023
rect 786 -26083 846 -26023
rect 922 -26083 982 -26023
rect 1242 -26083 1302 -26023
rect 1380 -26083 1440 -26023
rect 1700 -26083 1760 -26023
rect 1836 -26083 1896 -26023
rect 2156 -26083 2216 -26023
rect 2292 -26083 2352 -26023
rect 2612 -26083 2672 -26023
rect 2750 -26083 2810 -26023
rect 3070 -26083 3130 -26023
rect 3206 -26083 3266 -26023
rect 3526 -26083 3586 -26023
rect 3662 -26083 3722 -26023
rect 3982 -26083 4042 -26023
rect 466 -26433 526 -26373
rect 786 -26433 846 -26373
rect 922 -26433 982 -26373
rect 1242 -26433 1302 -26373
rect 1380 -26433 1440 -26373
rect 1700 -26433 1760 -26373
rect 1836 -26433 1896 -26373
rect 2156 -26433 2216 -26373
rect 2292 -26433 2352 -26373
rect 2612 -26433 2672 -26373
rect 2750 -26433 2810 -26373
rect 3070 -26433 3130 -26373
rect 3206 -26433 3266 -26373
rect 3526 -26433 3586 -26373
rect 3662 -26433 3722 -26373
rect 3982 -26433 4042 -26373
rect 4120 -26083 4180 -26023
rect 4440 -26083 4500 -26023
rect 4576 -26083 4636 -26023
rect 4896 -26083 4956 -26023
rect 5032 -26083 5092 -26023
rect 5352 -26083 5412 -26023
rect 5490 -26083 5550 -26023
rect 5810 -26083 5870 -26023
rect 5946 -26083 6006 -26023
rect 6266 -26083 6326 -26023
rect 6402 -26083 6462 -26023
rect 6722 -26083 6782 -26023
rect 6860 -26083 6920 -26023
rect 7180 -26083 7240 -26023
rect 7316 -26083 7376 -26023
rect 7636 -26083 7696 -26023
rect 7772 -26083 7832 -26023
rect 8092 -26083 8152 -26023
rect 8246 -26083 8306 -26023
rect 8566 -26083 8626 -26023
rect 8702 -26083 8762 -26023
rect 9022 -26083 9082 -26023
rect 9160 -26083 9220 -26023
rect 9480 -26083 9540 -26023
rect 9616 -26083 9676 -26023
rect 9936 -26083 9996 -26023
rect 10072 -26083 10132 -26023
rect 10392 -26083 10452 -26023
rect 10530 -26083 10590 -26023
rect 10850 -26083 10910 -26023
rect 10986 -26083 11046 -26023
rect 11306 -26083 11366 -26023
rect 11442 -26083 11502 -26023
rect 11762 -26083 11822 -26023
rect 11900 -26083 11960 -26023
rect 12220 -26083 12280 -26023
rect 12356 -26083 12416 -26023
rect 12676 -26083 12736 -26023
rect 12812 -26083 12872 -26023
rect 13132 -26083 13192 -26023
rect 13270 -26083 13330 -26023
rect 13590 -26083 13650 -26023
rect 13726 -26083 13786 -26023
rect 14046 -26083 14106 -26023
rect 14182 -26083 14242 -26023
rect 14502 -26083 14562 -26023
rect 14640 -26083 14700 -26023
rect 14960 -26083 15020 -26023
rect 15096 -26083 15156 -26023
rect 15416 -26083 15476 -26023
rect 4120 -26433 4180 -26373
rect 4440 -26433 4500 -26373
rect 4576 -26433 4636 -26373
rect 4896 -26433 4956 -26373
rect 5032 -26433 5092 -26373
rect 5352 -26433 5412 -26373
rect 5490 -26433 5550 -26373
rect 5810 -26433 5870 -26373
rect 5946 -26433 6006 -26373
rect 6266 -26433 6326 -26373
rect 6402 -26433 6462 -26373
rect 6722 -26433 6782 -26373
rect 6860 -26433 6920 -26373
rect 7180 -26433 7240 -26373
rect 7316 -26433 7376 -26373
rect 7636 -26433 7696 -26373
rect 7772 -26433 7832 -26373
rect 8092 -26433 8152 -26373
rect 8246 -26433 8306 -26373
rect 8566 -26433 8626 -26373
rect 8702 -26433 8762 -26373
rect 9022 -26433 9082 -26373
rect 9160 -26433 9220 -26373
rect 9480 -26433 9540 -26373
rect 9616 -26433 9676 -26373
rect 9936 -26433 9996 -26373
rect 10072 -26433 10132 -26373
rect 10392 -26433 10452 -26373
rect 10530 -26433 10590 -26373
rect 10850 -26433 10910 -26373
rect 10986 -26433 11046 -26373
rect 11306 -26433 11366 -26373
rect 11442 -26433 11502 -26373
rect 11762 -26433 11822 -26373
rect 11900 -26433 11960 -26373
rect 12220 -26433 12280 -26373
rect 12356 -26433 12416 -26373
rect 12676 -26433 12736 -26373
rect 12812 -26433 12872 -26373
rect 13132 -26433 13192 -26373
rect 13270 -26433 13330 -26373
rect 13590 -26433 13650 -26373
rect 13726 -26433 13786 -26373
rect 14046 -26433 14106 -26373
rect 14182 -26433 14242 -26373
rect 14502 -26433 14562 -26373
rect 14640 -26433 14700 -26373
rect 14960 -26433 15020 -26373
rect 15096 -26433 15156 -26373
rect 15416 -26433 15476 -26373
rect 10 -26575 14 -26515
rect 14 -26575 66 -26515
rect 66 -26575 70 -26515
rect 330 -26575 390 -26515
rect 10 -26925 14 -26865
rect 14 -26925 66 -26865
rect 66 -26925 70 -26865
rect 330 -26925 390 -26865
rect 466 -26575 526 -26515
rect 786 -26575 846 -26515
rect 922 -26575 982 -26515
rect 1242 -26575 1302 -26515
rect 1380 -26575 1440 -26515
rect 1700 -26575 1760 -26515
rect 1836 -26575 1896 -26515
rect 2156 -26575 2216 -26515
rect 2292 -26575 2352 -26515
rect 2612 -26575 2672 -26515
rect 2750 -26575 2810 -26515
rect 3070 -26575 3130 -26515
rect 3206 -26575 3266 -26515
rect 3526 -26575 3586 -26515
rect 3662 -26575 3722 -26515
rect 3982 -26575 4042 -26515
rect 4120 -26575 4180 -26515
rect 4440 -26575 4500 -26515
rect 4576 -26575 4636 -26515
rect 4896 -26575 4956 -26515
rect 5032 -26575 5092 -26515
rect 5352 -26575 5412 -26515
rect 5490 -26575 5550 -26515
rect 5810 -26575 5870 -26515
rect 5946 -26575 6006 -26515
rect 6266 -26575 6326 -26515
rect 6402 -26575 6462 -26515
rect 6722 -26575 6782 -26515
rect 6860 -26575 6920 -26515
rect 7180 -26575 7240 -26515
rect 7316 -26575 7376 -26515
rect 7636 -26575 7696 -26515
rect 7772 -26575 7832 -26515
rect 8092 -26575 8152 -26515
rect 8246 -26575 8306 -26515
rect 8566 -26575 8626 -26515
rect 8702 -26575 8762 -26515
rect 9022 -26575 9082 -26515
rect 9160 -26575 9220 -26515
rect 9480 -26575 9540 -26515
rect 9616 -26575 9676 -26515
rect 9936 -26575 9996 -26515
rect 10072 -26575 10132 -26515
rect 10392 -26575 10452 -26515
rect 10530 -26575 10590 -26515
rect 10850 -26575 10910 -26515
rect 10986 -26575 11046 -26515
rect 11306 -26575 11366 -26515
rect 11442 -26575 11502 -26515
rect 11762 -26575 11822 -26515
rect 11900 -26575 11960 -26515
rect 12220 -26575 12280 -26515
rect 12356 -26575 12416 -26515
rect 12676 -26575 12736 -26515
rect 12812 -26575 12872 -26515
rect 13132 -26575 13192 -26515
rect 13270 -26575 13330 -26515
rect 13590 -26575 13650 -26515
rect 13726 -26575 13786 -26515
rect 14046 -26575 14106 -26515
rect 14182 -26575 14242 -26515
rect 14502 -26575 14562 -26515
rect 14640 -26575 14700 -26515
rect 14960 -26575 15020 -26515
rect 15096 -26575 15156 -26515
rect 15416 -26575 15476 -26515
rect 466 -26925 526 -26865
rect 786 -26925 846 -26865
rect 922 -26925 982 -26865
rect 1242 -26925 1302 -26865
rect 1380 -26925 1440 -26865
rect 1700 -26925 1760 -26865
rect 1836 -26925 1896 -26865
rect 2156 -26925 2216 -26865
rect 2292 -26925 2352 -26865
rect 2612 -26925 2672 -26865
rect 2750 -26925 2810 -26865
rect 3070 -26925 3130 -26865
rect 3206 -26925 3266 -26865
rect 3526 -26925 3586 -26865
rect 3662 -26925 3722 -26865
rect 3982 -26925 4042 -26865
rect 4120 -26925 4180 -26865
rect 4440 -26925 4500 -26865
rect 4576 -26925 4636 -26865
rect 4896 -26925 4956 -26865
rect 5032 -26925 5092 -26865
rect 5352 -26925 5412 -26865
rect 5490 -26925 5550 -26865
rect 5810 -26925 5870 -26865
rect 5946 -26925 6006 -26865
rect 6266 -26925 6326 -26865
rect 6402 -26925 6462 -26865
rect 6722 -26925 6782 -26865
rect 6860 -26925 6920 -26865
rect 7180 -26925 7240 -26865
rect 7316 -26925 7376 -26865
rect 7636 -26925 7696 -26865
rect 7772 -26925 7832 -26865
rect 8092 -26925 8152 -26865
rect 8246 -26925 8306 -26865
rect 8566 -26925 8626 -26865
rect 8702 -26925 8762 -26865
rect 9022 -26925 9082 -26865
rect 9160 -26925 9220 -26865
rect 9480 -26925 9540 -26865
rect 9616 -26925 9676 -26865
rect 9936 -26925 9996 -26865
rect 10072 -26925 10132 -26865
rect 10392 -26925 10452 -26865
rect 10530 -26925 10590 -26865
rect 10850 -26925 10910 -26865
rect 10986 -26925 11046 -26865
rect 11306 -26925 11366 -26865
rect 11442 -26925 11502 -26865
rect 11762 -26925 11822 -26865
rect 11900 -26925 11960 -26865
rect 12220 -26925 12280 -26865
rect 12356 -26925 12416 -26865
rect 12676 -26925 12736 -26865
rect 12812 -26925 12872 -26865
rect 13132 -26925 13192 -26865
rect 13270 -26925 13330 -26865
rect 13590 -26925 13650 -26865
rect 13726 -26925 13786 -26865
rect 14046 -26925 14106 -26865
rect 14182 -26925 14242 -26865
rect 14502 -26925 14562 -26865
rect 14640 -26925 14700 -26865
rect 14960 -26925 15020 -26865
rect 15096 -26925 15156 -26865
rect 15416 -26925 15476 -26865
rect 10 -27077 14 -27017
rect 14 -27077 66 -27017
rect 66 -27077 70 -27017
rect 330 -27077 390 -27017
rect 10 -27427 14 -27367
rect 14 -27427 66 -27367
rect 66 -27427 70 -27367
rect 330 -27427 390 -27367
rect 466 -27077 526 -27017
rect 786 -27077 846 -27017
rect 922 -27077 982 -27017
rect 1242 -27077 1302 -27017
rect 1380 -27077 1440 -27017
rect 1700 -27077 1760 -27017
rect 1836 -27077 1896 -27017
rect 2156 -27077 2216 -27017
rect 2292 -27077 2352 -27017
rect 2612 -27077 2672 -27017
rect 2750 -27077 2810 -27017
rect 3070 -27077 3130 -27017
rect 3206 -27077 3266 -27017
rect 3526 -27077 3586 -27017
rect 3662 -27077 3722 -27017
rect 3982 -27077 4042 -27017
rect 4120 -27077 4180 -27017
rect 4440 -27077 4500 -27017
rect 4576 -27077 4636 -27017
rect 4896 -27077 4956 -27017
rect 5032 -27077 5092 -27017
rect 5352 -27077 5412 -27017
rect 5490 -27077 5550 -27017
rect 5810 -27077 5870 -27017
rect 5946 -27077 6006 -27017
rect 6266 -27077 6326 -27017
rect 6402 -27077 6462 -27017
rect 6722 -27077 6782 -27017
rect 6860 -27077 6920 -27017
rect 7180 -27077 7240 -27017
rect 7316 -27077 7376 -27017
rect 7636 -27077 7696 -27017
rect 7772 -27077 7832 -27017
rect 8092 -27077 8152 -27017
rect 8246 -27077 8306 -27017
rect 8566 -27077 8626 -27017
rect 8702 -27077 8762 -27017
rect 9022 -27077 9082 -27017
rect 9160 -27077 9220 -27017
rect 9480 -27077 9540 -27017
rect 9616 -27077 9676 -27017
rect 9936 -27077 9996 -27017
rect 10072 -27077 10132 -27017
rect 10392 -27077 10452 -27017
rect 10530 -27077 10590 -27017
rect 10850 -27077 10910 -27017
rect 10986 -27077 11046 -27017
rect 11306 -27077 11366 -27017
rect 11442 -27077 11502 -27017
rect 11762 -27077 11822 -27017
rect 11900 -27077 11960 -27017
rect 12220 -27077 12280 -27017
rect 12356 -27077 12416 -27017
rect 12676 -27077 12736 -27017
rect 12812 -27077 12872 -27017
rect 13132 -27077 13192 -27017
rect 13270 -27077 13330 -27017
rect 13590 -27077 13650 -27017
rect 13726 -27077 13786 -27017
rect 14046 -27077 14106 -27017
rect 14182 -27077 14242 -27017
rect 14502 -27077 14562 -27017
rect 14640 -27077 14700 -27017
rect 14960 -27077 15020 -27017
rect 15096 -27077 15156 -27017
rect 15416 -27077 15476 -27017
rect 466 -27427 526 -27367
rect 786 -27427 846 -27367
rect 922 -27427 982 -27367
rect 1242 -27427 1302 -27367
rect 1380 -27427 1440 -27367
rect 1700 -27427 1760 -27367
rect 1836 -27427 1896 -27367
rect 2156 -27427 2216 -27367
rect 2292 -27427 2352 -27367
rect 2612 -27427 2672 -27367
rect 2750 -27427 2810 -27367
rect 3070 -27427 3130 -27367
rect 3206 -27427 3266 -27367
rect 3526 -27427 3586 -27367
rect 3662 -27427 3722 -27367
rect 3982 -27427 4042 -27367
rect 4120 -27427 4180 -27367
rect 4440 -27427 4500 -27367
rect 4576 -27427 4636 -27367
rect 4896 -27427 4956 -27367
rect 5032 -27427 5092 -27367
rect 5352 -27427 5412 -27367
rect 5490 -27427 5550 -27367
rect 5810 -27427 5870 -27367
rect 5946 -27427 6006 -27367
rect 6266 -27427 6326 -27367
rect 6402 -27427 6462 -27367
rect 6722 -27427 6782 -27367
rect 6860 -27427 6920 -27367
rect 7180 -27427 7240 -27367
rect 7316 -27427 7376 -27367
rect 7636 -27427 7696 -27367
rect 7772 -27427 7832 -27367
rect 8092 -27427 8152 -27367
rect 8246 -27427 8306 -27367
rect 8566 -27427 8626 -27367
rect 8702 -27427 8762 -27367
rect 9022 -27427 9082 -27367
rect 9160 -27427 9220 -27367
rect 9480 -27427 9540 -27367
rect 9616 -27427 9676 -27367
rect 9936 -27427 9996 -27367
rect 10072 -27427 10132 -27367
rect 10392 -27427 10452 -27367
rect 10530 -27427 10590 -27367
rect 10850 -27427 10910 -27367
rect 10986 -27427 11046 -27367
rect 11306 -27427 11366 -27367
rect 11442 -27427 11502 -27367
rect 11762 -27427 11822 -27367
rect 11900 -27427 11960 -27367
rect 12220 -27427 12280 -27367
rect 12356 -27427 12416 -27367
rect 12676 -27427 12736 -27367
rect 12812 -27427 12872 -27367
rect 13132 -27427 13192 -27367
rect 13270 -27427 13330 -27367
rect 13590 -27427 13650 -27367
rect 13726 -27427 13786 -27367
rect 14046 -27427 14106 -27367
rect 14182 -27427 14242 -27367
rect 14502 -27427 14562 -27367
rect 14640 -27427 14700 -27367
rect 14960 -27427 15020 -27367
rect 15096 -27427 15156 -27367
rect 15416 -27427 15476 -27367
rect 10 -27593 14 -27533
rect 14 -27593 66 -27533
rect 66 -27593 70 -27533
rect 330 -27593 390 -27533
rect 10 -27943 14 -27883
rect 14 -27943 66 -27883
rect 66 -27943 70 -27883
rect 330 -27943 390 -27883
rect 466 -27593 526 -27533
rect 786 -27593 846 -27533
rect 922 -27593 982 -27533
rect 1242 -27593 1302 -27533
rect 1380 -27593 1440 -27533
rect 1700 -27593 1760 -27533
rect 1836 -27593 1896 -27533
rect 2156 -27593 2216 -27533
rect 2292 -27593 2352 -27533
rect 2612 -27593 2672 -27533
rect 2750 -27593 2810 -27533
rect 3070 -27593 3130 -27533
rect 3206 -27593 3266 -27533
rect 3526 -27593 3586 -27533
rect 3662 -27593 3722 -27533
rect 3982 -27593 4042 -27533
rect 4120 -27593 4180 -27533
rect 4440 -27593 4500 -27533
rect 4576 -27593 4636 -27533
rect 4896 -27593 4956 -27533
rect 5032 -27593 5092 -27533
rect 5352 -27593 5412 -27533
rect 5490 -27593 5550 -27533
rect 5810 -27593 5870 -27533
rect 5946 -27593 6006 -27533
rect 6266 -27593 6326 -27533
rect 6402 -27593 6462 -27533
rect 6722 -27593 6782 -27533
rect 6860 -27593 6920 -27533
rect 7180 -27593 7240 -27533
rect 7316 -27593 7376 -27533
rect 7636 -27593 7696 -27533
rect 7772 -27593 7832 -27533
rect 8092 -27593 8152 -27533
rect 8246 -27593 8306 -27533
rect 8566 -27593 8626 -27533
rect 8702 -27593 8762 -27533
rect 9022 -27593 9082 -27533
rect 9160 -27593 9220 -27533
rect 9480 -27593 9540 -27533
rect 9616 -27593 9676 -27533
rect 9936 -27593 9996 -27533
rect 10072 -27593 10132 -27533
rect 10392 -27593 10452 -27533
rect 10530 -27593 10590 -27533
rect 10850 -27593 10910 -27533
rect 10986 -27593 11046 -27533
rect 11306 -27593 11366 -27533
rect 11442 -27593 11502 -27533
rect 11762 -27593 11822 -27533
rect 11900 -27593 11960 -27533
rect 12220 -27593 12280 -27533
rect 12356 -27593 12416 -27533
rect 12676 -27593 12736 -27533
rect 12812 -27593 12872 -27533
rect 13132 -27593 13192 -27533
rect 13270 -27593 13330 -27533
rect 13590 -27593 13650 -27533
rect 13726 -27593 13786 -27533
rect 14046 -27593 14106 -27533
rect 14182 -27593 14242 -27533
rect 14502 -27593 14562 -27533
rect 14640 -27593 14700 -27533
rect 14960 -27593 15020 -27533
rect 15096 -27593 15156 -27533
rect 15416 -27593 15476 -27533
rect 466 -27943 526 -27883
rect 786 -27943 846 -27883
rect 922 -27943 982 -27883
rect 1242 -27943 1302 -27883
rect 1380 -27943 1440 -27883
rect 1700 -27943 1760 -27883
rect 1836 -27943 1896 -27883
rect 2156 -27943 2216 -27883
rect 2292 -27943 2352 -27883
rect 2612 -27943 2672 -27883
rect 2750 -27943 2810 -27883
rect 3070 -27943 3130 -27883
rect 3206 -27943 3266 -27883
rect 3526 -27943 3586 -27883
rect 3662 -27943 3722 -27883
rect 3982 -27943 4042 -27883
rect 4120 -27943 4180 -27883
rect 4440 -27943 4500 -27883
rect 4576 -27943 4636 -27883
rect 4896 -27943 4956 -27883
rect 5032 -27943 5092 -27883
rect 5352 -27943 5412 -27883
rect 5490 -27943 5550 -27883
rect 5810 -27943 5870 -27883
rect 5946 -27943 6006 -27883
rect 6266 -27943 6326 -27883
rect 6402 -27943 6462 -27883
rect 6722 -27943 6782 -27883
rect 6860 -27943 6920 -27883
rect 7180 -27943 7240 -27883
rect 7316 -27943 7376 -27883
rect 7636 -27943 7696 -27883
rect 7772 -27943 7832 -27883
rect 8092 -27943 8152 -27883
rect 8246 -27943 8306 -27883
rect 8566 -27943 8626 -27883
rect 8702 -27943 8762 -27883
rect 9022 -27943 9082 -27883
rect 9160 -27943 9220 -27883
rect 9480 -27943 9540 -27883
rect 9616 -27943 9676 -27883
rect 9936 -27943 9996 -27883
rect 10072 -27943 10132 -27883
rect 10392 -27943 10452 -27883
rect 10530 -27943 10590 -27883
rect 10850 -27943 10910 -27883
rect 10986 -27943 11046 -27883
rect 11306 -27943 11366 -27883
rect 11442 -27943 11502 -27883
rect 11762 -27943 11822 -27883
rect 11900 -27943 11960 -27883
rect 12220 -27943 12280 -27883
rect 12356 -27943 12416 -27883
rect 12676 -27943 12736 -27883
rect 12812 -27943 12872 -27883
rect 13132 -27943 13192 -27883
rect 13270 -27943 13330 -27883
rect 13590 -27943 13650 -27883
rect 13726 -27943 13786 -27883
rect 14046 -27943 14106 -27883
rect 14182 -27943 14242 -27883
rect 14502 -27943 14562 -27883
rect 14640 -27943 14700 -27883
rect 14960 -27943 15020 -27883
rect 15096 -27943 15156 -27883
rect 15416 -27943 15476 -27883
rect 10 -28085 14 -28025
rect 14 -28085 66 -28025
rect 66 -28085 70 -28025
rect 330 -28085 390 -28025
rect 10 -28435 14 -28375
rect 14 -28435 66 -28375
rect 66 -28435 70 -28375
rect 330 -28435 390 -28375
rect 466 -28085 526 -28025
rect 786 -28085 846 -28025
rect 922 -28085 982 -28025
rect 1242 -28085 1302 -28025
rect 1380 -28085 1440 -28025
rect 1700 -28085 1760 -28025
rect 1836 -28085 1896 -28025
rect 2156 -28085 2216 -28025
rect 2292 -28085 2352 -28025
rect 2612 -28085 2672 -28025
rect 2750 -28085 2810 -28025
rect 3070 -28085 3130 -28025
rect 3206 -28085 3266 -28025
rect 3526 -28085 3586 -28025
rect 3662 -28085 3722 -28025
rect 3982 -28085 4042 -28025
rect 4120 -28085 4180 -28025
rect 4440 -28085 4500 -28025
rect 4576 -28085 4636 -28025
rect 4896 -28085 4956 -28025
rect 5032 -28085 5092 -28025
rect 5352 -28085 5412 -28025
rect 5490 -28085 5550 -28025
rect 5810 -28085 5870 -28025
rect 5946 -28085 6006 -28025
rect 6266 -28085 6326 -28025
rect 6402 -28085 6462 -28025
rect 6722 -28085 6782 -28025
rect 6860 -28085 6920 -28025
rect 7180 -28085 7240 -28025
rect 7316 -28085 7376 -28025
rect 7636 -28085 7696 -28025
rect 7772 -28085 7832 -28025
rect 8092 -28085 8152 -28025
rect 8246 -28085 8306 -28025
rect 8566 -28085 8626 -28025
rect 8702 -28085 8762 -28025
rect 9022 -28085 9082 -28025
rect 9160 -28085 9220 -28025
rect 9480 -28085 9540 -28025
rect 9616 -28085 9676 -28025
rect 9936 -28085 9996 -28025
rect 10072 -28085 10132 -28025
rect 10392 -28085 10452 -28025
rect 10530 -28085 10590 -28025
rect 10850 -28085 10910 -28025
rect 10986 -28085 11046 -28025
rect 11306 -28085 11366 -28025
rect 11442 -28085 11502 -28025
rect 11762 -28085 11822 -28025
rect 11900 -28085 11960 -28025
rect 12220 -28085 12280 -28025
rect 12356 -28085 12416 -28025
rect 12676 -28085 12736 -28025
rect 12812 -28085 12872 -28025
rect 13132 -28085 13192 -28025
rect 13270 -28085 13330 -28025
rect 13590 -28085 13650 -28025
rect 13726 -28085 13786 -28025
rect 14046 -28085 14106 -28025
rect 14182 -28085 14242 -28025
rect 14502 -28085 14562 -28025
rect 14640 -28085 14700 -28025
rect 14960 -28085 15020 -28025
rect 15096 -28085 15156 -28025
rect 15416 -28085 15476 -28025
rect 466 -28435 526 -28375
rect 786 -28435 846 -28375
rect 922 -28435 982 -28375
rect 1242 -28435 1302 -28375
rect 1380 -28435 1440 -28375
rect 1700 -28435 1760 -28375
rect 1836 -28435 1896 -28375
rect 2156 -28435 2216 -28375
rect 2292 -28435 2352 -28375
rect 2612 -28435 2672 -28375
rect 2750 -28435 2810 -28375
rect 3070 -28435 3130 -28375
rect 3206 -28435 3266 -28375
rect 3526 -28435 3586 -28375
rect 3662 -28435 3722 -28375
rect 3982 -28435 4042 -28375
rect 4120 -28435 4180 -28375
rect 4440 -28435 4500 -28375
rect 4576 -28435 4636 -28375
rect 4896 -28435 4956 -28375
rect 5032 -28435 5092 -28375
rect 5352 -28435 5412 -28375
rect 5490 -28435 5550 -28375
rect 5810 -28435 5870 -28375
rect 5946 -28435 6006 -28375
rect 6266 -28435 6326 -28375
rect 6402 -28435 6462 -28375
rect 6722 -28435 6782 -28375
rect 6860 -28435 6920 -28375
rect 7180 -28435 7240 -28375
rect 7316 -28435 7376 -28375
rect 7636 -28435 7696 -28375
rect 7772 -28435 7832 -28375
rect 8092 -28435 8152 -28375
rect 8246 -28435 8306 -28375
rect 8566 -28435 8626 -28375
rect 8702 -28435 8762 -28375
rect 9022 -28435 9082 -28375
rect 9160 -28435 9220 -28375
rect 9480 -28435 9540 -28375
rect 9616 -28435 9676 -28375
rect 9936 -28435 9996 -28375
rect 10072 -28435 10132 -28375
rect 10392 -28435 10452 -28375
rect 10530 -28435 10590 -28375
rect 10850 -28435 10910 -28375
rect 10986 -28435 11046 -28375
rect 11306 -28435 11366 -28375
rect 11442 -28435 11502 -28375
rect 11762 -28435 11822 -28375
rect 11900 -28435 11960 -28375
rect 12220 -28435 12280 -28375
rect 12356 -28435 12416 -28375
rect 12676 -28435 12736 -28375
rect 12812 -28435 12872 -28375
rect 13132 -28435 13192 -28375
rect 13270 -28435 13330 -28375
rect 13590 -28435 13650 -28375
rect 13726 -28435 13786 -28375
rect 14046 -28435 14106 -28375
rect 14182 -28435 14242 -28375
rect 14502 -28435 14562 -28375
rect 14640 -28435 14700 -28375
rect 14960 -28435 15020 -28375
rect 15096 -28435 15156 -28375
rect 15416 -28435 15476 -28375
rect 10 -28587 14 -28527
rect 14 -28587 66 -28527
rect 66 -28587 70 -28527
rect 330 -28587 390 -28527
rect 10 -28937 14 -28877
rect 14 -28937 66 -28877
rect 66 -28937 70 -28877
rect 330 -28937 390 -28877
rect 466 -28587 526 -28527
rect 786 -28587 846 -28527
rect 922 -28587 982 -28527
rect 1242 -28587 1302 -28527
rect 1380 -28587 1440 -28527
rect 1700 -28587 1760 -28527
rect 1836 -28587 1896 -28527
rect 2156 -28587 2216 -28527
rect 2292 -28587 2352 -28527
rect 2612 -28587 2672 -28527
rect 2750 -28587 2810 -28527
rect 3070 -28587 3130 -28527
rect 3206 -28587 3266 -28527
rect 3526 -28587 3586 -28527
rect 3662 -28587 3722 -28527
rect 3982 -28587 4042 -28527
rect 4120 -28587 4180 -28527
rect 4440 -28587 4500 -28527
rect 4576 -28587 4636 -28527
rect 4896 -28587 4956 -28527
rect 5032 -28587 5092 -28527
rect 5352 -28587 5412 -28527
rect 5490 -28587 5550 -28527
rect 5810 -28587 5870 -28527
rect 5946 -28587 6006 -28527
rect 6266 -28587 6326 -28527
rect 6402 -28587 6462 -28527
rect 6722 -28587 6782 -28527
rect 6860 -28587 6920 -28527
rect 7180 -28587 7240 -28527
rect 7316 -28587 7376 -28527
rect 7636 -28587 7696 -28527
rect 7772 -28587 7832 -28527
rect 8092 -28587 8152 -28527
rect 8246 -28587 8306 -28527
rect 8566 -28587 8626 -28527
rect 8702 -28587 8762 -28527
rect 9022 -28587 9082 -28527
rect 9160 -28587 9220 -28527
rect 9480 -28587 9540 -28527
rect 9616 -28587 9676 -28527
rect 9936 -28587 9996 -28527
rect 10072 -28587 10132 -28527
rect 10392 -28587 10452 -28527
rect 10530 -28587 10590 -28527
rect 10850 -28587 10910 -28527
rect 10986 -28587 11046 -28527
rect 11306 -28587 11366 -28527
rect 11442 -28587 11502 -28527
rect 11762 -28587 11822 -28527
rect 11900 -28587 11960 -28527
rect 12220 -28587 12280 -28527
rect 12356 -28587 12416 -28527
rect 12676 -28587 12736 -28527
rect 12812 -28587 12872 -28527
rect 13132 -28587 13192 -28527
rect 13270 -28587 13330 -28527
rect 13590 -28587 13650 -28527
rect 13726 -28587 13786 -28527
rect 14046 -28587 14106 -28527
rect 14182 -28587 14242 -28527
rect 14502 -28587 14562 -28527
rect 14640 -28587 14700 -28527
rect 14960 -28587 15020 -28527
rect 15096 -28587 15156 -28527
rect 15416 -28587 15476 -28527
rect 466 -28937 526 -28877
rect 786 -28937 846 -28877
rect 922 -28937 982 -28877
rect 1242 -28937 1302 -28877
rect 1380 -28937 1440 -28877
rect 1700 -28937 1760 -28877
rect 1836 -28937 1896 -28877
rect 2156 -28937 2216 -28877
rect 2292 -28937 2352 -28877
rect 2612 -28937 2672 -28877
rect 2750 -28937 2810 -28877
rect 3070 -28937 3130 -28877
rect 3206 -28937 3266 -28877
rect 3526 -28937 3586 -28877
rect 3662 -28937 3722 -28877
rect 3982 -28937 4042 -28877
rect 4120 -28937 4180 -28877
rect 4440 -28937 4500 -28877
rect 4576 -28937 4636 -28877
rect 4896 -28937 4956 -28877
rect 5032 -28937 5092 -28877
rect 5352 -28937 5412 -28877
rect 5490 -28937 5550 -28877
rect 5810 -28937 5870 -28877
rect 5946 -28937 6006 -28877
rect 6266 -28937 6326 -28877
rect 6402 -28937 6462 -28877
rect 6722 -28937 6782 -28877
rect 6860 -28937 6920 -28877
rect 7180 -28937 7240 -28877
rect 7316 -28937 7376 -28877
rect 7636 -28937 7696 -28877
rect 7772 -28937 7832 -28877
rect 8092 -28937 8152 -28877
rect 8246 -28937 8306 -28877
rect 8566 -28937 8626 -28877
rect 8702 -28937 8762 -28877
rect 9022 -28937 9082 -28877
rect 9160 -28937 9220 -28877
rect 9480 -28937 9540 -28877
rect 9616 -28937 9676 -28877
rect 9936 -28937 9996 -28877
rect 10072 -28937 10132 -28877
rect 10392 -28937 10452 -28877
rect 10530 -28937 10590 -28877
rect 10850 -28937 10910 -28877
rect 10986 -28937 11046 -28877
rect 11306 -28937 11366 -28877
rect 11442 -28937 11502 -28877
rect 11762 -28937 11822 -28877
rect 11900 -28937 11960 -28877
rect 12220 -28937 12280 -28877
rect 12356 -28937 12416 -28877
rect 12676 -28937 12736 -28877
rect 12812 -28937 12872 -28877
rect 13132 -28937 13192 -28877
rect 13270 -28937 13330 -28877
rect 13590 -28937 13650 -28877
rect 13726 -28937 13786 -28877
rect 14046 -28937 14106 -28877
rect 14182 -28937 14242 -28877
rect 14502 -28937 14562 -28877
rect 14640 -28937 14700 -28877
rect 14960 -28937 15020 -28877
rect 15096 -28937 15156 -28877
rect 15416 -28937 15476 -28877
rect 10 -29081 14 -29021
rect 14 -29081 66 -29021
rect 66 -29081 70 -29021
rect 330 -29081 390 -29021
rect 10 -29431 14 -29371
rect 14 -29431 66 -29371
rect 66 -29431 70 -29371
rect 330 -29431 390 -29371
rect 466 -29081 526 -29021
rect 786 -29081 846 -29021
rect 922 -29081 982 -29021
rect 1242 -29081 1302 -29021
rect 1380 -29081 1440 -29021
rect 1700 -29081 1760 -29021
rect 1836 -29081 1896 -29021
rect 2156 -29081 2216 -29021
rect 2292 -29081 2352 -29021
rect 2612 -29081 2672 -29021
rect 2750 -29081 2810 -29021
rect 3070 -29081 3130 -29021
rect 3206 -29081 3266 -29021
rect 3526 -29081 3586 -29021
rect 3662 -29081 3722 -29021
rect 3982 -29081 4042 -29021
rect 4120 -29081 4180 -29021
rect 4440 -29081 4500 -29021
rect 4576 -29081 4636 -29021
rect 4896 -29081 4956 -29021
rect 5032 -29081 5092 -29021
rect 5352 -29081 5412 -29021
rect 5490 -29081 5550 -29021
rect 5810 -29081 5870 -29021
rect 5946 -29081 6006 -29021
rect 6266 -29081 6326 -29021
rect 6402 -29081 6462 -29021
rect 6722 -29081 6782 -29021
rect 6860 -29081 6920 -29021
rect 7180 -29081 7240 -29021
rect 7316 -29081 7376 -29021
rect 7636 -29081 7696 -29021
rect 7772 -29081 7832 -29021
rect 8092 -29081 8152 -29021
rect 8246 -29081 8306 -29021
rect 8566 -29081 8626 -29021
rect 8702 -29081 8762 -29021
rect 9022 -29081 9082 -29021
rect 9160 -29081 9220 -29021
rect 9480 -29081 9540 -29021
rect 9616 -29081 9676 -29021
rect 9936 -29081 9996 -29021
rect 10072 -29081 10132 -29021
rect 10392 -29081 10452 -29021
rect 10530 -29081 10590 -29021
rect 10850 -29081 10910 -29021
rect 10986 -29081 11046 -29021
rect 11306 -29081 11366 -29021
rect 11442 -29081 11502 -29021
rect 11762 -29081 11822 -29021
rect 11900 -29081 11960 -29021
rect 12220 -29081 12280 -29021
rect 12356 -29081 12416 -29021
rect 12676 -29081 12736 -29021
rect 12812 -29081 12872 -29021
rect 13132 -29081 13192 -29021
rect 13270 -29081 13330 -29021
rect 13590 -29081 13650 -29021
rect 13726 -29081 13786 -29021
rect 14046 -29081 14106 -29021
rect 14182 -29081 14242 -29021
rect 14502 -29081 14562 -29021
rect 14640 -29081 14700 -29021
rect 14960 -29081 15020 -29021
rect 15096 -29081 15156 -29021
rect 15416 -29081 15476 -29021
rect 466 -29431 526 -29371
rect 786 -29431 846 -29371
rect 922 -29431 982 -29371
rect 1242 -29431 1302 -29371
rect 1380 -29431 1440 -29371
rect 1700 -29431 1760 -29371
rect 1836 -29431 1896 -29371
rect 2156 -29431 2216 -29371
rect 2292 -29431 2352 -29371
rect 2612 -29431 2672 -29371
rect 2750 -29431 2810 -29371
rect 3070 -29431 3130 -29371
rect 3206 -29431 3266 -29371
rect 3526 -29431 3586 -29371
rect 3662 -29431 3722 -29371
rect 3982 -29431 4042 -29371
rect 4120 -29431 4180 -29371
rect 4440 -29431 4500 -29371
rect 4576 -29431 4636 -29371
rect 4896 -29431 4956 -29371
rect 5032 -29431 5092 -29371
rect 5352 -29431 5412 -29371
rect 5490 -29431 5550 -29371
rect 5810 -29431 5870 -29371
rect 5946 -29431 6006 -29371
rect 6266 -29431 6326 -29371
rect 6402 -29431 6462 -29371
rect 6722 -29431 6782 -29371
rect 6860 -29431 6920 -29371
rect 7180 -29431 7240 -29371
rect 7316 -29431 7376 -29371
rect 7636 -29431 7696 -29371
rect 7772 -29431 7832 -29371
rect 8092 -29431 8152 -29371
rect 8246 -29431 8306 -29371
rect 8566 -29431 8626 -29371
rect 8702 -29431 8762 -29371
rect 9022 -29431 9082 -29371
rect 9160 -29431 9220 -29371
rect 9480 -29431 9540 -29371
rect 9616 -29431 9676 -29371
rect 9936 -29431 9996 -29371
rect 10072 -29431 10132 -29371
rect 10392 -29431 10452 -29371
rect 10530 -29431 10590 -29371
rect 10850 -29431 10910 -29371
rect 10986 -29431 11046 -29371
rect 11306 -29431 11366 -29371
rect 11442 -29431 11502 -29371
rect 11762 -29431 11822 -29371
rect 11900 -29431 11960 -29371
rect 12220 -29431 12280 -29371
rect 12356 -29431 12416 -29371
rect 12676 -29431 12736 -29371
rect 12812 -29431 12872 -29371
rect 13132 -29431 13192 -29371
rect 13270 -29431 13330 -29371
rect 13590 -29431 13650 -29371
rect 13726 -29431 13786 -29371
rect 14046 -29431 14106 -29371
rect 14182 -29431 14242 -29371
rect 14502 -29431 14562 -29371
rect 14640 -29431 14700 -29371
rect 14960 -29431 15020 -29371
rect 15096 -29431 15156 -29371
rect 15416 -29431 15476 -29371
rect 10 -29573 14 -29513
rect 14 -29573 66 -29513
rect 66 -29573 70 -29513
rect 330 -29573 390 -29513
rect 10 -29923 14 -29863
rect 14 -29923 66 -29863
rect 66 -29923 70 -29863
rect 330 -29923 390 -29863
rect 466 -29573 526 -29513
rect 786 -29573 846 -29513
rect 922 -29573 982 -29513
rect 1242 -29573 1302 -29513
rect 1380 -29573 1440 -29513
rect 1700 -29573 1760 -29513
rect 1836 -29573 1896 -29513
rect 2156 -29573 2216 -29513
rect 2292 -29573 2352 -29513
rect 2612 -29573 2672 -29513
rect 2750 -29573 2810 -29513
rect 3070 -29573 3130 -29513
rect 3206 -29573 3266 -29513
rect 3526 -29573 3586 -29513
rect 3662 -29573 3722 -29513
rect 3982 -29573 4042 -29513
rect 4120 -29573 4180 -29513
rect 4440 -29573 4500 -29513
rect 4576 -29573 4636 -29513
rect 4896 -29573 4956 -29513
rect 5032 -29573 5092 -29513
rect 5352 -29573 5412 -29513
rect 5490 -29573 5550 -29513
rect 5810 -29573 5870 -29513
rect 5946 -29573 6006 -29513
rect 6266 -29573 6326 -29513
rect 6402 -29573 6462 -29513
rect 6722 -29573 6782 -29513
rect 6860 -29573 6920 -29513
rect 7180 -29573 7240 -29513
rect 7316 -29573 7376 -29513
rect 7636 -29573 7696 -29513
rect 7772 -29573 7832 -29513
rect 8092 -29573 8152 -29513
rect 8246 -29573 8306 -29513
rect 8566 -29573 8626 -29513
rect 8702 -29573 8762 -29513
rect 9022 -29573 9082 -29513
rect 9160 -29573 9220 -29513
rect 9480 -29573 9540 -29513
rect 9616 -29573 9676 -29513
rect 9936 -29573 9996 -29513
rect 10072 -29573 10132 -29513
rect 10392 -29573 10452 -29513
rect 10530 -29573 10590 -29513
rect 10850 -29573 10910 -29513
rect 10986 -29573 11046 -29513
rect 11306 -29573 11366 -29513
rect 11442 -29573 11502 -29513
rect 11762 -29573 11822 -29513
rect 11900 -29573 11960 -29513
rect 12220 -29573 12280 -29513
rect 12356 -29573 12416 -29513
rect 12676 -29573 12736 -29513
rect 12812 -29573 12872 -29513
rect 13132 -29573 13192 -29513
rect 13270 -29573 13330 -29513
rect 13590 -29573 13650 -29513
rect 13726 -29573 13786 -29513
rect 14046 -29573 14106 -29513
rect 14182 -29573 14242 -29513
rect 14502 -29573 14562 -29513
rect 14640 -29573 14700 -29513
rect 14960 -29573 15020 -29513
rect 15096 -29573 15156 -29513
rect 15416 -29573 15476 -29513
rect 466 -29923 526 -29863
rect 786 -29923 846 -29863
rect 922 -29923 982 -29863
rect 1242 -29923 1302 -29863
rect 1380 -29923 1440 -29863
rect 1700 -29923 1760 -29863
rect 1836 -29923 1896 -29863
rect 2156 -29923 2216 -29863
rect 2292 -29923 2352 -29863
rect 2612 -29923 2672 -29863
rect 2750 -29923 2810 -29863
rect 3070 -29923 3130 -29863
rect 3206 -29923 3266 -29863
rect 3526 -29923 3586 -29863
rect 3662 -29923 3722 -29863
rect 3982 -29923 4042 -29863
rect 4120 -29923 4180 -29863
rect 4440 -29923 4500 -29863
rect 4576 -29923 4636 -29863
rect 4896 -29923 4956 -29863
rect 5032 -29923 5092 -29863
rect 5352 -29923 5412 -29863
rect 5490 -29923 5550 -29863
rect 5810 -29923 5870 -29863
rect 5946 -29923 6006 -29863
rect 6266 -29923 6326 -29863
rect 6402 -29923 6462 -29863
rect 6722 -29923 6782 -29863
rect 6860 -29923 6920 -29863
rect 7180 -29923 7240 -29863
rect 7316 -29923 7376 -29863
rect 7636 -29923 7696 -29863
rect 7772 -29923 7832 -29863
rect 8092 -29923 8152 -29863
rect 8246 -29923 8306 -29863
rect 8566 -29923 8626 -29863
rect 8702 -29923 8762 -29863
rect 9022 -29923 9082 -29863
rect 9160 -29923 9220 -29863
rect 9480 -29923 9540 -29863
rect 9616 -29923 9676 -29863
rect 9936 -29923 9996 -29863
rect 10072 -29923 10132 -29863
rect 10392 -29923 10452 -29863
rect 10530 -29923 10590 -29863
rect 10850 -29923 10910 -29863
rect 10986 -29923 11046 -29863
rect 11306 -29923 11366 -29863
rect 11442 -29923 11502 -29863
rect 11762 -29923 11822 -29863
rect 11900 -29923 11960 -29863
rect 12220 -29923 12280 -29863
rect 12356 -29923 12416 -29863
rect 12676 -29923 12736 -29863
rect 12812 -29923 12872 -29863
rect 13132 -29923 13192 -29863
rect 13270 -29923 13330 -29863
rect 13590 -29923 13650 -29863
rect 13726 -29923 13786 -29863
rect 14046 -29923 14106 -29863
rect 14182 -29923 14242 -29863
rect 14502 -29923 14562 -29863
rect 14640 -29923 14700 -29863
rect 14960 -29923 15020 -29863
rect 15096 -29923 15156 -29863
rect 15416 -29923 15476 -29863
rect 10 -30075 14 -30015
rect 14 -30075 66 -30015
rect 66 -30075 70 -30015
rect 330 -30075 390 -30015
rect 10 -30425 14 -30365
rect 14 -30425 66 -30365
rect 66 -30425 70 -30365
rect 330 -30425 390 -30365
rect 466 -30075 526 -30015
rect 786 -30075 846 -30015
rect 922 -30075 982 -30015
rect 1242 -30075 1302 -30015
rect 1380 -30075 1440 -30015
rect 1700 -30075 1760 -30015
rect 1836 -30075 1896 -30015
rect 2156 -30075 2216 -30015
rect 2292 -30075 2352 -30015
rect 2612 -30075 2672 -30015
rect 2750 -30075 2810 -30015
rect 3070 -30075 3130 -30015
rect 3206 -30075 3266 -30015
rect 3526 -30075 3586 -30015
rect 3662 -30075 3722 -30015
rect 3982 -30075 4042 -30015
rect 4120 -30075 4180 -30015
rect 4440 -30075 4500 -30015
rect 4576 -30075 4636 -30015
rect 4896 -30075 4956 -30015
rect 5032 -30075 5092 -30015
rect 5352 -30075 5412 -30015
rect 5490 -30075 5550 -30015
rect 5810 -30075 5870 -30015
rect 5946 -30075 6006 -30015
rect 6266 -30075 6326 -30015
rect 6402 -30075 6462 -30015
rect 6722 -30075 6782 -30015
rect 6860 -30075 6920 -30015
rect 7180 -30075 7240 -30015
rect 7316 -30075 7376 -30015
rect 7636 -30075 7696 -30015
rect 7772 -30075 7832 -30015
rect 8092 -30075 8152 -30015
rect 8246 -30075 8306 -30015
rect 8566 -30075 8626 -30015
rect 8702 -30075 8762 -30015
rect 9022 -30075 9082 -30015
rect 9160 -30075 9220 -30015
rect 9480 -30075 9540 -30015
rect 9616 -30075 9676 -30015
rect 9936 -30075 9996 -30015
rect 10072 -30075 10132 -30015
rect 10392 -30075 10452 -30015
rect 10530 -30075 10590 -30015
rect 10850 -30075 10910 -30015
rect 10986 -30075 11046 -30015
rect 11306 -30075 11366 -30015
rect 11442 -30075 11502 -30015
rect 11762 -30075 11822 -30015
rect 11900 -30075 11960 -30015
rect 12220 -30075 12280 -30015
rect 12356 -30075 12416 -30015
rect 12676 -30075 12736 -30015
rect 12812 -30075 12872 -30015
rect 13132 -30075 13192 -30015
rect 13270 -30075 13330 -30015
rect 13590 -30075 13650 -30015
rect 13726 -30075 13786 -30015
rect 14046 -30075 14106 -30015
rect 14182 -30075 14242 -30015
rect 14502 -30075 14562 -30015
rect 14640 -30075 14700 -30015
rect 14960 -30075 15020 -30015
rect 15096 -30075 15156 -30015
rect 15416 -30075 15476 -30015
rect 466 -30425 526 -30365
rect 786 -30425 846 -30365
rect 922 -30425 982 -30365
rect 1242 -30425 1302 -30365
rect 1380 -30425 1440 -30365
rect 1700 -30425 1760 -30365
rect 1836 -30425 1896 -30365
rect 2156 -30425 2216 -30365
rect 2292 -30425 2352 -30365
rect 2612 -30425 2672 -30365
rect 2750 -30425 2810 -30365
rect 3070 -30425 3130 -30365
rect 3206 -30425 3266 -30365
rect 3526 -30425 3586 -30365
rect 3662 -30425 3722 -30365
rect 3982 -30425 4042 -30365
rect 4120 -30425 4180 -30365
rect 4440 -30425 4500 -30365
rect 4576 -30425 4636 -30365
rect 4896 -30425 4956 -30365
rect 5032 -30425 5092 -30365
rect 5352 -30425 5412 -30365
rect 5490 -30425 5550 -30365
rect 5810 -30425 5870 -30365
rect 5946 -30425 6006 -30365
rect 6266 -30425 6326 -30365
rect 6402 -30425 6462 -30365
rect 6722 -30425 6782 -30365
rect 6860 -30425 6920 -30365
rect 7180 -30425 7240 -30365
rect 7316 -30425 7376 -30365
rect 7636 -30425 7696 -30365
rect 7772 -30425 7832 -30365
rect 8092 -30425 8152 -30365
rect 8246 -30425 8306 -30365
rect 8566 -30425 8626 -30365
rect 8702 -30425 8762 -30365
rect 9022 -30425 9082 -30365
rect 9160 -30425 9220 -30365
rect 9480 -30425 9540 -30365
rect 9616 -30425 9676 -30365
rect 9936 -30425 9996 -30365
rect 10072 -30425 10132 -30365
rect 10392 -30425 10452 -30365
rect 10530 -30425 10590 -30365
rect 10850 -30425 10910 -30365
rect 10986 -30425 11046 -30365
rect 11306 -30425 11366 -30365
rect 11442 -30425 11502 -30365
rect 11762 -30425 11822 -30365
rect 11900 -30425 11960 -30365
rect 12220 -30425 12280 -30365
rect 12356 -30425 12416 -30365
rect 12676 -30425 12736 -30365
rect 12812 -30425 12872 -30365
rect 13132 -30425 13192 -30365
rect 13270 -30425 13330 -30365
rect 13590 -30425 13650 -30365
rect 13726 -30425 13786 -30365
rect 14046 -30425 14106 -30365
rect 14182 -30425 14242 -30365
rect 14502 -30425 14562 -30365
rect 14640 -30425 14700 -30365
rect 14960 -30425 15020 -30365
rect 15096 -30425 15156 -30365
rect 15416 -30425 15476 -30365
rect 10 -30591 14 -30531
rect 14 -30591 66 -30531
rect 66 -30591 70 -30531
rect 330 -30591 390 -30531
rect 10 -30941 14 -30881
rect 14 -30941 66 -30881
rect 66 -30941 70 -30881
rect 330 -30941 390 -30881
rect 466 -30591 526 -30531
rect 786 -30591 846 -30531
rect 922 -30591 982 -30531
rect 1242 -30591 1302 -30531
rect 1380 -30591 1440 -30531
rect 1700 -30591 1760 -30531
rect 1836 -30591 1896 -30531
rect 2156 -30591 2216 -30531
rect 2292 -30591 2352 -30531
rect 2612 -30591 2672 -30531
rect 2750 -30591 2810 -30531
rect 3070 -30591 3130 -30531
rect 3206 -30591 3266 -30531
rect 3526 -30591 3586 -30531
rect 3662 -30591 3722 -30531
rect 3982 -30591 4042 -30531
rect 4120 -30591 4180 -30531
rect 4440 -30591 4500 -30531
rect 4576 -30591 4636 -30531
rect 4896 -30591 4956 -30531
rect 5032 -30591 5092 -30531
rect 5352 -30591 5412 -30531
rect 5490 -30591 5550 -30531
rect 5810 -30591 5870 -30531
rect 5946 -30591 6006 -30531
rect 6266 -30591 6326 -30531
rect 6402 -30591 6462 -30531
rect 6722 -30591 6782 -30531
rect 6860 -30591 6920 -30531
rect 7180 -30591 7240 -30531
rect 7316 -30591 7376 -30531
rect 7636 -30591 7696 -30531
rect 7772 -30591 7832 -30531
rect 8092 -30591 8152 -30531
rect 8246 -30591 8306 -30531
rect 8566 -30591 8626 -30531
rect 8702 -30591 8762 -30531
rect 9022 -30591 9082 -30531
rect 9160 -30591 9220 -30531
rect 9480 -30591 9540 -30531
rect 9616 -30591 9676 -30531
rect 9936 -30591 9996 -30531
rect 10072 -30591 10132 -30531
rect 10392 -30591 10452 -30531
rect 10530 -30591 10590 -30531
rect 10850 -30591 10910 -30531
rect 10986 -30591 11046 -30531
rect 11306 -30591 11366 -30531
rect 11442 -30591 11502 -30531
rect 11762 -30591 11822 -30531
rect 11900 -30591 11960 -30531
rect 12220 -30591 12280 -30531
rect 12356 -30591 12416 -30531
rect 12676 -30591 12736 -30531
rect 12812 -30591 12872 -30531
rect 13132 -30591 13192 -30531
rect 13270 -30591 13330 -30531
rect 13590 -30591 13650 -30531
rect 13726 -30591 13786 -30531
rect 14046 -30591 14106 -30531
rect 14182 -30591 14242 -30531
rect 14502 -30591 14562 -30531
rect 14640 -30591 14700 -30531
rect 14960 -30591 15020 -30531
rect 15096 -30591 15156 -30531
rect 15416 -30591 15476 -30531
rect 466 -30941 526 -30881
rect 786 -30941 846 -30881
rect 922 -30941 982 -30881
rect 1242 -30941 1302 -30881
rect 1380 -30941 1440 -30881
rect 1700 -30941 1760 -30881
rect 1836 -30941 1896 -30881
rect 2156 -30941 2216 -30881
rect 2292 -30941 2352 -30881
rect 2612 -30941 2672 -30881
rect 2750 -30941 2810 -30881
rect 3070 -30941 3130 -30881
rect 3206 -30941 3266 -30881
rect 3526 -30941 3586 -30881
rect 3662 -30941 3722 -30881
rect 3982 -30941 4042 -30881
rect 4120 -30941 4180 -30881
rect 4440 -30941 4500 -30881
rect 4576 -30941 4636 -30881
rect 4896 -30941 4956 -30881
rect 5032 -30941 5092 -30881
rect 5352 -30941 5412 -30881
rect 5490 -30941 5550 -30881
rect 5810 -30941 5870 -30881
rect 5946 -30941 6006 -30881
rect 6266 -30941 6326 -30881
rect 6402 -30941 6462 -30881
rect 6722 -30941 6782 -30881
rect 6860 -30941 6920 -30881
rect 7180 -30941 7240 -30881
rect 7316 -30941 7376 -30881
rect 7636 -30941 7696 -30881
rect 7772 -30941 7832 -30881
rect 8092 -30941 8152 -30881
rect 8246 -30941 8306 -30881
rect 8566 -30941 8626 -30881
rect 8702 -30941 8762 -30881
rect 9022 -30941 9082 -30881
rect 9160 -30941 9220 -30881
rect 9480 -30941 9540 -30881
rect 9616 -30941 9676 -30881
rect 9936 -30941 9996 -30881
rect 10072 -30941 10132 -30881
rect 10392 -30941 10452 -30881
rect 10530 -30941 10590 -30881
rect 10850 -30941 10910 -30881
rect 10986 -30941 11046 -30881
rect 11306 -30941 11366 -30881
rect 11442 -30941 11502 -30881
rect 11762 -30941 11822 -30881
rect 11900 -30941 11960 -30881
rect 12220 -30941 12280 -30881
rect 12356 -30941 12416 -30881
rect 12676 -30941 12736 -30881
rect 12812 -30941 12872 -30881
rect 13132 -30941 13192 -30881
rect 13270 -30941 13330 -30881
rect 13590 -30941 13650 -30881
rect 13726 -30941 13786 -30881
rect 14046 -30941 14106 -30881
rect 14182 -30941 14242 -30881
rect 14502 -30941 14562 -30881
rect 14640 -30941 14700 -30881
rect 14960 -30941 15020 -30881
rect 15096 -30941 15156 -30881
rect 15416 -30941 15476 -30881
rect 10 -31083 14 -31023
rect 14 -31083 66 -31023
rect 66 -31083 70 -31023
rect 330 -31083 390 -31023
rect 10 -31433 14 -31373
rect 14 -31433 66 -31373
rect 66 -31433 70 -31373
rect 330 -31433 390 -31373
rect 466 -31083 526 -31023
rect 786 -31083 846 -31023
rect 922 -31083 982 -31023
rect 1242 -31083 1302 -31023
rect 1380 -31083 1440 -31023
rect 1700 -31083 1760 -31023
rect 1836 -31083 1896 -31023
rect 2156 -31083 2216 -31023
rect 2292 -31083 2352 -31023
rect 2612 -31083 2672 -31023
rect 2750 -31083 2810 -31023
rect 3070 -31083 3130 -31023
rect 3206 -31083 3266 -31023
rect 3526 -31083 3586 -31023
rect 3662 -31083 3722 -31023
rect 3982 -31083 4042 -31023
rect 4120 -31083 4180 -31023
rect 4440 -31083 4500 -31023
rect 4576 -31083 4636 -31023
rect 4896 -31083 4956 -31023
rect 5032 -31083 5092 -31023
rect 5352 -31083 5412 -31023
rect 5490 -31083 5550 -31023
rect 5810 -31083 5870 -31023
rect 5946 -31083 6006 -31023
rect 6266 -31083 6326 -31023
rect 6402 -31083 6462 -31023
rect 6722 -31083 6782 -31023
rect 6860 -31083 6920 -31023
rect 7180 -31083 7240 -31023
rect 7316 -31083 7376 -31023
rect 7636 -31083 7696 -31023
rect 7772 -31083 7832 -31023
rect 8092 -31083 8152 -31023
rect 8246 -31083 8306 -31023
rect 8566 -31083 8626 -31023
rect 8702 -31083 8762 -31023
rect 9022 -31083 9082 -31023
rect 9160 -31083 9220 -31023
rect 9480 -31083 9540 -31023
rect 9616 -31083 9676 -31023
rect 9936 -31083 9996 -31023
rect 10072 -31083 10132 -31023
rect 10392 -31083 10452 -31023
rect 10530 -31083 10590 -31023
rect 10850 -31083 10910 -31023
rect 10986 -31083 11046 -31023
rect 11306 -31083 11366 -31023
rect 11442 -31083 11502 -31023
rect 11762 -31083 11822 -31023
rect 11900 -31083 11960 -31023
rect 12220 -31083 12280 -31023
rect 12356 -31083 12416 -31023
rect 12676 -31083 12736 -31023
rect 12812 -31083 12872 -31023
rect 13132 -31083 13192 -31023
rect 13270 -31083 13330 -31023
rect 13590 -31083 13650 -31023
rect 13726 -31083 13786 -31023
rect 14046 -31083 14106 -31023
rect 14182 -31083 14242 -31023
rect 14502 -31083 14562 -31023
rect 14640 -31083 14700 -31023
rect 14960 -31083 15020 -31023
rect 15096 -31083 15156 -31023
rect 15416 -31083 15476 -31023
rect 466 -31433 526 -31373
rect 786 -31433 846 -31373
rect 922 -31433 982 -31373
rect 1242 -31433 1302 -31373
rect 1380 -31433 1440 -31373
rect 1700 -31433 1760 -31373
rect 1836 -31433 1896 -31373
rect 2156 -31433 2216 -31373
rect 2292 -31433 2352 -31373
rect 2612 -31433 2672 -31373
rect 2750 -31433 2810 -31373
rect 3070 -31433 3130 -31373
rect 3206 -31433 3266 -31373
rect 3526 -31433 3586 -31373
rect 3662 -31433 3722 -31373
rect 3982 -31433 4042 -31373
rect 4120 -31433 4180 -31373
rect 4440 -31433 4500 -31373
rect 4576 -31433 4636 -31373
rect 4896 -31433 4956 -31373
rect 5032 -31433 5092 -31373
rect 5352 -31433 5412 -31373
rect 5490 -31433 5550 -31373
rect 5810 -31433 5870 -31373
rect 5946 -31433 6006 -31373
rect 6266 -31433 6326 -31373
rect 6402 -31433 6462 -31373
rect 6722 -31433 6782 -31373
rect 6860 -31433 6920 -31373
rect 7180 -31433 7240 -31373
rect 7316 -31433 7376 -31373
rect 7636 -31433 7696 -31373
rect 7772 -31433 7832 -31373
rect 8092 -31433 8152 -31373
rect 8246 -31433 8306 -31373
rect 8566 -31433 8626 -31373
rect 8702 -31433 8762 -31373
rect 9022 -31433 9082 -31373
rect 9160 -31433 9220 -31373
rect 9480 -31433 9540 -31373
rect 9616 -31433 9676 -31373
rect 9936 -31433 9996 -31373
rect 10072 -31433 10132 -31373
rect 10392 -31433 10452 -31373
rect 10530 -31433 10590 -31373
rect 10850 -31433 10910 -31373
rect 10986 -31433 11046 -31373
rect 11306 -31433 11366 -31373
rect 11442 -31433 11502 -31373
rect 11762 -31433 11822 -31373
rect 11900 -31433 11960 -31373
rect 12220 -31433 12280 -31373
rect 12356 -31433 12416 -31373
rect 12676 -31433 12736 -31373
rect 12812 -31433 12872 -31373
rect 13132 -31433 13192 -31373
rect 13270 -31433 13330 -31373
rect 13590 -31433 13650 -31373
rect 13726 -31433 13786 -31373
rect 14046 -31433 14106 -31373
rect 14182 -31433 14242 -31373
rect 14502 -31433 14562 -31373
rect 14640 -31433 14700 -31373
rect 14960 -31433 15020 -31373
rect 15096 -31433 15156 -31373
rect 15416 -31433 15476 -31373
rect 10 -31585 14 -31525
rect 14 -31585 66 -31525
rect 66 -31585 70 -31525
rect 330 -31585 390 -31525
rect 10 -31935 14 -31875
rect 14 -31935 66 -31875
rect 66 -31935 70 -31875
rect 330 -31935 390 -31875
rect 466 -31585 526 -31525
rect 786 -31585 846 -31525
rect 922 -31585 982 -31525
rect 1242 -31585 1302 -31525
rect 1380 -31585 1440 -31525
rect 1700 -31585 1760 -31525
rect 1836 -31585 1896 -31525
rect 2156 -31585 2216 -31525
rect 2292 -31585 2352 -31525
rect 2612 -31585 2672 -31525
rect 2750 -31585 2810 -31525
rect 3070 -31585 3130 -31525
rect 3206 -31585 3266 -31525
rect 3526 -31585 3586 -31525
rect 3662 -31585 3722 -31525
rect 3982 -31585 4042 -31525
rect 4120 -31585 4180 -31525
rect 4440 -31585 4500 -31525
rect 4576 -31585 4636 -31525
rect 4896 -31585 4956 -31525
rect 5032 -31585 5092 -31525
rect 5352 -31585 5412 -31525
rect 5490 -31585 5550 -31525
rect 5810 -31585 5870 -31525
rect 5946 -31585 6006 -31525
rect 6266 -31585 6326 -31525
rect 6402 -31585 6462 -31525
rect 6722 -31585 6782 -31525
rect 6860 -31585 6920 -31525
rect 7180 -31585 7240 -31525
rect 7316 -31585 7376 -31525
rect 7636 -31585 7696 -31525
rect 7772 -31585 7832 -31525
rect 8092 -31585 8152 -31525
rect 8246 -31585 8306 -31525
rect 8566 -31585 8626 -31525
rect 8702 -31585 8762 -31525
rect 9022 -31585 9082 -31525
rect 9160 -31585 9220 -31525
rect 9480 -31585 9540 -31525
rect 9616 -31585 9676 -31525
rect 9936 -31585 9996 -31525
rect 10072 -31585 10132 -31525
rect 10392 -31585 10452 -31525
rect 10530 -31585 10590 -31525
rect 10850 -31585 10910 -31525
rect 10986 -31585 11046 -31525
rect 11306 -31585 11366 -31525
rect 11442 -31585 11502 -31525
rect 11762 -31585 11822 -31525
rect 11900 -31585 11960 -31525
rect 12220 -31585 12280 -31525
rect 12356 -31585 12416 -31525
rect 12676 -31585 12736 -31525
rect 12812 -31585 12872 -31525
rect 13132 -31585 13192 -31525
rect 13270 -31585 13330 -31525
rect 13590 -31585 13650 -31525
rect 13726 -31585 13786 -31525
rect 14046 -31585 14106 -31525
rect 14182 -31585 14242 -31525
rect 14502 -31585 14562 -31525
rect 14640 -31585 14700 -31525
rect 14960 -31585 15020 -31525
rect 15096 -31585 15156 -31525
rect 15416 -31585 15476 -31525
rect 466 -31935 526 -31875
rect 786 -31935 846 -31875
rect 922 -31935 982 -31875
rect 1242 -31935 1302 -31875
rect 1380 -31935 1440 -31875
rect 1700 -31935 1760 -31875
rect 1836 -31935 1896 -31875
rect 2156 -31935 2216 -31875
rect 2292 -31935 2352 -31875
rect 2612 -31935 2672 -31875
rect 2750 -31935 2810 -31875
rect 3070 -31935 3130 -31875
rect 3206 -31935 3266 -31875
rect 3526 -31935 3586 -31875
rect 3662 -31935 3722 -31875
rect 3982 -31935 4042 -31875
rect 4120 -31935 4180 -31875
rect 4440 -31935 4500 -31875
rect 4576 -31935 4636 -31875
rect 4896 -31935 4956 -31875
rect 5032 -31935 5092 -31875
rect 5352 -31935 5412 -31875
rect 5490 -31935 5550 -31875
rect 5810 -31935 5870 -31875
rect 5946 -31935 6006 -31875
rect 6266 -31935 6326 -31875
rect 6402 -31935 6462 -31875
rect 6722 -31935 6782 -31875
rect 6860 -31935 6920 -31875
rect 7180 -31935 7240 -31875
rect 7316 -31935 7376 -31875
rect 7636 -31935 7696 -31875
rect 7772 -31935 7832 -31875
rect 8092 -31935 8152 -31875
rect 8246 -31935 8306 -31875
rect 8566 -31935 8626 -31875
rect 8702 -31935 8762 -31875
rect 9022 -31935 9082 -31875
rect 9160 -31935 9220 -31875
rect 9480 -31935 9540 -31875
rect 9616 -31935 9676 -31875
rect 9936 -31935 9996 -31875
rect 10072 -31935 10132 -31875
rect 10392 -31935 10452 -31875
rect 10530 -31935 10590 -31875
rect 10850 -31935 10910 -31875
rect 10986 -31935 11046 -31875
rect 11306 -31935 11366 -31875
rect 11442 -31935 11502 -31875
rect 11762 -31935 11822 -31875
rect 11900 -31935 11960 -31875
rect 12220 -31935 12280 -31875
rect 12356 -31935 12416 -31875
rect 12676 -31935 12736 -31875
rect 12812 -31935 12872 -31875
rect 13132 -31935 13192 -31875
rect 13270 -31935 13330 -31875
rect 13590 -31935 13650 -31875
rect 13726 -31935 13786 -31875
rect 14046 -31935 14106 -31875
rect 14182 -31935 14242 -31875
rect 14502 -31935 14562 -31875
rect 14640 -31935 14700 -31875
rect 14960 -31935 15020 -31875
rect 15096 -31935 15156 -31875
rect 15416 -31935 15476 -31875
rect 10 -32077 14 -32017
rect 14 -32077 66 -32017
rect 66 -32077 70 -32017
rect 330 -32077 390 -32017
rect 466 -32077 526 -32017
rect 786 -32077 846 -32017
rect 922 -32077 982 -32017
rect 1242 -32077 1302 -32017
rect 1380 -32077 1440 -32017
rect 1700 -32077 1760 -32017
rect 1836 -32077 1896 -32017
rect 2156 -32077 2216 -32017
rect 2292 -32077 2352 -32017
rect 2612 -32077 2672 -32017
rect 2750 -32077 2810 -32017
rect 3070 -32077 3130 -32017
rect 3206 -32077 3266 -32017
rect 3526 -32077 3586 -32017
rect 3662 -32077 3722 -32017
rect 3982 -32077 4042 -32017
rect 4120 -32077 4180 -32017
rect 4440 -32077 4500 -32017
rect 4576 -32077 4636 -32017
rect 4896 -32077 4956 -32017
rect 5032 -32077 5092 -32017
rect 5352 -32077 5412 -32017
rect 5490 -32077 5550 -32017
rect 5810 -32077 5870 -32017
rect 5946 -32077 6006 -32017
rect 6266 -32077 6326 -32017
rect 6402 -32077 6462 -32017
rect 6722 -32077 6782 -32017
rect 6860 -32077 6920 -32017
rect 7180 -32077 7240 -32017
rect 7316 -32077 7376 -32017
rect 7636 -32077 7696 -32017
rect 7772 -32077 7832 -32017
rect 8092 -32077 8152 -32017
rect 8246 -32077 8306 -32017
rect 8566 -32077 8626 -32017
rect 8702 -32077 8762 -32017
rect 9022 -32077 9082 -32017
rect 9160 -32077 9220 -32017
rect 9480 -32077 9540 -32017
rect 9616 -32077 9676 -32017
rect 9936 -32077 9996 -32017
rect 10072 -32077 10132 -32017
rect 10392 -32077 10452 -32017
rect 10530 -32077 10590 -32017
rect 10850 -32077 10910 -32017
rect 10986 -32077 11046 -32017
rect 11306 -32077 11366 -32017
rect 11442 -32077 11502 -32017
rect 11762 -32077 11822 -32017
rect 11900 -32077 11960 -32017
rect 12220 -32077 12280 -32017
rect 12356 -32077 12416 -32017
rect 12676 -32077 12736 -32017
rect 12812 -32077 12872 -32017
rect 13132 -32077 13192 -32017
rect 13270 -32077 13330 -32017
rect 13590 -32077 13650 -32017
rect 13726 -32077 13786 -32017
rect 14046 -32077 14106 -32017
rect 14182 -32077 14242 -32017
rect 14502 -32077 14562 -32017
rect 14640 -32077 14700 -32017
rect 14960 -32077 15020 -32017
rect 15096 -32077 15156 -32017
rect 15416 -32077 15476 -32017
rect 10 -32427 70 -32367
rect 330 -32427 390 -32367
rect 466 -32427 526 -32367
rect 786 -32427 846 -32367
rect 922 -32427 982 -32367
rect 1242 -32427 1302 -32367
rect 1380 -32427 1440 -32367
rect 1700 -32427 1760 -32367
rect 1836 -32427 1896 -32367
rect 2156 -32427 2216 -32367
rect 2292 -32427 2352 -32367
rect 2612 -32427 2672 -32367
rect 2750 -32427 2810 -32367
rect 3070 -32427 3130 -32367
rect 3206 -32427 3266 -32367
rect 3526 -32427 3586 -32367
rect 3662 -32427 3722 -32367
rect 3982 -32427 4042 -32367
rect 4120 -32427 4180 -32367
rect 4440 -32427 4500 -32367
rect 4576 -32427 4636 -32367
rect 4896 -32427 4956 -32367
rect 5032 -32427 5092 -32367
rect 5352 -32427 5412 -32367
rect 5490 -32427 5550 -32367
rect 5810 -32427 5870 -32367
rect 5946 -32427 6006 -32367
rect 6266 -32427 6326 -32367
rect 6402 -32427 6462 -32367
rect 6722 -32427 6782 -32367
rect 6860 -32427 6920 -32367
rect 7180 -32427 7240 -32367
rect 7316 -32427 7376 -32367
rect 7636 -32427 7696 -32367
rect 7772 -32427 7832 -32367
rect 8092 -32427 8152 -32367
rect 8246 -32427 8306 -32367
rect 8566 -32427 8626 -32367
rect 8702 -32427 8762 -32367
rect 9022 -32427 9082 -32367
rect 9160 -32427 9220 -32367
rect 9480 -32427 9540 -32367
rect 9616 -32427 9676 -32367
rect 9936 -32427 9996 -32367
rect 10072 -32427 10132 -32367
rect 10392 -32427 10452 -32367
rect 10530 -32427 10590 -32367
rect 10850 -32427 10910 -32367
rect 10986 -32427 11046 -32367
rect 11306 -32427 11366 -32367
rect 11442 -32427 11502 -32367
rect 11762 -32427 11822 -32367
rect 11900 -32427 11960 -32367
rect 12220 -32427 12280 -32367
rect 12356 -32427 12416 -32367
rect 12676 -32427 12736 -32367
rect 12812 -32427 12872 -32367
rect 13132 -32427 13192 -32367
rect 13270 -32427 13330 -32367
rect 13590 -32427 13650 -32367
rect 13726 -32427 13786 -32367
rect 14046 -32427 14106 -32367
rect 14182 -32427 14242 -32367
rect 14502 -32427 14562 -32367
rect 14640 -32427 14700 -32367
rect 14960 -32427 15020 -32367
rect 15096 -32427 15156 -32367
rect 15416 -32427 15476 -32367
<< metal3 >>
rect 78 651 321 661
rect 78 590 89 651
rect 150 590 250 651
rect 311 590 321 651
rect 78 580 321 590
rect 15111 611 15452 623
rect 15111 551 15127 611
rect 15201 551 15358 611
rect 15432 551 15452 611
rect 15111 539 15452 551
rect 1370 440 1770 450
rect 1370 380 1380 440
rect 1440 390 1700 440
rect 1440 380 1450 390
rect 1370 370 1450 380
rect 1690 380 1700 390
rect 1760 380 1770 440
rect 1690 370 1770 380
rect 1370 100 1430 370
rect 1700 360 1770 370
rect 1510 310 1540 330
rect 1490 270 1540 310
rect 1600 310 1630 330
rect 1600 270 1650 310
rect 1490 200 1650 270
rect 1490 160 1540 200
rect 1510 140 1540 160
rect 1600 160 1650 200
rect 1600 140 1630 160
rect 1710 100 1770 360
rect 1370 90 1450 100
rect 1370 30 1380 90
rect 1440 80 1450 90
rect 1690 90 1770 100
rect 1690 80 1700 90
rect 1440 30 1700 80
rect 1760 30 1770 90
rect 1370 20 1770 30
rect 1826 440 2226 450
rect 1826 380 1836 440
rect 1896 390 2156 440
rect 1896 380 1906 390
rect 1826 370 1906 380
rect 2146 380 2156 390
rect 2216 380 2226 440
rect 2146 370 2226 380
rect 1826 100 1886 370
rect 2156 360 2226 370
rect 1966 310 1996 330
rect 1946 270 1996 310
rect 2056 310 2086 330
rect 2056 270 2106 310
rect 1946 200 2106 270
rect 1946 160 1996 200
rect 1966 140 1996 160
rect 2056 160 2106 200
rect 2056 140 2086 160
rect 2166 100 2226 360
rect 1826 90 1906 100
rect 1826 30 1836 90
rect 1896 80 1906 90
rect 2146 90 2226 100
rect 2146 80 2156 90
rect 1896 30 2156 80
rect 2216 30 2226 90
rect 1826 20 2226 30
rect 2282 440 2682 450
rect 2282 380 2292 440
rect 2352 390 2612 440
rect 2352 380 2362 390
rect 2282 370 2362 380
rect 2602 380 2612 390
rect 2672 380 2682 440
rect 2602 370 2682 380
rect 2282 100 2342 370
rect 2612 360 2682 370
rect 2422 310 2452 330
rect 2402 270 2452 310
rect 2512 310 2542 330
rect 2512 270 2562 310
rect 2402 200 2562 270
rect 2402 160 2452 200
rect 2422 140 2452 160
rect 2512 160 2562 200
rect 2512 140 2542 160
rect 2622 100 2682 360
rect 2282 90 2362 100
rect 2282 30 2292 90
rect 2352 80 2362 90
rect 2602 90 2682 100
rect 2602 80 2612 90
rect 2352 30 2612 80
rect 2672 30 2682 90
rect 2282 20 2682 30
rect 2740 440 3140 450
rect 2740 380 2750 440
rect 2810 390 3070 440
rect 2810 380 2820 390
rect 2740 370 2820 380
rect 3060 380 3070 390
rect 3130 380 3140 440
rect 3060 370 3140 380
rect 2740 100 2800 370
rect 3070 360 3140 370
rect 2880 310 2910 330
rect 2860 270 2910 310
rect 2970 310 3000 330
rect 2970 270 3020 310
rect 2860 200 3020 270
rect 2860 160 2910 200
rect 2880 140 2910 160
rect 2970 160 3020 200
rect 2970 140 3000 160
rect 3080 100 3140 360
rect 2740 90 2820 100
rect 2740 30 2750 90
rect 2810 80 2820 90
rect 3060 90 3140 100
rect 3060 80 3070 90
rect 2810 30 3070 80
rect 3130 30 3140 90
rect 2740 20 3140 30
rect 3196 440 3596 450
rect 3196 380 3206 440
rect 3266 390 3526 440
rect 3266 380 3276 390
rect 3196 370 3276 380
rect 3516 380 3526 390
rect 3586 380 3596 440
rect 3516 370 3596 380
rect 3196 100 3256 370
rect 3526 360 3596 370
rect 3336 310 3366 330
rect 3316 270 3366 310
rect 3426 310 3456 330
rect 3426 270 3476 310
rect 3316 200 3476 270
rect 3316 160 3366 200
rect 3336 140 3366 160
rect 3426 160 3476 200
rect 3426 140 3456 160
rect 3536 100 3596 360
rect 3196 90 3276 100
rect 3196 30 3206 90
rect 3266 80 3276 90
rect 3516 90 3596 100
rect 3516 80 3526 90
rect 3266 30 3526 80
rect 3586 30 3596 90
rect 3196 20 3596 30
rect 3652 440 4052 450
rect 3652 380 3662 440
rect 3722 390 3982 440
rect 3722 380 3732 390
rect 3652 370 3732 380
rect 3972 380 3982 390
rect 4042 380 4052 440
rect 3972 370 4052 380
rect 3652 100 3712 370
rect 3982 360 4052 370
rect 3792 310 3822 330
rect 3772 270 3822 310
rect 3882 310 3912 330
rect 3882 270 3932 310
rect 3772 200 3932 270
rect 3772 160 3822 200
rect 3792 140 3822 160
rect 3882 160 3932 200
rect 3882 140 3912 160
rect 3992 100 4052 360
rect 3652 90 3732 100
rect 3652 30 3662 90
rect 3722 80 3732 90
rect 3972 90 4052 100
rect 3972 80 3982 90
rect 3722 30 3982 80
rect 4042 30 4052 90
rect 3652 20 4052 30
rect 4110 440 4510 450
rect 4110 380 4120 440
rect 4180 390 4440 440
rect 4180 380 4190 390
rect 4110 370 4190 380
rect 4430 380 4440 390
rect 4500 380 4510 440
rect 4430 370 4510 380
rect 4110 100 4170 370
rect 4440 360 4510 370
rect 4250 310 4280 330
rect 4230 270 4280 310
rect 4340 310 4370 330
rect 4340 270 4390 310
rect 4230 200 4390 270
rect 4230 160 4280 200
rect 4250 140 4280 160
rect 4340 160 4390 200
rect 4340 140 4370 160
rect 4450 100 4510 360
rect 4110 90 4190 100
rect 4110 30 4120 90
rect 4180 80 4190 90
rect 4430 90 4510 100
rect 4430 80 4440 90
rect 4180 30 4440 80
rect 4500 30 4510 90
rect 4110 20 4510 30
rect 4566 440 4966 450
rect 4566 380 4576 440
rect 4636 390 4896 440
rect 4636 380 4646 390
rect 4566 370 4646 380
rect 4886 380 4896 390
rect 4956 380 4966 440
rect 4886 370 4966 380
rect 4566 100 4626 370
rect 4896 360 4966 370
rect 4706 310 4736 330
rect 4686 270 4736 310
rect 4796 310 4826 330
rect 4796 270 4846 310
rect 4686 200 4846 270
rect 4686 160 4736 200
rect 4706 140 4736 160
rect 4796 160 4846 200
rect 4796 140 4826 160
rect 4906 100 4966 360
rect 4566 90 4646 100
rect 4566 30 4576 90
rect 4636 80 4646 90
rect 4886 90 4966 100
rect 4886 80 4896 90
rect 4636 30 4896 80
rect 4956 30 4966 90
rect 4566 20 4966 30
rect 5022 440 5422 450
rect 5022 380 5032 440
rect 5092 390 5352 440
rect 5092 380 5102 390
rect 5022 370 5102 380
rect 5342 380 5352 390
rect 5412 380 5422 440
rect 5342 370 5422 380
rect 5022 100 5082 370
rect 5352 360 5422 370
rect 5162 310 5192 330
rect 5142 270 5192 310
rect 5252 310 5282 330
rect 5252 270 5302 310
rect 5142 200 5302 270
rect 5142 160 5192 200
rect 5162 140 5192 160
rect 5252 160 5302 200
rect 5252 140 5282 160
rect 5362 100 5422 360
rect 5022 90 5102 100
rect 5022 30 5032 90
rect 5092 80 5102 90
rect 5342 90 5422 100
rect 5342 80 5352 90
rect 5092 30 5352 80
rect 5412 30 5422 90
rect 5022 20 5422 30
rect 5480 440 5880 450
rect 5480 380 5490 440
rect 5550 390 5810 440
rect 5550 380 5560 390
rect 5480 370 5560 380
rect 5800 380 5810 390
rect 5870 380 5880 440
rect 5800 370 5880 380
rect 5480 100 5540 370
rect 5810 360 5880 370
rect 5620 310 5650 330
rect 5600 270 5650 310
rect 5710 310 5740 330
rect 5710 270 5760 310
rect 5600 200 5760 270
rect 5600 160 5650 200
rect 5620 140 5650 160
rect 5710 160 5760 200
rect 5710 140 5740 160
rect 5820 100 5880 360
rect 5480 90 5560 100
rect 5480 30 5490 90
rect 5550 80 5560 90
rect 5800 90 5880 100
rect 5800 80 5810 90
rect 5550 30 5810 80
rect 5870 30 5880 90
rect 5480 20 5880 30
rect 5936 440 6336 450
rect 5936 380 5946 440
rect 6006 390 6266 440
rect 6006 380 6016 390
rect 5936 370 6016 380
rect 6256 380 6266 390
rect 6326 380 6336 440
rect 6256 370 6336 380
rect 5936 100 5996 370
rect 6266 360 6336 370
rect 6076 310 6106 330
rect 6056 270 6106 310
rect 6166 310 6196 330
rect 6166 270 6216 310
rect 6056 200 6216 270
rect 6056 160 6106 200
rect 6076 140 6106 160
rect 6166 160 6216 200
rect 6166 140 6196 160
rect 6276 100 6336 360
rect 5936 90 6016 100
rect 5936 30 5946 90
rect 6006 80 6016 90
rect 6256 90 6336 100
rect 6256 80 6266 90
rect 6006 30 6266 80
rect 6326 30 6336 90
rect 5936 20 6336 30
rect 6392 440 6792 450
rect 6392 380 6402 440
rect 6462 390 6722 440
rect 6462 380 6472 390
rect 6392 370 6472 380
rect 6712 380 6722 390
rect 6782 380 6792 440
rect 6712 370 6792 380
rect 6392 100 6452 370
rect 6722 360 6792 370
rect 6532 310 6562 330
rect 6512 270 6562 310
rect 6622 310 6652 330
rect 6622 270 6672 310
rect 6512 200 6672 270
rect 6512 160 6562 200
rect 6532 140 6562 160
rect 6622 160 6672 200
rect 6622 140 6652 160
rect 6732 100 6792 360
rect 6392 90 6472 100
rect 6392 30 6402 90
rect 6462 80 6472 90
rect 6712 90 6792 100
rect 6712 80 6722 90
rect 6462 30 6722 80
rect 6782 30 6792 90
rect 6392 20 6792 30
rect 6850 440 7250 450
rect 6850 380 6860 440
rect 6920 390 7180 440
rect 6920 380 6930 390
rect 6850 370 6930 380
rect 7170 380 7180 390
rect 7240 380 7250 440
rect 7170 370 7250 380
rect 6850 100 6910 370
rect 7180 360 7250 370
rect 6990 310 7020 330
rect 6970 270 7020 310
rect 7080 310 7110 330
rect 7080 270 7130 310
rect 6970 200 7130 270
rect 6970 160 7020 200
rect 6990 140 7020 160
rect 7080 160 7130 200
rect 7080 140 7110 160
rect 7190 100 7250 360
rect 6850 90 6930 100
rect 6850 30 6860 90
rect 6920 80 6930 90
rect 7170 90 7250 100
rect 7170 80 7180 90
rect 6920 30 7180 80
rect 7240 30 7250 90
rect 6850 20 7250 30
rect 7306 440 7706 450
rect 7306 380 7316 440
rect 7376 390 7636 440
rect 7376 380 7386 390
rect 7306 370 7386 380
rect 7626 380 7636 390
rect 7696 380 7706 440
rect 7626 370 7706 380
rect 7306 100 7366 370
rect 7636 360 7706 370
rect 7446 310 7476 330
rect 7426 270 7476 310
rect 7536 310 7566 330
rect 7536 270 7586 310
rect 7426 200 7586 270
rect 7426 160 7476 200
rect 7446 140 7476 160
rect 7536 160 7586 200
rect 7536 140 7566 160
rect 7646 100 7706 360
rect 7306 90 7386 100
rect 7306 30 7316 90
rect 7376 80 7386 90
rect 7626 90 7706 100
rect 7626 80 7636 90
rect 7376 30 7636 80
rect 7696 30 7706 90
rect 7306 20 7706 30
rect 7762 440 8162 450
rect 7762 380 7772 440
rect 7832 390 8092 440
rect 7832 380 7842 390
rect 7762 370 7842 380
rect 8082 380 8092 390
rect 8152 380 8162 440
rect 8082 370 8162 380
rect 7762 100 7822 370
rect 8092 360 8162 370
rect 7902 310 7932 330
rect 7882 270 7932 310
rect 7992 310 8022 330
rect 7992 270 8042 310
rect 7882 200 8042 270
rect 7882 160 7932 200
rect 7902 140 7932 160
rect 7992 160 8042 200
rect 7992 140 8022 160
rect 8102 100 8162 360
rect 7762 90 7842 100
rect 7762 30 7772 90
rect 7832 80 7842 90
rect 8082 90 8162 100
rect 8082 80 8092 90
rect 7832 30 8092 80
rect 8152 30 8162 90
rect 7762 20 8162 30
rect 8236 440 8636 450
rect 8236 380 8246 440
rect 8306 390 8566 440
rect 8306 380 8316 390
rect 8236 370 8316 380
rect 8556 380 8566 390
rect 8626 380 8636 440
rect 8556 370 8636 380
rect 8236 100 8296 370
rect 8566 360 8636 370
rect 8376 310 8406 330
rect 8356 270 8406 310
rect 8466 310 8496 330
rect 8466 270 8516 310
rect 8356 200 8516 270
rect 8356 160 8406 200
rect 8376 140 8406 160
rect 8466 160 8516 200
rect 8466 140 8496 160
rect 8576 100 8636 360
rect 8236 90 8316 100
rect 8236 30 8246 90
rect 8306 80 8316 90
rect 8556 90 8636 100
rect 8556 80 8566 90
rect 8306 30 8566 80
rect 8626 30 8636 90
rect 8236 20 8636 30
rect 8692 440 9092 450
rect 8692 380 8702 440
rect 8762 390 9022 440
rect 8762 380 8772 390
rect 8692 370 8772 380
rect 9012 380 9022 390
rect 9082 380 9092 440
rect 9012 370 9092 380
rect 8692 100 8752 370
rect 9022 360 9092 370
rect 8832 310 8862 330
rect 8812 270 8862 310
rect 8922 310 8952 330
rect 8922 270 8972 310
rect 8812 200 8972 270
rect 8812 160 8862 200
rect 8832 140 8862 160
rect 8922 160 8972 200
rect 8922 140 8952 160
rect 9032 100 9092 360
rect 8692 90 8772 100
rect 8692 30 8702 90
rect 8762 80 8772 90
rect 9012 90 9092 100
rect 9012 80 9022 90
rect 8762 30 9022 80
rect 9082 30 9092 90
rect 8692 20 9092 30
rect 9150 440 9550 450
rect 9150 380 9160 440
rect 9220 390 9480 440
rect 9220 380 9230 390
rect 9150 370 9230 380
rect 9470 380 9480 390
rect 9540 380 9550 440
rect 9470 370 9550 380
rect 9150 100 9210 370
rect 9480 360 9550 370
rect 9290 310 9320 330
rect 9270 270 9320 310
rect 9380 310 9410 330
rect 9380 270 9430 310
rect 9270 200 9430 270
rect 9270 160 9320 200
rect 9290 140 9320 160
rect 9380 160 9430 200
rect 9380 140 9410 160
rect 9490 100 9550 360
rect 9150 90 9230 100
rect 9150 30 9160 90
rect 9220 80 9230 90
rect 9470 90 9550 100
rect 9470 80 9480 90
rect 9220 30 9480 80
rect 9540 30 9550 90
rect 9150 20 9550 30
rect 9606 440 10006 450
rect 9606 380 9616 440
rect 9676 390 9936 440
rect 9676 380 9686 390
rect 9606 370 9686 380
rect 9926 380 9936 390
rect 9996 380 10006 440
rect 9926 370 10006 380
rect 9606 100 9666 370
rect 9936 360 10006 370
rect 9746 310 9776 330
rect 9726 270 9776 310
rect 9836 310 9866 330
rect 9836 270 9886 310
rect 9726 200 9886 270
rect 9726 160 9776 200
rect 9746 140 9776 160
rect 9836 160 9886 200
rect 9836 140 9866 160
rect 9946 100 10006 360
rect 9606 90 9686 100
rect 9606 30 9616 90
rect 9676 80 9686 90
rect 9926 90 10006 100
rect 9926 80 9936 90
rect 9676 30 9936 80
rect 9996 30 10006 90
rect 9606 20 10006 30
rect 10062 440 10462 450
rect 10062 380 10072 440
rect 10132 390 10392 440
rect 10132 380 10142 390
rect 10062 370 10142 380
rect 10382 380 10392 390
rect 10452 380 10462 440
rect 10382 370 10462 380
rect 10062 100 10122 370
rect 10392 360 10462 370
rect 10202 310 10232 330
rect 10182 270 10232 310
rect 10292 310 10322 330
rect 10292 270 10342 310
rect 10182 200 10342 270
rect 10182 160 10232 200
rect 10202 140 10232 160
rect 10292 160 10342 200
rect 10292 140 10322 160
rect 10402 100 10462 360
rect 10062 90 10142 100
rect 10062 30 10072 90
rect 10132 80 10142 90
rect 10382 90 10462 100
rect 10382 80 10392 90
rect 10132 30 10392 80
rect 10452 30 10462 90
rect 10062 20 10462 30
rect 10520 440 10920 450
rect 10520 380 10530 440
rect 10590 390 10850 440
rect 10590 380 10600 390
rect 10520 370 10600 380
rect 10840 380 10850 390
rect 10910 380 10920 440
rect 10840 370 10920 380
rect 10520 100 10580 370
rect 10850 360 10920 370
rect 10660 310 10690 330
rect 10640 270 10690 310
rect 10750 310 10780 330
rect 10750 270 10800 310
rect 10640 200 10800 270
rect 10640 160 10690 200
rect 10660 140 10690 160
rect 10750 160 10800 200
rect 10750 140 10780 160
rect 10860 100 10920 360
rect 10520 90 10600 100
rect 10520 30 10530 90
rect 10590 80 10600 90
rect 10840 90 10920 100
rect 10840 80 10850 90
rect 10590 30 10850 80
rect 10910 30 10920 90
rect 10520 20 10920 30
rect 10976 440 11376 450
rect 10976 380 10986 440
rect 11046 390 11306 440
rect 11046 380 11056 390
rect 10976 370 11056 380
rect 11296 380 11306 390
rect 11366 380 11376 440
rect 11296 370 11376 380
rect 10976 100 11036 370
rect 11306 360 11376 370
rect 11116 310 11146 330
rect 11096 270 11146 310
rect 11206 310 11236 330
rect 11206 270 11256 310
rect 11096 200 11256 270
rect 11096 160 11146 200
rect 11116 140 11146 160
rect 11206 160 11256 200
rect 11206 140 11236 160
rect 11316 100 11376 360
rect 10976 90 11056 100
rect 10976 30 10986 90
rect 11046 80 11056 90
rect 11296 90 11376 100
rect 11296 80 11306 90
rect 11046 30 11306 80
rect 11366 30 11376 90
rect 10976 20 11376 30
rect 11432 440 11832 450
rect 11432 380 11442 440
rect 11502 390 11762 440
rect 11502 380 11512 390
rect 11432 370 11512 380
rect 11752 380 11762 390
rect 11822 380 11832 440
rect 11752 370 11832 380
rect 11432 100 11492 370
rect 11762 360 11832 370
rect 11572 310 11602 330
rect 11552 270 11602 310
rect 11662 310 11692 330
rect 11662 270 11712 310
rect 11552 200 11712 270
rect 11552 160 11602 200
rect 11572 140 11602 160
rect 11662 160 11712 200
rect 11662 140 11692 160
rect 11772 100 11832 360
rect 11432 90 11512 100
rect 11432 30 11442 90
rect 11502 80 11512 90
rect 11752 90 11832 100
rect 11752 80 11762 90
rect 11502 30 11762 80
rect 11822 30 11832 90
rect 11432 20 11832 30
rect 11890 440 12290 450
rect 11890 380 11900 440
rect 11960 390 12220 440
rect 11960 380 11970 390
rect 11890 370 11970 380
rect 12210 380 12220 390
rect 12280 380 12290 440
rect 12210 370 12290 380
rect 11890 100 11950 370
rect 12220 360 12290 370
rect 12030 310 12060 330
rect 12010 270 12060 310
rect 12120 310 12150 330
rect 12120 270 12170 310
rect 12010 200 12170 270
rect 12010 160 12060 200
rect 12030 140 12060 160
rect 12120 160 12170 200
rect 12120 140 12150 160
rect 12230 100 12290 360
rect 11890 90 11970 100
rect 11890 30 11900 90
rect 11960 80 11970 90
rect 12210 90 12290 100
rect 12210 80 12220 90
rect 11960 30 12220 80
rect 12280 30 12290 90
rect 11890 20 12290 30
rect 12346 440 12746 450
rect 12346 380 12356 440
rect 12416 390 12676 440
rect 12416 380 12426 390
rect 12346 370 12426 380
rect 12666 380 12676 390
rect 12736 380 12746 440
rect 12666 370 12746 380
rect 12346 100 12406 370
rect 12676 360 12746 370
rect 12486 310 12516 330
rect 12466 270 12516 310
rect 12576 310 12606 330
rect 12576 270 12626 310
rect 12466 200 12626 270
rect 12466 160 12516 200
rect 12486 140 12516 160
rect 12576 160 12626 200
rect 12576 140 12606 160
rect 12686 100 12746 360
rect 12346 90 12426 100
rect 12346 30 12356 90
rect 12416 80 12426 90
rect 12666 90 12746 100
rect 12666 80 12676 90
rect 12416 30 12676 80
rect 12736 30 12746 90
rect 12346 20 12746 30
rect 12802 440 13202 450
rect 12802 380 12812 440
rect 12872 390 13132 440
rect 12872 380 12882 390
rect 12802 370 12882 380
rect 13122 380 13132 390
rect 13192 380 13202 440
rect 13122 370 13202 380
rect 12802 100 12862 370
rect 13132 360 13202 370
rect 12942 310 12972 330
rect 12922 270 12972 310
rect 13032 310 13062 330
rect 13032 270 13082 310
rect 12922 200 13082 270
rect 12922 160 12972 200
rect 12942 140 12972 160
rect 13032 160 13082 200
rect 13032 140 13062 160
rect 13142 100 13202 360
rect 12802 90 12882 100
rect 12802 30 12812 90
rect 12872 80 12882 90
rect 13122 90 13202 100
rect 13122 80 13132 90
rect 12872 30 13132 80
rect 13192 30 13202 90
rect 12802 20 13202 30
rect 13260 440 13660 450
rect 13260 380 13270 440
rect 13330 390 13590 440
rect 13330 380 13340 390
rect 13260 370 13340 380
rect 13580 380 13590 390
rect 13650 380 13660 440
rect 13580 370 13660 380
rect 13260 100 13320 370
rect 13590 360 13660 370
rect 13400 310 13430 330
rect 13380 270 13430 310
rect 13490 310 13520 330
rect 13490 270 13540 310
rect 13380 200 13540 270
rect 13380 160 13430 200
rect 13400 140 13430 160
rect 13490 160 13540 200
rect 13490 140 13520 160
rect 13600 100 13660 360
rect 13260 90 13340 100
rect 13260 30 13270 90
rect 13330 80 13340 90
rect 13580 90 13660 100
rect 13580 80 13590 90
rect 13330 30 13590 80
rect 13650 30 13660 90
rect 13260 20 13660 30
rect 13716 440 14116 450
rect 13716 380 13726 440
rect 13786 390 14046 440
rect 13786 380 13796 390
rect 13716 370 13796 380
rect 14036 380 14046 390
rect 14106 380 14116 440
rect 14036 370 14116 380
rect 13716 100 13776 370
rect 14046 360 14116 370
rect 13856 310 13886 330
rect 13836 270 13886 310
rect 13946 310 13976 330
rect 13946 270 13996 310
rect 13836 200 13996 270
rect 13836 160 13886 200
rect 13856 140 13886 160
rect 13946 160 13996 200
rect 13946 140 13976 160
rect 14056 100 14116 360
rect 13716 90 13796 100
rect 13716 30 13726 90
rect 13786 80 13796 90
rect 14036 90 14116 100
rect 14036 80 14046 90
rect 13786 30 14046 80
rect 14106 30 14116 90
rect 13716 20 14116 30
rect 14172 440 14572 450
rect 14172 380 14182 440
rect 14242 390 14502 440
rect 14242 380 14252 390
rect 14172 370 14252 380
rect 14492 380 14502 390
rect 14562 380 14572 440
rect 14492 370 14572 380
rect 14172 100 14232 370
rect 14502 360 14572 370
rect 14312 310 14342 330
rect 14292 270 14342 310
rect 14402 310 14432 330
rect 14402 270 14452 310
rect 14292 200 14452 270
rect 14292 160 14342 200
rect 14312 140 14342 160
rect 14402 160 14452 200
rect 14402 140 14432 160
rect 14512 100 14572 360
rect 14172 90 14252 100
rect 14172 30 14182 90
rect 14242 80 14252 90
rect 14492 90 14572 100
rect 14492 80 14502 90
rect 14242 30 14502 80
rect 14562 30 14572 90
rect 14172 20 14572 30
rect 14630 440 15030 450
rect 14630 380 14640 440
rect 14700 390 14960 440
rect 14700 380 14710 390
rect 14630 370 14710 380
rect 14950 380 14960 390
rect 15020 380 15030 440
rect 14950 370 15030 380
rect 14630 100 14690 370
rect 14960 360 15030 370
rect 14770 310 14800 330
rect 14750 270 14800 310
rect 14860 310 14890 330
rect 14860 270 14910 310
rect 14750 200 14910 270
rect 14750 160 14800 200
rect 14770 140 14800 160
rect 14860 160 14910 200
rect 14860 140 14890 160
rect 14970 100 15030 360
rect 14630 90 14710 100
rect 14630 30 14640 90
rect 14700 80 14710 90
rect 14950 90 15030 100
rect 14950 80 14960 90
rect 14700 30 14960 80
rect 15020 30 15030 90
rect 14630 20 15030 30
rect 15086 440 15486 450
rect 15086 380 15096 440
rect 15156 390 15416 440
rect 15156 380 15166 390
rect 15086 370 15166 380
rect 15406 380 15416 390
rect 15476 380 15486 440
rect 15406 370 15486 380
rect 15086 100 15146 370
rect 15416 360 15486 370
rect 15226 310 15256 330
rect 15206 270 15256 310
rect 15316 310 15346 330
rect 15316 270 15366 310
rect 15206 200 15366 270
rect 15206 160 15256 200
rect 15226 140 15256 160
rect 15316 160 15366 200
rect 15316 140 15346 160
rect 15426 100 15486 360
rect 15086 90 15166 100
rect 15086 30 15096 90
rect 15156 80 15166 90
rect 15406 90 15486 100
rect 15406 80 15416 90
rect 15156 30 15416 80
rect 15476 30 15486 90
rect 15086 20 15486 30
rect 0 -52 400 -42
rect 0 -112 10 -52
rect 70 -102 330 -52
rect 70 -112 80 -102
rect 0 -122 80 -112
rect 320 -112 330 -102
rect 390 -112 400 -52
rect 320 -122 400 -112
rect 0 -392 60 -122
rect 330 -132 400 -122
rect 140 -182 170 -162
rect 120 -222 170 -182
rect 230 -182 260 -162
rect 230 -222 280 -182
rect 120 -292 280 -222
rect 120 -332 170 -292
rect 140 -352 170 -332
rect 230 -332 280 -292
rect 230 -352 260 -332
rect 340 -392 400 -132
rect 0 -402 80 -392
rect 0 -462 10 -402
rect 70 -412 80 -402
rect 320 -402 400 -392
rect 320 -412 330 -402
rect 70 -462 330 -412
rect 390 -462 400 -402
rect 0 -472 400 -462
rect 456 -52 856 -42
rect 456 -112 466 -52
rect 526 -102 786 -52
rect 526 -112 536 -102
rect 456 -122 536 -112
rect 776 -112 786 -102
rect 846 -112 856 -52
rect 776 -122 856 -112
rect 456 -392 516 -122
rect 786 -132 856 -122
rect 596 -182 626 -162
rect 576 -222 626 -182
rect 686 -182 716 -162
rect 686 -222 736 -182
rect 576 -292 736 -222
rect 576 -332 626 -292
rect 596 -352 626 -332
rect 686 -332 736 -292
rect 686 -352 716 -332
rect 796 -392 856 -132
rect 456 -402 536 -392
rect 456 -462 466 -402
rect 526 -412 536 -402
rect 776 -402 856 -392
rect 776 -412 786 -402
rect 526 -462 786 -412
rect 846 -462 856 -402
rect 456 -472 856 -462
rect 912 -52 1312 -42
rect 912 -112 922 -52
rect 982 -102 1242 -52
rect 982 -112 992 -102
rect 912 -122 992 -112
rect 1232 -112 1242 -102
rect 1302 -112 1312 -52
rect 1232 -122 1312 -112
rect 912 -392 972 -122
rect 1242 -132 1312 -122
rect 1052 -182 1082 -162
rect 1032 -222 1082 -182
rect 1142 -182 1172 -162
rect 1142 -222 1192 -182
rect 1032 -292 1192 -222
rect 1032 -332 1082 -292
rect 1052 -352 1082 -332
rect 1142 -332 1192 -292
rect 1142 -352 1172 -332
rect 1252 -392 1312 -132
rect 912 -402 992 -392
rect 912 -462 922 -402
rect 982 -412 992 -402
rect 1232 -402 1312 -392
rect 1232 -412 1242 -402
rect 982 -462 1242 -412
rect 1302 -462 1312 -402
rect 912 -472 1312 -462
rect 1370 -52 1770 -42
rect 1370 -112 1380 -52
rect 1440 -102 1700 -52
rect 1440 -112 1450 -102
rect 1370 -122 1450 -112
rect 1690 -112 1700 -102
rect 1760 -112 1770 -52
rect 1690 -122 1770 -112
rect 1370 -392 1430 -122
rect 1700 -132 1770 -122
rect 1510 -182 1540 -162
rect 1490 -222 1540 -182
rect 1600 -182 1630 -162
rect 1600 -222 1650 -182
rect 1490 -292 1650 -222
rect 1490 -332 1540 -292
rect 1510 -352 1540 -332
rect 1600 -332 1650 -292
rect 1600 -352 1630 -332
rect 1710 -392 1770 -132
rect 1370 -402 1450 -392
rect 1370 -462 1380 -402
rect 1440 -412 1450 -402
rect 1690 -402 1770 -392
rect 1690 -412 1700 -402
rect 1440 -462 1700 -412
rect 1760 -462 1770 -402
rect 1370 -472 1770 -462
rect 1826 -52 2226 -42
rect 1826 -112 1836 -52
rect 1896 -102 2156 -52
rect 1896 -112 1906 -102
rect 1826 -122 1906 -112
rect 2146 -112 2156 -102
rect 2216 -112 2226 -52
rect 2146 -122 2226 -112
rect 1826 -392 1886 -122
rect 2156 -132 2226 -122
rect 1966 -182 1996 -162
rect 1946 -222 1996 -182
rect 2056 -182 2086 -162
rect 2056 -222 2106 -182
rect 1946 -292 2106 -222
rect 1946 -332 1996 -292
rect 1966 -352 1996 -332
rect 2056 -332 2106 -292
rect 2056 -352 2086 -332
rect 2166 -392 2226 -132
rect 1826 -402 1906 -392
rect 1826 -462 1836 -402
rect 1896 -412 1906 -402
rect 2146 -402 2226 -392
rect 2146 -412 2156 -402
rect 1896 -462 2156 -412
rect 2216 -462 2226 -402
rect 1826 -472 2226 -462
rect 2282 -52 2682 -42
rect 2282 -112 2292 -52
rect 2352 -102 2612 -52
rect 2352 -112 2362 -102
rect 2282 -122 2362 -112
rect 2602 -112 2612 -102
rect 2672 -112 2682 -52
rect 2602 -122 2682 -112
rect 2282 -392 2342 -122
rect 2612 -132 2682 -122
rect 2422 -182 2452 -162
rect 2402 -222 2452 -182
rect 2512 -182 2542 -162
rect 2512 -222 2562 -182
rect 2402 -292 2562 -222
rect 2402 -332 2452 -292
rect 2422 -352 2452 -332
rect 2512 -332 2562 -292
rect 2512 -352 2542 -332
rect 2622 -392 2682 -132
rect 2282 -402 2362 -392
rect 2282 -462 2292 -402
rect 2352 -412 2362 -402
rect 2602 -402 2682 -392
rect 2602 -412 2612 -402
rect 2352 -462 2612 -412
rect 2672 -462 2682 -402
rect 2282 -472 2682 -462
rect 2740 -52 3140 -42
rect 2740 -112 2750 -52
rect 2810 -102 3070 -52
rect 2810 -112 2820 -102
rect 2740 -122 2820 -112
rect 3060 -112 3070 -102
rect 3130 -112 3140 -52
rect 3060 -122 3140 -112
rect 2740 -392 2800 -122
rect 3070 -132 3140 -122
rect 2880 -182 2910 -162
rect 2860 -222 2910 -182
rect 2970 -182 3000 -162
rect 2970 -222 3020 -182
rect 2860 -292 3020 -222
rect 2860 -332 2910 -292
rect 2880 -352 2910 -332
rect 2970 -332 3020 -292
rect 2970 -352 3000 -332
rect 3080 -392 3140 -132
rect 2740 -402 2820 -392
rect 2740 -462 2750 -402
rect 2810 -412 2820 -402
rect 3060 -402 3140 -392
rect 3060 -412 3070 -402
rect 2810 -462 3070 -412
rect 3130 -462 3140 -402
rect 2740 -472 3140 -462
rect 3196 -52 3596 -42
rect 3196 -112 3206 -52
rect 3266 -102 3526 -52
rect 3266 -112 3276 -102
rect 3196 -122 3276 -112
rect 3516 -112 3526 -102
rect 3586 -112 3596 -52
rect 3516 -122 3596 -112
rect 3196 -392 3256 -122
rect 3526 -132 3596 -122
rect 3336 -182 3366 -162
rect 3316 -222 3366 -182
rect 3426 -182 3456 -162
rect 3426 -222 3476 -182
rect 3316 -292 3476 -222
rect 3316 -332 3366 -292
rect 3336 -352 3366 -332
rect 3426 -332 3476 -292
rect 3426 -352 3456 -332
rect 3536 -392 3596 -132
rect 3196 -402 3276 -392
rect 3196 -462 3206 -402
rect 3266 -412 3276 -402
rect 3516 -402 3596 -392
rect 3516 -412 3526 -402
rect 3266 -462 3526 -412
rect 3586 -462 3596 -402
rect 3196 -472 3596 -462
rect 3652 -52 4052 -42
rect 3652 -112 3662 -52
rect 3722 -102 3982 -52
rect 3722 -112 3732 -102
rect 3652 -122 3732 -112
rect 3972 -112 3982 -102
rect 4042 -112 4052 -52
rect 3972 -122 4052 -112
rect 3652 -392 3712 -122
rect 3982 -132 4052 -122
rect 3792 -182 3822 -162
rect 3772 -222 3822 -182
rect 3882 -182 3912 -162
rect 3882 -222 3932 -182
rect 3772 -292 3932 -222
rect 3772 -332 3822 -292
rect 3792 -352 3822 -332
rect 3882 -332 3932 -292
rect 3882 -352 3912 -332
rect 3992 -392 4052 -132
rect 3652 -402 3732 -392
rect 3652 -462 3662 -402
rect 3722 -412 3732 -402
rect 3972 -402 4052 -392
rect 3972 -412 3982 -402
rect 3722 -462 3982 -412
rect 4042 -462 4052 -402
rect 3652 -472 4052 -462
rect 4110 -52 4510 -42
rect 4110 -112 4120 -52
rect 4180 -102 4440 -52
rect 4180 -112 4190 -102
rect 4110 -122 4190 -112
rect 4430 -112 4440 -102
rect 4500 -112 4510 -52
rect 4430 -122 4510 -112
rect 4110 -392 4170 -122
rect 4440 -132 4510 -122
rect 4250 -182 4280 -162
rect 4230 -222 4280 -182
rect 4340 -182 4370 -162
rect 4340 -222 4390 -182
rect 4230 -292 4390 -222
rect 4230 -332 4280 -292
rect 4250 -352 4280 -332
rect 4340 -332 4390 -292
rect 4340 -352 4370 -332
rect 4450 -392 4510 -132
rect 4110 -402 4190 -392
rect 4110 -462 4120 -402
rect 4180 -412 4190 -402
rect 4430 -402 4510 -392
rect 4430 -412 4440 -402
rect 4180 -462 4440 -412
rect 4500 -462 4510 -402
rect 4110 -472 4510 -462
rect 4566 -52 4966 -42
rect 4566 -112 4576 -52
rect 4636 -102 4896 -52
rect 4636 -112 4646 -102
rect 4566 -122 4646 -112
rect 4886 -112 4896 -102
rect 4956 -112 4966 -52
rect 4886 -122 4966 -112
rect 4566 -392 4626 -122
rect 4896 -132 4966 -122
rect 4706 -182 4736 -162
rect 4686 -222 4736 -182
rect 4796 -182 4826 -162
rect 4796 -222 4846 -182
rect 4686 -292 4846 -222
rect 4686 -332 4736 -292
rect 4706 -352 4736 -332
rect 4796 -332 4846 -292
rect 4796 -352 4826 -332
rect 4906 -392 4966 -132
rect 4566 -402 4646 -392
rect 4566 -462 4576 -402
rect 4636 -412 4646 -402
rect 4886 -402 4966 -392
rect 4886 -412 4896 -402
rect 4636 -462 4896 -412
rect 4956 -462 4966 -402
rect 4566 -472 4966 -462
rect 5022 -52 5422 -42
rect 5022 -112 5032 -52
rect 5092 -102 5352 -52
rect 5092 -112 5102 -102
rect 5022 -122 5102 -112
rect 5342 -112 5352 -102
rect 5412 -112 5422 -52
rect 5342 -122 5422 -112
rect 5022 -392 5082 -122
rect 5352 -132 5422 -122
rect 5162 -182 5192 -162
rect 5142 -222 5192 -182
rect 5252 -182 5282 -162
rect 5252 -222 5302 -182
rect 5142 -292 5302 -222
rect 5142 -332 5192 -292
rect 5162 -352 5192 -332
rect 5252 -332 5302 -292
rect 5252 -352 5282 -332
rect 5362 -392 5422 -132
rect 5022 -402 5102 -392
rect 5022 -462 5032 -402
rect 5092 -412 5102 -402
rect 5342 -402 5422 -392
rect 5342 -412 5352 -402
rect 5092 -462 5352 -412
rect 5412 -462 5422 -402
rect 5022 -472 5422 -462
rect 5480 -52 5880 -42
rect 5480 -112 5490 -52
rect 5550 -102 5810 -52
rect 5550 -112 5560 -102
rect 5480 -122 5560 -112
rect 5800 -112 5810 -102
rect 5870 -112 5880 -52
rect 5800 -122 5880 -112
rect 5480 -392 5540 -122
rect 5810 -132 5880 -122
rect 5620 -182 5650 -162
rect 5600 -222 5650 -182
rect 5710 -182 5740 -162
rect 5710 -222 5760 -182
rect 5600 -292 5760 -222
rect 5600 -332 5650 -292
rect 5620 -352 5650 -332
rect 5710 -332 5760 -292
rect 5710 -352 5740 -332
rect 5820 -392 5880 -132
rect 5480 -402 5560 -392
rect 5480 -462 5490 -402
rect 5550 -412 5560 -402
rect 5800 -402 5880 -392
rect 5800 -412 5810 -402
rect 5550 -462 5810 -412
rect 5870 -462 5880 -402
rect 5480 -472 5880 -462
rect 5936 -52 6336 -42
rect 5936 -112 5946 -52
rect 6006 -102 6266 -52
rect 6006 -112 6016 -102
rect 5936 -122 6016 -112
rect 6256 -112 6266 -102
rect 6326 -112 6336 -52
rect 6256 -122 6336 -112
rect 5936 -392 5996 -122
rect 6266 -132 6336 -122
rect 6076 -182 6106 -162
rect 6056 -222 6106 -182
rect 6166 -182 6196 -162
rect 6166 -222 6216 -182
rect 6056 -292 6216 -222
rect 6056 -332 6106 -292
rect 6076 -352 6106 -332
rect 6166 -332 6216 -292
rect 6166 -352 6196 -332
rect 6276 -392 6336 -132
rect 5936 -402 6016 -392
rect 5936 -462 5946 -402
rect 6006 -412 6016 -402
rect 6256 -402 6336 -392
rect 6256 -412 6266 -402
rect 6006 -462 6266 -412
rect 6326 -462 6336 -402
rect 5936 -472 6336 -462
rect 6392 -52 6792 -42
rect 6392 -112 6402 -52
rect 6462 -102 6722 -52
rect 6462 -112 6472 -102
rect 6392 -122 6472 -112
rect 6712 -112 6722 -102
rect 6782 -112 6792 -52
rect 6712 -122 6792 -112
rect 6392 -392 6452 -122
rect 6722 -132 6792 -122
rect 6532 -182 6562 -162
rect 6512 -222 6562 -182
rect 6622 -182 6652 -162
rect 6622 -222 6672 -182
rect 6512 -292 6672 -222
rect 6512 -332 6562 -292
rect 6532 -352 6562 -332
rect 6622 -332 6672 -292
rect 6622 -352 6652 -332
rect 6732 -392 6792 -132
rect 6392 -402 6472 -392
rect 6392 -462 6402 -402
rect 6462 -412 6472 -402
rect 6712 -402 6792 -392
rect 6712 -412 6722 -402
rect 6462 -462 6722 -412
rect 6782 -462 6792 -402
rect 6392 -472 6792 -462
rect 6850 -52 7250 -42
rect 6850 -112 6860 -52
rect 6920 -102 7180 -52
rect 6920 -112 6930 -102
rect 6850 -122 6930 -112
rect 7170 -112 7180 -102
rect 7240 -112 7250 -52
rect 7170 -122 7250 -112
rect 6850 -392 6910 -122
rect 7180 -132 7250 -122
rect 6990 -182 7020 -162
rect 6970 -222 7020 -182
rect 7080 -182 7110 -162
rect 7080 -222 7130 -182
rect 6970 -292 7130 -222
rect 6970 -332 7020 -292
rect 6990 -352 7020 -332
rect 7080 -332 7130 -292
rect 7080 -352 7110 -332
rect 7190 -392 7250 -132
rect 6850 -402 6930 -392
rect 6850 -462 6860 -402
rect 6920 -412 6930 -402
rect 7170 -402 7250 -392
rect 7170 -412 7180 -402
rect 6920 -462 7180 -412
rect 7240 -462 7250 -402
rect 6850 -472 7250 -462
rect 7306 -52 7706 -42
rect 7306 -112 7316 -52
rect 7376 -102 7636 -52
rect 7376 -112 7386 -102
rect 7306 -122 7386 -112
rect 7626 -112 7636 -102
rect 7696 -112 7706 -52
rect 7626 -122 7706 -112
rect 7306 -392 7366 -122
rect 7636 -132 7706 -122
rect 7446 -182 7476 -162
rect 7426 -222 7476 -182
rect 7536 -182 7566 -162
rect 7536 -222 7586 -182
rect 7426 -292 7586 -222
rect 7426 -332 7476 -292
rect 7446 -352 7476 -332
rect 7536 -332 7586 -292
rect 7536 -352 7566 -332
rect 7646 -392 7706 -132
rect 7306 -402 7386 -392
rect 7306 -462 7316 -402
rect 7376 -412 7386 -402
rect 7626 -402 7706 -392
rect 7626 -412 7636 -402
rect 7376 -462 7636 -412
rect 7696 -462 7706 -402
rect 7306 -472 7706 -462
rect 7762 -52 8162 -42
rect 7762 -112 7772 -52
rect 7832 -102 8092 -52
rect 7832 -112 7842 -102
rect 7762 -122 7842 -112
rect 8082 -112 8092 -102
rect 8152 -112 8162 -52
rect 8082 -122 8162 -112
rect 7762 -392 7822 -122
rect 8092 -132 8162 -122
rect 7902 -182 7932 -162
rect 7882 -222 7932 -182
rect 7992 -182 8022 -162
rect 7992 -222 8042 -182
rect 7882 -292 8042 -222
rect 7882 -332 7932 -292
rect 7902 -352 7932 -332
rect 7992 -332 8042 -292
rect 7992 -352 8022 -332
rect 8102 -392 8162 -132
rect 7762 -402 7842 -392
rect 7762 -462 7772 -402
rect 7832 -412 7842 -402
rect 8082 -402 8162 -392
rect 8082 -412 8092 -402
rect 7832 -462 8092 -412
rect 8152 -462 8162 -402
rect 7762 -472 8162 -462
rect 8236 -52 8636 -42
rect 8236 -112 8246 -52
rect 8306 -102 8566 -52
rect 8306 -112 8316 -102
rect 8236 -122 8316 -112
rect 8556 -112 8566 -102
rect 8626 -112 8636 -52
rect 8556 -122 8636 -112
rect 8236 -392 8296 -122
rect 8566 -132 8636 -122
rect 8376 -182 8406 -162
rect 8356 -222 8406 -182
rect 8466 -182 8496 -162
rect 8466 -222 8516 -182
rect 8356 -292 8516 -222
rect 8356 -332 8406 -292
rect 8376 -352 8406 -332
rect 8466 -332 8516 -292
rect 8466 -352 8496 -332
rect 8576 -392 8636 -132
rect 8236 -402 8316 -392
rect 8236 -462 8246 -402
rect 8306 -412 8316 -402
rect 8556 -402 8636 -392
rect 8556 -412 8566 -402
rect 8306 -462 8566 -412
rect 8626 -462 8636 -402
rect 8236 -472 8636 -462
rect 8692 -52 9092 -42
rect 8692 -112 8702 -52
rect 8762 -102 9022 -52
rect 8762 -112 8772 -102
rect 8692 -122 8772 -112
rect 9012 -112 9022 -102
rect 9082 -112 9092 -52
rect 9012 -122 9092 -112
rect 8692 -392 8752 -122
rect 9022 -132 9092 -122
rect 8832 -182 8862 -162
rect 8812 -222 8862 -182
rect 8922 -182 8952 -162
rect 8922 -222 8972 -182
rect 8812 -292 8972 -222
rect 8812 -332 8862 -292
rect 8832 -352 8862 -332
rect 8922 -332 8972 -292
rect 8922 -352 8952 -332
rect 9032 -392 9092 -132
rect 8692 -402 8772 -392
rect 8692 -462 8702 -402
rect 8762 -412 8772 -402
rect 9012 -402 9092 -392
rect 9012 -412 9022 -402
rect 8762 -462 9022 -412
rect 9082 -462 9092 -402
rect 8692 -472 9092 -462
rect 9150 -52 9550 -42
rect 9150 -112 9160 -52
rect 9220 -102 9480 -52
rect 9220 -112 9230 -102
rect 9150 -122 9230 -112
rect 9470 -112 9480 -102
rect 9540 -112 9550 -52
rect 9470 -122 9550 -112
rect 9150 -392 9210 -122
rect 9480 -132 9550 -122
rect 9290 -182 9320 -162
rect 9270 -222 9320 -182
rect 9380 -182 9410 -162
rect 9380 -222 9430 -182
rect 9270 -292 9430 -222
rect 9270 -332 9320 -292
rect 9290 -352 9320 -332
rect 9380 -332 9430 -292
rect 9380 -352 9410 -332
rect 9490 -392 9550 -132
rect 9150 -402 9230 -392
rect 9150 -462 9160 -402
rect 9220 -412 9230 -402
rect 9470 -402 9550 -392
rect 9470 -412 9480 -402
rect 9220 -462 9480 -412
rect 9540 -462 9550 -402
rect 9150 -472 9550 -462
rect 9606 -52 10006 -42
rect 9606 -112 9616 -52
rect 9676 -102 9936 -52
rect 9676 -112 9686 -102
rect 9606 -122 9686 -112
rect 9926 -112 9936 -102
rect 9996 -112 10006 -52
rect 9926 -122 10006 -112
rect 9606 -392 9666 -122
rect 9936 -132 10006 -122
rect 9746 -182 9776 -162
rect 9726 -222 9776 -182
rect 9836 -182 9866 -162
rect 9836 -222 9886 -182
rect 9726 -292 9886 -222
rect 9726 -332 9776 -292
rect 9746 -352 9776 -332
rect 9836 -332 9886 -292
rect 9836 -352 9866 -332
rect 9946 -392 10006 -132
rect 9606 -402 9686 -392
rect 9606 -462 9616 -402
rect 9676 -412 9686 -402
rect 9926 -402 10006 -392
rect 9926 -412 9936 -402
rect 9676 -462 9936 -412
rect 9996 -462 10006 -402
rect 9606 -472 10006 -462
rect 10062 -52 10462 -42
rect 10062 -112 10072 -52
rect 10132 -102 10392 -52
rect 10132 -112 10142 -102
rect 10062 -122 10142 -112
rect 10382 -112 10392 -102
rect 10452 -112 10462 -52
rect 10382 -122 10462 -112
rect 10062 -392 10122 -122
rect 10392 -132 10462 -122
rect 10202 -182 10232 -162
rect 10182 -222 10232 -182
rect 10292 -182 10322 -162
rect 10292 -222 10342 -182
rect 10182 -292 10342 -222
rect 10182 -332 10232 -292
rect 10202 -352 10232 -332
rect 10292 -332 10342 -292
rect 10292 -352 10322 -332
rect 10402 -392 10462 -132
rect 10062 -402 10142 -392
rect 10062 -462 10072 -402
rect 10132 -412 10142 -402
rect 10382 -402 10462 -392
rect 10382 -412 10392 -402
rect 10132 -462 10392 -412
rect 10452 -462 10462 -402
rect 10062 -472 10462 -462
rect 10520 -52 10920 -42
rect 10520 -112 10530 -52
rect 10590 -102 10850 -52
rect 10590 -112 10600 -102
rect 10520 -122 10600 -112
rect 10840 -112 10850 -102
rect 10910 -112 10920 -52
rect 10840 -122 10920 -112
rect 10520 -392 10580 -122
rect 10850 -132 10920 -122
rect 10660 -182 10690 -162
rect 10640 -222 10690 -182
rect 10750 -182 10780 -162
rect 10750 -222 10800 -182
rect 10640 -292 10800 -222
rect 10640 -332 10690 -292
rect 10660 -352 10690 -332
rect 10750 -332 10800 -292
rect 10750 -352 10780 -332
rect 10860 -392 10920 -132
rect 10520 -402 10600 -392
rect 10520 -462 10530 -402
rect 10590 -412 10600 -402
rect 10840 -402 10920 -392
rect 10840 -412 10850 -402
rect 10590 -462 10850 -412
rect 10910 -462 10920 -402
rect 10520 -472 10920 -462
rect 10976 -52 11376 -42
rect 10976 -112 10986 -52
rect 11046 -102 11306 -52
rect 11046 -112 11056 -102
rect 10976 -122 11056 -112
rect 11296 -112 11306 -102
rect 11366 -112 11376 -52
rect 11296 -122 11376 -112
rect 10976 -392 11036 -122
rect 11306 -132 11376 -122
rect 11116 -182 11146 -162
rect 11096 -222 11146 -182
rect 11206 -182 11236 -162
rect 11206 -222 11256 -182
rect 11096 -292 11256 -222
rect 11096 -332 11146 -292
rect 11116 -352 11146 -332
rect 11206 -332 11256 -292
rect 11206 -352 11236 -332
rect 11316 -392 11376 -132
rect 10976 -402 11056 -392
rect 10976 -462 10986 -402
rect 11046 -412 11056 -402
rect 11296 -402 11376 -392
rect 11296 -412 11306 -402
rect 11046 -462 11306 -412
rect 11366 -462 11376 -402
rect 10976 -472 11376 -462
rect 11432 -52 11832 -42
rect 11432 -112 11442 -52
rect 11502 -102 11762 -52
rect 11502 -112 11512 -102
rect 11432 -122 11512 -112
rect 11752 -112 11762 -102
rect 11822 -112 11832 -52
rect 11752 -122 11832 -112
rect 11432 -392 11492 -122
rect 11762 -132 11832 -122
rect 11572 -182 11602 -162
rect 11552 -222 11602 -182
rect 11662 -182 11692 -162
rect 11662 -222 11712 -182
rect 11552 -292 11712 -222
rect 11552 -332 11602 -292
rect 11572 -352 11602 -332
rect 11662 -332 11712 -292
rect 11662 -352 11692 -332
rect 11772 -392 11832 -132
rect 11432 -402 11512 -392
rect 11432 -462 11442 -402
rect 11502 -412 11512 -402
rect 11752 -402 11832 -392
rect 11752 -412 11762 -402
rect 11502 -462 11762 -412
rect 11822 -462 11832 -402
rect 11432 -472 11832 -462
rect 11890 -52 12290 -42
rect 11890 -112 11900 -52
rect 11960 -102 12220 -52
rect 11960 -112 11970 -102
rect 11890 -122 11970 -112
rect 12210 -112 12220 -102
rect 12280 -112 12290 -52
rect 12210 -122 12290 -112
rect 11890 -392 11950 -122
rect 12220 -132 12290 -122
rect 12030 -182 12060 -162
rect 12010 -222 12060 -182
rect 12120 -182 12150 -162
rect 12120 -222 12170 -182
rect 12010 -292 12170 -222
rect 12010 -332 12060 -292
rect 12030 -352 12060 -332
rect 12120 -332 12170 -292
rect 12120 -352 12150 -332
rect 12230 -392 12290 -132
rect 11890 -402 11970 -392
rect 11890 -462 11900 -402
rect 11960 -412 11970 -402
rect 12210 -402 12290 -392
rect 12210 -412 12220 -402
rect 11960 -462 12220 -412
rect 12280 -462 12290 -402
rect 11890 -472 12290 -462
rect 12346 -52 12746 -42
rect 12346 -112 12356 -52
rect 12416 -102 12676 -52
rect 12416 -112 12426 -102
rect 12346 -122 12426 -112
rect 12666 -112 12676 -102
rect 12736 -112 12746 -52
rect 12666 -122 12746 -112
rect 12346 -392 12406 -122
rect 12676 -132 12746 -122
rect 12486 -182 12516 -162
rect 12466 -222 12516 -182
rect 12576 -182 12606 -162
rect 12576 -222 12626 -182
rect 12466 -292 12626 -222
rect 12466 -332 12516 -292
rect 12486 -352 12516 -332
rect 12576 -332 12626 -292
rect 12576 -352 12606 -332
rect 12686 -392 12746 -132
rect 12346 -402 12426 -392
rect 12346 -462 12356 -402
rect 12416 -412 12426 -402
rect 12666 -402 12746 -392
rect 12666 -412 12676 -402
rect 12416 -462 12676 -412
rect 12736 -462 12746 -402
rect 12346 -472 12746 -462
rect 12802 -52 13202 -42
rect 12802 -112 12812 -52
rect 12872 -102 13132 -52
rect 12872 -112 12882 -102
rect 12802 -122 12882 -112
rect 13122 -112 13132 -102
rect 13192 -112 13202 -52
rect 13122 -122 13202 -112
rect 12802 -392 12862 -122
rect 13132 -132 13202 -122
rect 12942 -182 12972 -162
rect 12922 -222 12972 -182
rect 13032 -182 13062 -162
rect 13032 -222 13082 -182
rect 12922 -292 13082 -222
rect 12922 -332 12972 -292
rect 12942 -352 12972 -332
rect 13032 -332 13082 -292
rect 13032 -352 13062 -332
rect 13142 -392 13202 -132
rect 12802 -402 12882 -392
rect 12802 -462 12812 -402
rect 12872 -412 12882 -402
rect 13122 -402 13202 -392
rect 13122 -412 13132 -402
rect 12872 -462 13132 -412
rect 13192 -462 13202 -402
rect 12802 -472 13202 -462
rect 13260 -52 13660 -42
rect 13260 -112 13270 -52
rect 13330 -102 13590 -52
rect 13330 -112 13340 -102
rect 13260 -122 13340 -112
rect 13580 -112 13590 -102
rect 13650 -112 13660 -52
rect 13580 -122 13660 -112
rect 13260 -392 13320 -122
rect 13590 -132 13660 -122
rect 13400 -182 13430 -162
rect 13380 -222 13430 -182
rect 13490 -182 13520 -162
rect 13490 -222 13540 -182
rect 13380 -292 13540 -222
rect 13380 -332 13430 -292
rect 13400 -352 13430 -332
rect 13490 -332 13540 -292
rect 13490 -352 13520 -332
rect 13600 -392 13660 -132
rect 13260 -402 13340 -392
rect 13260 -462 13270 -402
rect 13330 -412 13340 -402
rect 13580 -402 13660 -392
rect 13580 -412 13590 -402
rect 13330 -462 13590 -412
rect 13650 -462 13660 -402
rect 13260 -472 13660 -462
rect 13716 -52 14116 -42
rect 13716 -112 13726 -52
rect 13786 -102 14046 -52
rect 13786 -112 13796 -102
rect 13716 -122 13796 -112
rect 14036 -112 14046 -102
rect 14106 -112 14116 -52
rect 14036 -122 14116 -112
rect 13716 -392 13776 -122
rect 14046 -132 14116 -122
rect 13856 -182 13886 -162
rect 13836 -222 13886 -182
rect 13946 -182 13976 -162
rect 13946 -222 13996 -182
rect 13836 -292 13996 -222
rect 13836 -332 13886 -292
rect 13856 -352 13886 -332
rect 13946 -332 13996 -292
rect 13946 -352 13976 -332
rect 14056 -392 14116 -132
rect 13716 -402 13796 -392
rect 13716 -462 13726 -402
rect 13786 -412 13796 -402
rect 14036 -402 14116 -392
rect 14036 -412 14046 -402
rect 13786 -462 14046 -412
rect 14106 -462 14116 -402
rect 13716 -472 14116 -462
rect 14172 -52 14572 -42
rect 14172 -112 14182 -52
rect 14242 -102 14502 -52
rect 14242 -112 14252 -102
rect 14172 -122 14252 -112
rect 14492 -112 14502 -102
rect 14562 -112 14572 -52
rect 14492 -122 14572 -112
rect 14172 -392 14232 -122
rect 14502 -132 14572 -122
rect 14312 -182 14342 -162
rect 14292 -222 14342 -182
rect 14402 -182 14432 -162
rect 14402 -222 14452 -182
rect 14292 -292 14452 -222
rect 14292 -332 14342 -292
rect 14312 -352 14342 -332
rect 14402 -332 14452 -292
rect 14402 -352 14432 -332
rect 14512 -392 14572 -132
rect 14172 -402 14252 -392
rect 14172 -462 14182 -402
rect 14242 -412 14252 -402
rect 14492 -402 14572 -392
rect 14492 -412 14502 -402
rect 14242 -462 14502 -412
rect 14562 -462 14572 -402
rect 14172 -472 14572 -462
rect 14630 -52 15030 -42
rect 14630 -112 14640 -52
rect 14700 -102 14960 -52
rect 14700 -112 14710 -102
rect 14630 -122 14710 -112
rect 14950 -112 14960 -102
rect 15020 -112 15030 -52
rect 14950 -122 15030 -112
rect 14630 -392 14690 -122
rect 14960 -132 15030 -122
rect 14770 -182 14800 -162
rect 14750 -222 14800 -182
rect 14860 -182 14890 -162
rect 14860 -222 14910 -182
rect 14750 -292 14910 -222
rect 14750 -332 14800 -292
rect 14770 -352 14800 -332
rect 14860 -332 14910 -292
rect 14860 -352 14890 -332
rect 14970 -392 15030 -132
rect 14630 -402 14710 -392
rect 14630 -462 14640 -402
rect 14700 -412 14710 -402
rect 14950 -402 15030 -392
rect 14950 -412 14960 -402
rect 14700 -462 14960 -412
rect 15020 -462 15030 -402
rect 14630 -472 15030 -462
rect 15086 -52 15486 -42
rect 15086 -112 15096 -52
rect 15156 -102 15416 -52
rect 15156 -112 15166 -102
rect 15086 -122 15166 -112
rect 15406 -112 15416 -102
rect 15476 -112 15486 -52
rect 15406 -122 15486 -112
rect 15086 -392 15146 -122
rect 15416 -132 15486 -122
rect 15226 -182 15256 -162
rect 15206 -222 15256 -182
rect 15316 -182 15346 -162
rect 15316 -222 15366 -182
rect 15206 -292 15366 -222
rect 15206 -332 15256 -292
rect 15226 -352 15256 -332
rect 15316 -332 15366 -292
rect 15316 -352 15346 -332
rect 15426 -392 15486 -132
rect 15086 -402 15166 -392
rect 15086 -462 15096 -402
rect 15156 -412 15166 -402
rect 15406 -402 15486 -392
rect 15406 -412 15416 -402
rect 15156 -462 15416 -412
rect 15476 -462 15486 -402
rect 15086 -472 15486 -462
rect 0 -554 400 -544
rect 0 -614 10 -554
rect 70 -604 330 -554
rect 70 -614 80 -604
rect 0 -624 80 -614
rect 320 -614 330 -604
rect 390 -614 400 -554
rect 320 -624 400 -614
rect 0 -894 60 -624
rect 330 -634 400 -624
rect 140 -684 170 -664
rect 120 -724 170 -684
rect 230 -684 260 -664
rect 230 -724 280 -684
rect 120 -794 280 -724
rect 120 -834 170 -794
rect 140 -854 170 -834
rect 230 -834 280 -794
rect 230 -854 260 -834
rect 340 -894 400 -634
rect 0 -904 80 -894
rect 0 -964 10 -904
rect 70 -914 80 -904
rect 320 -904 400 -894
rect 320 -914 330 -904
rect 70 -964 330 -914
rect 390 -964 400 -904
rect 0 -974 400 -964
rect 456 -554 856 -544
rect 456 -614 466 -554
rect 526 -604 786 -554
rect 526 -614 536 -604
rect 456 -624 536 -614
rect 776 -614 786 -604
rect 846 -614 856 -554
rect 776 -624 856 -614
rect 456 -894 516 -624
rect 786 -634 856 -624
rect 596 -684 626 -664
rect 576 -724 626 -684
rect 686 -684 716 -664
rect 686 -724 736 -684
rect 576 -794 736 -724
rect 576 -834 626 -794
rect 596 -854 626 -834
rect 686 -834 736 -794
rect 686 -854 716 -834
rect 796 -894 856 -634
rect 456 -904 536 -894
rect 456 -964 466 -904
rect 526 -914 536 -904
rect 776 -904 856 -894
rect 776 -914 786 -904
rect 526 -964 786 -914
rect 846 -964 856 -904
rect 456 -974 856 -964
rect 912 -554 1312 -544
rect 912 -614 922 -554
rect 982 -604 1242 -554
rect 982 -614 992 -604
rect 912 -624 992 -614
rect 1232 -614 1242 -604
rect 1302 -614 1312 -554
rect 1232 -624 1312 -614
rect 912 -894 972 -624
rect 1242 -634 1312 -624
rect 1052 -684 1082 -664
rect 1032 -724 1082 -684
rect 1142 -684 1172 -664
rect 1142 -724 1192 -684
rect 1032 -794 1192 -724
rect 1032 -834 1082 -794
rect 1052 -854 1082 -834
rect 1142 -834 1192 -794
rect 1142 -854 1172 -834
rect 1252 -894 1312 -634
rect 912 -904 992 -894
rect 912 -964 922 -904
rect 982 -914 992 -904
rect 1232 -904 1312 -894
rect 1232 -914 1242 -904
rect 982 -964 1242 -914
rect 1302 -964 1312 -904
rect 912 -974 1312 -964
rect 1370 -554 1770 -544
rect 1370 -614 1380 -554
rect 1440 -604 1700 -554
rect 1440 -614 1450 -604
rect 1370 -624 1450 -614
rect 1690 -614 1700 -604
rect 1760 -614 1770 -554
rect 1690 -624 1770 -614
rect 1370 -894 1430 -624
rect 1700 -634 1770 -624
rect 1510 -684 1540 -664
rect 1490 -724 1540 -684
rect 1600 -684 1630 -664
rect 1600 -724 1650 -684
rect 1490 -794 1650 -724
rect 1490 -834 1540 -794
rect 1510 -854 1540 -834
rect 1600 -834 1650 -794
rect 1600 -854 1630 -834
rect 1710 -894 1770 -634
rect 1370 -904 1450 -894
rect 1370 -964 1380 -904
rect 1440 -914 1450 -904
rect 1690 -904 1770 -894
rect 1690 -914 1700 -904
rect 1440 -964 1700 -914
rect 1760 -964 1770 -904
rect 1370 -974 1770 -964
rect 1826 -554 2226 -544
rect 1826 -614 1836 -554
rect 1896 -604 2156 -554
rect 1896 -614 1906 -604
rect 1826 -624 1906 -614
rect 2146 -614 2156 -604
rect 2216 -614 2226 -554
rect 2146 -624 2226 -614
rect 1826 -894 1886 -624
rect 2156 -634 2226 -624
rect 1966 -684 1996 -664
rect 1946 -724 1996 -684
rect 2056 -684 2086 -664
rect 2056 -724 2106 -684
rect 1946 -794 2106 -724
rect 1946 -834 1996 -794
rect 1966 -854 1996 -834
rect 2056 -834 2106 -794
rect 2056 -854 2086 -834
rect 2166 -894 2226 -634
rect 1826 -904 1906 -894
rect 1826 -964 1836 -904
rect 1896 -914 1906 -904
rect 2146 -904 2226 -894
rect 2146 -914 2156 -904
rect 1896 -964 2156 -914
rect 2216 -964 2226 -904
rect 1826 -974 2226 -964
rect 2282 -554 2682 -544
rect 2282 -614 2292 -554
rect 2352 -604 2612 -554
rect 2352 -614 2362 -604
rect 2282 -624 2362 -614
rect 2602 -614 2612 -604
rect 2672 -614 2682 -554
rect 2602 -624 2682 -614
rect 2282 -894 2342 -624
rect 2612 -634 2682 -624
rect 2422 -684 2452 -664
rect 2402 -724 2452 -684
rect 2512 -684 2542 -664
rect 2512 -724 2562 -684
rect 2402 -794 2562 -724
rect 2402 -834 2452 -794
rect 2422 -854 2452 -834
rect 2512 -834 2562 -794
rect 2512 -854 2542 -834
rect 2622 -894 2682 -634
rect 2282 -904 2362 -894
rect 2282 -964 2292 -904
rect 2352 -914 2362 -904
rect 2602 -904 2682 -894
rect 2602 -914 2612 -904
rect 2352 -964 2612 -914
rect 2672 -964 2682 -904
rect 2282 -974 2682 -964
rect 2740 -554 3140 -544
rect 2740 -614 2750 -554
rect 2810 -604 3070 -554
rect 2810 -614 2820 -604
rect 2740 -624 2820 -614
rect 3060 -614 3070 -604
rect 3130 -614 3140 -554
rect 3060 -624 3140 -614
rect 2740 -894 2800 -624
rect 3070 -634 3140 -624
rect 2880 -684 2910 -664
rect 2860 -724 2910 -684
rect 2970 -684 3000 -664
rect 2970 -724 3020 -684
rect 2860 -794 3020 -724
rect 2860 -834 2910 -794
rect 2880 -854 2910 -834
rect 2970 -834 3020 -794
rect 2970 -854 3000 -834
rect 3080 -894 3140 -634
rect 2740 -904 2820 -894
rect 2740 -964 2750 -904
rect 2810 -914 2820 -904
rect 3060 -904 3140 -894
rect 3060 -914 3070 -904
rect 2810 -964 3070 -914
rect 3130 -964 3140 -904
rect 2740 -974 3140 -964
rect 3196 -554 3596 -544
rect 3196 -614 3206 -554
rect 3266 -604 3526 -554
rect 3266 -614 3276 -604
rect 3196 -624 3276 -614
rect 3516 -614 3526 -604
rect 3586 -614 3596 -554
rect 3516 -624 3596 -614
rect 3196 -894 3256 -624
rect 3526 -634 3596 -624
rect 3336 -684 3366 -664
rect 3316 -724 3366 -684
rect 3426 -684 3456 -664
rect 3426 -724 3476 -684
rect 3316 -794 3476 -724
rect 3316 -834 3366 -794
rect 3336 -854 3366 -834
rect 3426 -834 3476 -794
rect 3426 -854 3456 -834
rect 3536 -894 3596 -634
rect 3196 -904 3276 -894
rect 3196 -964 3206 -904
rect 3266 -914 3276 -904
rect 3516 -904 3596 -894
rect 3516 -914 3526 -904
rect 3266 -964 3526 -914
rect 3586 -964 3596 -904
rect 3196 -974 3596 -964
rect 3652 -554 4052 -544
rect 3652 -614 3662 -554
rect 3722 -604 3982 -554
rect 3722 -614 3732 -604
rect 3652 -624 3732 -614
rect 3972 -614 3982 -604
rect 4042 -614 4052 -554
rect 3972 -624 4052 -614
rect 3652 -894 3712 -624
rect 3982 -634 4052 -624
rect 3792 -684 3822 -664
rect 3772 -724 3822 -684
rect 3882 -684 3912 -664
rect 3882 -724 3932 -684
rect 3772 -794 3932 -724
rect 3772 -834 3822 -794
rect 3792 -854 3822 -834
rect 3882 -834 3932 -794
rect 3882 -854 3912 -834
rect 3992 -894 4052 -634
rect 3652 -904 3732 -894
rect 3652 -964 3662 -904
rect 3722 -914 3732 -904
rect 3972 -904 4052 -894
rect 3972 -914 3982 -904
rect 3722 -964 3982 -914
rect 4042 -964 4052 -904
rect 3652 -974 4052 -964
rect 4110 -554 4510 -544
rect 4110 -614 4120 -554
rect 4180 -604 4440 -554
rect 4180 -614 4190 -604
rect 4110 -624 4190 -614
rect 4430 -614 4440 -604
rect 4500 -614 4510 -554
rect 4430 -624 4510 -614
rect 4110 -894 4170 -624
rect 4440 -634 4510 -624
rect 4250 -684 4280 -664
rect 4230 -724 4280 -684
rect 4340 -684 4370 -664
rect 4340 -724 4390 -684
rect 4230 -794 4390 -724
rect 4230 -834 4280 -794
rect 4250 -854 4280 -834
rect 4340 -834 4390 -794
rect 4340 -854 4370 -834
rect 4450 -894 4510 -634
rect 4110 -904 4190 -894
rect 4110 -964 4120 -904
rect 4180 -914 4190 -904
rect 4430 -904 4510 -894
rect 4430 -914 4440 -904
rect 4180 -964 4440 -914
rect 4500 -964 4510 -904
rect 4110 -974 4510 -964
rect 4566 -554 4966 -544
rect 4566 -614 4576 -554
rect 4636 -604 4896 -554
rect 4636 -614 4646 -604
rect 4566 -624 4646 -614
rect 4886 -614 4896 -604
rect 4956 -614 4966 -554
rect 4886 -624 4966 -614
rect 4566 -894 4626 -624
rect 4896 -634 4966 -624
rect 4706 -684 4736 -664
rect 4686 -724 4736 -684
rect 4796 -684 4826 -664
rect 4796 -724 4846 -684
rect 4686 -794 4846 -724
rect 4686 -834 4736 -794
rect 4706 -854 4736 -834
rect 4796 -834 4846 -794
rect 4796 -854 4826 -834
rect 4906 -894 4966 -634
rect 4566 -904 4646 -894
rect 4566 -964 4576 -904
rect 4636 -914 4646 -904
rect 4886 -904 4966 -894
rect 4886 -914 4896 -904
rect 4636 -964 4896 -914
rect 4956 -964 4966 -904
rect 4566 -974 4966 -964
rect 5022 -554 5422 -544
rect 5022 -614 5032 -554
rect 5092 -604 5352 -554
rect 5092 -614 5102 -604
rect 5022 -624 5102 -614
rect 5342 -614 5352 -604
rect 5412 -614 5422 -554
rect 5342 -624 5422 -614
rect 5022 -894 5082 -624
rect 5352 -634 5422 -624
rect 5162 -684 5192 -664
rect 5142 -724 5192 -684
rect 5252 -684 5282 -664
rect 5252 -724 5302 -684
rect 5142 -794 5302 -724
rect 5142 -834 5192 -794
rect 5162 -854 5192 -834
rect 5252 -834 5302 -794
rect 5252 -854 5282 -834
rect 5362 -894 5422 -634
rect 5022 -904 5102 -894
rect 5022 -964 5032 -904
rect 5092 -914 5102 -904
rect 5342 -904 5422 -894
rect 5342 -914 5352 -904
rect 5092 -964 5352 -914
rect 5412 -964 5422 -904
rect 5022 -974 5422 -964
rect 5480 -554 5880 -544
rect 5480 -614 5490 -554
rect 5550 -604 5810 -554
rect 5550 -614 5560 -604
rect 5480 -624 5560 -614
rect 5800 -614 5810 -604
rect 5870 -614 5880 -554
rect 5800 -624 5880 -614
rect 5480 -894 5540 -624
rect 5810 -634 5880 -624
rect 5620 -684 5650 -664
rect 5600 -724 5650 -684
rect 5710 -684 5740 -664
rect 5710 -724 5760 -684
rect 5600 -794 5760 -724
rect 5600 -834 5650 -794
rect 5620 -854 5650 -834
rect 5710 -834 5760 -794
rect 5710 -854 5740 -834
rect 5820 -894 5880 -634
rect 5480 -904 5560 -894
rect 5480 -964 5490 -904
rect 5550 -914 5560 -904
rect 5800 -904 5880 -894
rect 5800 -914 5810 -904
rect 5550 -964 5810 -914
rect 5870 -964 5880 -904
rect 5480 -974 5880 -964
rect 5936 -554 6336 -544
rect 5936 -614 5946 -554
rect 6006 -604 6266 -554
rect 6006 -614 6016 -604
rect 5936 -624 6016 -614
rect 6256 -614 6266 -604
rect 6326 -614 6336 -554
rect 6256 -624 6336 -614
rect 5936 -894 5996 -624
rect 6266 -634 6336 -624
rect 6076 -684 6106 -664
rect 6056 -724 6106 -684
rect 6166 -684 6196 -664
rect 6166 -724 6216 -684
rect 6056 -794 6216 -724
rect 6056 -834 6106 -794
rect 6076 -854 6106 -834
rect 6166 -834 6216 -794
rect 6166 -854 6196 -834
rect 6276 -894 6336 -634
rect 5936 -904 6016 -894
rect 5936 -964 5946 -904
rect 6006 -914 6016 -904
rect 6256 -904 6336 -894
rect 6256 -914 6266 -904
rect 6006 -964 6266 -914
rect 6326 -964 6336 -904
rect 5936 -974 6336 -964
rect 6392 -554 6792 -544
rect 6392 -614 6402 -554
rect 6462 -604 6722 -554
rect 6462 -614 6472 -604
rect 6392 -624 6472 -614
rect 6712 -614 6722 -604
rect 6782 -614 6792 -554
rect 6712 -624 6792 -614
rect 6392 -894 6452 -624
rect 6722 -634 6792 -624
rect 6532 -684 6562 -664
rect 6512 -724 6562 -684
rect 6622 -684 6652 -664
rect 6622 -724 6672 -684
rect 6512 -794 6672 -724
rect 6512 -834 6562 -794
rect 6532 -854 6562 -834
rect 6622 -834 6672 -794
rect 6622 -854 6652 -834
rect 6732 -894 6792 -634
rect 6392 -904 6472 -894
rect 6392 -964 6402 -904
rect 6462 -914 6472 -904
rect 6712 -904 6792 -894
rect 6712 -914 6722 -904
rect 6462 -964 6722 -914
rect 6782 -964 6792 -904
rect 6392 -974 6792 -964
rect 6850 -554 7250 -544
rect 6850 -614 6860 -554
rect 6920 -604 7180 -554
rect 6920 -614 6930 -604
rect 6850 -624 6930 -614
rect 7170 -614 7180 -604
rect 7240 -614 7250 -554
rect 7170 -624 7250 -614
rect 6850 -894 6910 -624
rect 7180 -634 7250 -624
rect 6990 -684 7020 -664
rect 6970 -724 7020 -684
rect 7080 -684 7110 -664
rect 7080 -724 7130 -684
rect 6970 -794 7130 -724
rect 6970 -834 7020 -794
rect 6990 -854 7020 -834
rect 7080 -834 7130 -794
rect 7080 -854 7110 -834
rect 7190 -894 7250 -634
rect 6850 -904 6930 -894
rect 6850 -964 6860 -904
rect 6920 -914 6930 -904
rect 7170 -904 7250 -894
rect 7170 -914 7180 -904
rect 6920 -964 7180 -914
rect 7240 -964 7250 -904
rect 6850 -974 7250 -964
rect 7306 -554 7706 -544
rect 7306 -614 7316 -554
rect 7376 -604 7636 -554
rect 7376 -614 7386 -604
rect 7306 -624 7386 -614
rect 7626 -614 7636 -604
rect 7696 -614 7706 -554
rect 7626 -624 7706 -614
rect 7306 -894 7366 -624
rect 7636 -634 7706 -624
rect 7446 -684 7476 -664
rect 7426 -724 7476 -684
rect 7536 -684 7566 -664
rect 7536 -724 7586 -684
rect 7426 -794 7586 -724
rect 7426 -834 7476 -794
rect 7446 -854 7476 -834
rect 7536 -834 7586 -794
rect 7536 -854 7566 -834
rect 7646 -894 7706 -634
rect 7306 -904 7386 -894
rect 7306 -964 7316 -904
rect 7376 -914 7386 -904
rect 7626 -904 7706 -894
rect 7626 -914 7636 -904
rect 7376 -964 7636 -914
rect 7696 -964 7706 -904
rect 7306 -974 7706 -964
rect 7762 -554 8162 -544
rect 7762 -614 7772 -554
rect 7832 -604 8092 -554
rect 7832 -614 7842 -604
rect 7762 -624 7842 -614
rect 8082 -614 8092 -604
rect 8152 -614 8162 -554
rect 8082 -624 8162 -614
rect 7762 -894 7822 -624
rect 8092 -634 8162 -624
rect 7902 -684 7932 -664
rect 7882 -724 7932 -684
rect 7992 -684 8022 -664
rect 7992 -724 8042 -684
rect 7882 -794 8042 -724
rect 7882 -834 7932 -794
rect 7902 -854 7932 -834
rect 7992 -834 8042 -794
rect 7992 -854 8022 -834
rect 8102 -894 8162 -634
rect 7762 -904 7842 -894
rect 7762 -964 7772 -904
rect 7832 -914 7842 -904
rect 8082 -904 8162 -894
rect 8082 -914 8092 -904
rect 7832 -964 8092 -914
rect 8152 -964 8162 -904
rect 7762 -974 8162 -964
rect 8236 -554 8636 -544
rect 8236 -614 8246 -554
rect 8306 -604 8566 -554
rect 8306 -614 8316 -604
rect 8236 -624 8316 -614
rect 8556 -614 8566 -604
rect 8626 -614 8636 -554
rect 8556 -624 8636 -614
rect 8236 -894 8296 -624
rect 8566 -634 8636 -624
rect 8376 -684 8406 -664
rect 8356 -724 8406 -684
rect 8466 -684 8496 -664
rect 8466 -724 8516 -684
rect 8356 -794 8516 -724
rect 8356 -834 8406 -794
rect 8376 -854 8406 -834
rect 8466 -834 8516 -794
rect 8466 -854 8496 -834
rect 8576 -894 8636 -634
rect 8236 -904 8316 -894
rect 8236 -964 8246 -904
rect 8306 -914 8316 -904
rect 8556 -904 8636 -894
rect 8556 -914 8566 -904
rect 8306 -964 8566 -914
rect 8626 -964 8636 -904
rect 8236 -974 8636 -964
rect 8692 -554 9092 -544
rect 8692 -614 8702 -554
rect 8762 -604 9022 -554
rect 8762 -614 8772 -604
rect 8692 -624 8772 -614
rect 9012 -614 9022 -604
rect 9082 -614 9092 -554
rect 9012 -624 9092 -614
rect 8692 -894 8752 -624
rect 9022 -634 9092 -624
rect 8832 -684 8862 -664
rect 8812 -724 8862 -684
rect 8922 -684 8952 -664
rect 8922 -724 8972 -684
rect 8812 -794 8972 -724
rect 8812 -834 8862 -794
rect 8832 -854 8862 -834
rect 8922 -834 8972 -794
rect 8922 -854 8952 -834
rect 9032 -894 9092 -634
rect 8692 -904 8772 -894
rect 8692 -964 8702 -904
rect 8762 -914 8772 -904
rect 9012 -904 9092 -894
rect 9012 -914 9022 -904
rect 8762 -964 9022 -914
rect 9082 -964 9092 -904
rect 8692 -974 9092 -964
rect 9150 -554 9550 -544
rect 9150 -614 9160 -554
rect 9220 -604 9480 -554
rect 9220 -614 9230 -604
rect 9150 -624 9230 -614
rect 9470 -614 9480 -604
rect 9540 -614 9550 -554
rect 9470 -624 9550 -614
rect 9150 -894 9210 -624
rect 9480 -634 9550 -624
rect 9290 -684 9320 -664
rect 9270 -724 9320 -684
rect 9380 -684 9410 -664
rect 9380 -724 9430 -684
rect 9270 -794 9430 -724
rect 9270 -834 9320 -794
rect 9290 -854 9320 -834
rect 9380 -834 9430 -794
rect 9380 -854 9410 -834
rect 9490 -894 9550 -634
rect 9150 -904 9230 -894
rect 9150 -964 9160 -904
rect 9220 -914 9230 -904
rect 9470 -904 9550 -894
rect 9470 -914 9480 -904
rect 9220 -964 9480 -914
rect 9540 -964 9550 -904
rect 9150 -974 9550 -964
rect 9606 -554 10006 -544
rect 9606 -614 9616 -554
rect 9676 -604 9936 -554
rect 9676 -614 9686 -604
rect 9606 -624 9686 -614
rect 9926 -614 9936 -604
rect 9996 -614 10006 -554
rect 9926 -624 10006 -614
rect 9606 -894 9666 -624
rect 9936 -634 10006 -624
rect 9746 -684 9776 -664
rect 9726 -724 9776 -684
rect 9836 -684 9866 -664
rect 9836 -724 9886 -684
rect 9726 -794 9886 -724
rect 9726 -834 9776 -794
rect 9746 -854 9776 -834
rect 9836 -834 9886 -794
rect 9836 -854 9866 -834
rect 9946 -894 10006 -634
rect 9606 -904 9686 -894
rect 9606 -964 9616 -904
rect 9676 -914 9686 -904
rect 9926 -904 10006 -894
rect 9926 -914 9936 -904
rect 9676 -964 9936 -914
rect 9996 -964 10006 -904
rect 9606 -974 10006 -964
rect 10062 -554 10462 -544
rect 10062 -614 10072 -554
rect 10132 -604 10392 -554
rect 10132 -614 10142 -604
rect 10062 -624 10142 -614
rect 10382 -614 10392 -604
rect 10452 -614 10462 -554
rect 10382 -624 10462 -614
rect 10062 -894 10122 -624
rect 10392 -634 10462 -624
rect 10202 -684 10232 -664
rect 10182 -724 10232 -684
rect 10292 -684 10322 -664
rect 10292 -724 10342 -684
rect 10182 -794 10342 -724
rect 10182 -834 10232 -794
rect 10202 -854 10232 -834
rect 10292 -834 10342 -794
rect 10292 -854 10322 -834
rect 10402 -894 10462 -634
rect 10062 -904 10142 -894
rect 10062 -964 10072 -904
rect 10132 -914 10142 -904
rect 10382 -904 10462 -894
rect 10382 -914 10392 -904
rect 10132 -964 10392 -914
rect 10452 -964 10462 -904
rect 10062 -974 10462 -964
rect 10520 -554 10920 -544
rect 10520 -614 10530 -554
rect 10590 -604 10850 -554
rect 10590 -614 10600 -604
rect 10520 -624 10600 -614
rect 10840 -614 10850 -604
rect 10910 -614 10920 -554
rect 10840 -624 10920 -614
rect 10520 -894 10580 -624
rect 10850 -634 10920 -624
rect 10660 -684 10690 -664
rect 10640 -724 10690 -684
rect 10750 -684 10780 -664
rect 10750 -724 10800 -684
rect 10640 -794 10800 -724
rect 10640 -834 10690 -794
rect 10660 -854 10690 -834
rect 10750 -834 10800 -794
rect 10750 -854 10780 -834
rect 10860 -894 10920 -634
rect 10520 -904 10600 -894
rect 10520 -964 10530 -904
rect 10590 -914 10600 -904
rect 10840 -904 10920 -894
rect 10840 -914 10850 -904
rect 10590 -964 10850 -914
rect 10910 -964 10920 -904
rect 10520 -974 10920 -964
rect 10976 -554 11376 -544
rect 10976 -614 10986 -554
rect 11046 -604 11306 -554
rect 11046 -614 11056 -604
rect 10976 -624 11056 -614
rect 11296 -614 11306 -604
rect 11366 -614 11376 -554
rect 11296 -624 11376 -614
rect 10976 -894 11036 -624
rect 11306 -634 11376 -624
rect 11116 -684 11146 -664
rect 11096 -724 11146 -684
rect 11206 -684 11236 -664
rect 11206 -724 11256 -684
rect 11096 -794 11256 -724
rect 11096 -834 11146 -794
rect 11116 -854 11146 -834
rect 11206 -834 11256 -794
rect 11206 -854 11236 -834
rect 11316 -894 11376 -634
rect 10976 -904 11056 -894
rect 10976 -964 10986 -904
rect 11046 -914 11056 -904
rect 11296 -904 11376 -894
rect 11296 -914 11306 -904
rect 11046 -964 11306 -914
rect 11366 -964 11376 -904
rect 10976 -974 11376 -964
rect 11432 -554 11832 -544
rect 11432 -614 11442 -554
rect 11502 -604 11762 -554
rect 11502 -614 11512 -604
rect 11432 -624 11512 -614
rect 11752 -614 11762 -604
rect 11822 -614 11832 -554
rect 11752 -624 11832 -614
rect 11432 -894 11492 -624
rect 11762 -634 11832 -624
rect 11572 -684 11602 -664
rect 11552 -724 11602 -684
rect 11662 -684 11692 -664
rect 11662 -724 11712 -684
rect 11552 -794 11712 -724
rect 11552 -834 11602 -794
rect 11572 -854 11602 -834
rect 11662 -834 11712 -794
rect 11662 -854 11692 -834
rect 11772 -894 11832 -634
rect 11432 -904 11512 -894
rect 11432 -964 11442 -904
rect 11502 -914 11512 -904
rect 11752 -904 11832 -894
rect 11752 -914 11762 -904
rect 11502 -964 11762 -914
rect 11822 -964 11832 -904
rect 11432 -974 11832 -964
rect 11890 -554 12290 -544
rect 11890 -614 11900 -554
rect 11960 -604 12220 -554
rect 11960 -614 11970 -604
rect 11890 -624 11970 -614
rect 12210 -614 12220 -604
rect 12280 -614 12290 -554
rect 12210 -624 12290 -614
rect 11890 -894 11950 -624
rect 12220 -634 12290 -624
rect 12030 -684 12060 -664
rect 12010 -724 12060 -684
rect 12120 -684 12150 -664
rect 12120 -724 12170 -684
rect 12010 -794 12170 -724
rect 12010 -834 12060 -794
rect 12030 -854 12060 -834
rect 12120 -834 12170 -794
rect 12120 -854 12150 -834
rect 12230 -894 12290 -634
rect 11890 -904 11970 -894
rect 11890 -964 11900 -904
rect 11960 -914 11970 -904
rect 12210 -904 12290 -894
rect 12210 -914 12220 -904
rect 11960 -964 12220 -914
rect 12280 -964 12290 -904
rect 11890 -974 12290 -964
rect 12346 -554 12746 -544
rect 12346 -614 12356 -554
rect 12416 -604 12676 -554
rect 12416 -614 12426 -604
rect 12346 -624 12426 -614
rect 12666 -614 12676 -604
rect 12736 -614 12746 -554
rect 12666 -624 12746 -614
rect 12346 -894 12406 -624
rect 12676 -634 12746 -624
rect 12486 -684 12516 -664
rect 12466 -724 12516 -684
rect 12576 -684 12606 -664
rect 12576 -724 12626 -684
rect 12466 -794 12626 -724
rect 12466 -834 12516 -794
rect 12486 -854 12516 -834
rect 12576 -834 12626 -794
rect 12576 -854 12606 -834
rect 12686 -894 12746 -634
rect 12346 -904 12426 -894
rect 12346 -964 12356 -904
rect 12416 -914 12426 -904
rect 12666 -904 12746 -894
rect 12666 -914 12676 -904
rect 12416 -964 12676 -914
rect 12736 -964 12746 -904
rect 12346 -974 12746 -964
rect 12802 -554 13202 -544
rect 12802 -614 12812 -554
rect 12872 -604 13132 -554
rect 12872 -614 12882 -604
rect 12802 -624 12882 -614
rect 13122 -614 13132 -604
rect 13192 -614 13202 -554
rect 13122 -624 13202 -614
rect 12802 -894 12862 -624
rect 13132 -634 13202 -624
rect 12942 -684 12972 -664
rect 12922 -724 12972 -684
rect 13032 -684 13062 -664
rect 13032 -724 13082 -684
rect 12922 -794 13082 -724
rect 12922 -834 12972 -794
rect 12942 -854 12972 -834
rect 13032 -834 13082 -794
rect 13032 -854 13062 -834
rect 13142 -894 13202 -634
rect 12802 -904 12882 -894
rect 12802 -964 12812 -904
rect 12872 -914 12882 -904
rect 13122 -904 13202 -894
rect 13122 -914 13132 -904
rect 12872 -964 13132 -914
rect 13192 -964 13202 -904
rect 12802 -974 13202 -964
rect 13260 -554 13660 -544
rect 13260 -614 13270 -554
rect 13330 -604 13590 -554
rect 13330 -614 13340 -604
rect 13260 -624 13340 -614
rect 13580 -614 13590 -604
rect 13650 -614 13660 -554
rect 13580 -624 13660 -614
rect 13260 -894 13320 -624
rect 13590 -634 13660 -624
rect 13400 -684 13430 -664
rect 13380 -724 13430 -684
rect 13490 -684 13520 -664
rect 13490 -724 13540 -684
rect 13380 -794 13540 -724
rect 13380 -834 13430 -794
rect 13400 -854 13430 -834
rect 13490 -834 13540 -794
rect 13490 -854 13520 -834
rect 13600 -894 13660 -634
rect 13260 -904 13340 -894
rect 13260 -964 13270 -904
rect 13330 -914 13340 -904
rect 13580 -904 13660 -894
rect 13580 -914 13590 -904
rect 13330 -964 13590 -914
rect 13650 -964 13660 -904
rect 13260 -974 13660 -964
rect 13716 -554 14116 -544
rect 13716 -614 13726 -554
rect 13786 -604 14046 -554
rect 13786 -614 13796 -604
rect 13716 -624 13796 -614
rect 14036 -614 14046 -604
rect 14106 -614 14116 -554
rect 14036 -624 14116 -614
rect 13716 -894 13776 -624
rect 14046 -634 14116 -624
rect 13856 -684 13886 -664
rect 13836 -724 13886 -684
rect 13946 -684 13976 -664
rect 13946 -724 13996 -684
rect 13836 -794 13996 -724
rect 13836 -834 13886 -794
rect 13856 -854 13886 -834
rect 13946 -834 13996 -794
rect 13946 -854 13976 -834
rect 14056 -894 14116 -634
rect 13716 -904 13796 -894
rect 13716 -964 13726 -904
rect 13786 -914 13796 -904
rect 14036 -904 14116 -894
rect 14036 -914 14046 -904
rect 13786 -964 14046 -914
rect 14106 -964 14116 -904
rect 13716 -974 14116 -964
rect 14172 -554 14572 -544
rect 14172 -614 14182 -554
rect 14242 -604 14502 -554
rect 14242 -614 14252 -604
rect 14172 -624 14252 -614
rect 14492 -614 14502 -604
rect 14562 -614 14572 -554
rect 14492 -624 14572 -614
rect 14172 -894 14232 -624
rect 14502 -634 14572 -624
rect 14312 -684 14342 -664
rect 14292 -724 14342 -684
rect 14402 -684 14432 -664
rect 14402 -724 14452 -684
rect 14292 -794 14452 -724
rect 14292 -834 14342 -794
rect 14312 -854 14342 -834
rect 14402 -834 14452 -794
rect 14402 -854 14432 -834
rect 14512 -894 14572 -634
rect 14172 -904 14252 -894
rect 14172 -964 14182 -904
rect 14242 -914 14252 -904
rect 14492 -904 14572 -894
rect 14492 -914 14502 -904
rect 14242 -964 14502 -914
rect 14562 -964 14572 -904
rect 14172 -974 14572 -964
rect 14630 -554 15030 -544
rect 14630 -614 14640 -554
rect 14700 -604 14960 -554
rect 14700 -614 14710 -604
rect 14630 -624 14710 -614
rect 14950 -614 14960 -604
rect 15020 -614 15030 -554
rect 14950 -624 15030 -614
rect 14630 -894 14690 -624
rect 14960 -634 15030 -624
rect 14770 -684 14800 -664
rect 14750 -724 14800 -684
rect 14860 -684 14890 -664
rect 14860 -724 14910 -684
rect 14750 -794 14910 -724
rect 14750 -834 14800 -794
rect 14770 -854 14800 -834
rect 14860 -834 14910 -794
rect 14860 -854 14890 -834
rect 14970 -894 15030 -634
rect 14630 -904 14710 -894
rect 14630 -964 14640 -904
rect 14700 -914 14710 -904
rect 14950 -904 15030 -894
rect 14950 -914 14960 -904
rect 14700 -964 14960 -914
rect 15020 -964 15030 -904
rect 14630 -974 15030 -964
rect 15086 -554 15486 -544
rect 15086 -614 15096 -554
rect 15156 -604 15416 -554
rect 15156 -614 15166 -604
rect 15086 -624 15166 -614
rect 15406 -614 15416 -604
rect 15476 -614 15486 -554
rect 15406 -624 15486 -614
rect 15086 -894 15146 -624
rect 15416 -634 15486 -624
rect 15226 -684 15256 -664
rect 15206 -724 15256 -684
rect 15316 -684 15346 -664
rect 15316 -724 15366 -684
rect 15206 -794 15366 -724
rect 15206 -834 15256 -794
rect 15226 -854 15256 -834
rect 15316 -834 15366 -794
rect 15316 -854 15346 -834
rect 15426 -894 15486 -634
rect 15086 -904 15166 -894
rect 15086 -964 15096 -904
rect 15156 -914 15166 -904
rect 15406 -904 15486 -894
rect 15406 -914 15416 -904
rect 15156 -964 15416 -914
rect 15476 -964 15486 -904
rect 15086 -974 15486 -964
rect 0 -1046 400 -1036
rect 0 -1106 10 -1046
rect 70 -1096 330 -1046
rect 70 -1106 80 -1096
rect 0 -1116 80 -1106
rect 320 -1106 330 -1096
rect 390 -1106 400 -1046
rect 320 -1116 400 -1106
rect 0 -1386 60 -1116
rect 330 -1126 400 -1116
rect 140 -1176 170 -1156
rect 120 -1216 170 -1176
rect 230 -1176 260 -1156
rect 230 -1216 280 -1176
rect 120 -1286 280 -1216
rect 120 -1326 170 -1286
rect 140 -1346 170 -1326
rect 230 -1326 280 -1286
rect 230 -1346 260 -1326
rect 340 -1386 400 -1126
rect 0 -1396 80 -1386
rect 0 -1456 10 -1396
rect 70 -1406 80 -1396
rect 320 -1396 400 -1386
rect 320 -1406 330 -1396
rect 70 -1456 330 -1406
rect 390 -1456 400 -1396
rect 0 -1466 400 -1456
rect 456 -1046 856 -1036
rect 456 -1106 466 -1046
rect 526 -1096 786 -1046
rect 526 -1106 536 -1096
rect 456 -1116 536 -1106
rect 776 -1106 786 -1096
rect 846 -1106 856 -1046
rect 776 -1116 856 -1106
rect 456 -1386 516 -1116
rect 786 -1126 856 -1116
rect 596 -1176 626 -1156
rect 576 -1216 626 -1176
rect 686 -1176 716 -1156
rect 686 -1216 736 -1176
rect 576 -1286 736 -1216
rect 576 -1326 626 -1286
rect 596 -1346 626 -1326
rect 686 -1326 736 -1286
rect 686 -1346 716 -1326
rect 796 -1386 856 -1126
rect 456 -1396 536 -1386
rect 456 -1456 466 -1396
rect 526 -1406 536 -1396
rect 776 -1396 856 -1386
rect 776 -1406 786 -1396
rect 526 -1456 786 -1406
rect 846 -1456 856 -1396
rect 456 -1466 856 -1456
rect 912 -1046 1312 -1036
rect 912 -1106 922 -1046
rect 982 -1096 1242 -1046
rect 982 -1106 992 -1096
rect 912 -1116 992 -1106
rect 1232 -1106 1242 -1096
rect 1302 -1106 1312 -1046
rect 1232 -1116 1312 -1106
rect 912 -1386 972 -1116
rect 1242 -1126 1312 -1116
rect 1052 -1176 1082 -1156
rect 1032 -1216 1082 -1176
rect 1142 -1176 1172 -1156
rect 1142 -1216 1192 -1176
rect 1032 -1286 1192 -1216
rect 1032 -1326 1082 -1286
rect 1052 -1346 1082 -1326
rect 1142 -1326 1192 -1286
rect 1142 -1346 1172 -1326
rect 1252 -1386 1312 -1126
rect 912 -1396 992 -1386
rect 912 -1456 922 -1396
rect 982 -1406 992 -1396
rect 1232 -1396 1312 -1386
rect 1232 -1406 1242 -1396
rect 982 -1456 1242 -1406
rect 1302 -1456 1312 -1396
rect 912 -1466 1312 -1456
rect 1370 -1046 1770 -1036
rect 1370 -1106 1380 -1046
rect 1440 -1096 1700 -1046
rect 1440 -1106 1450 -1096
rect 1370 -1116 1450 -1106
rect 1690 -1106 1700 -1096
rect 1760 -1106 1770 -1046
rect 1690 -1116 1770 -1106
rect 1370 -1386 1430 -1116
rect 1700 -1126 1770 -1116
rect 1510 -1176 1540 -1156
rect 1490 -1216 1540 -1176
rect 1600 -1176 1630 -1156
rect 1600 -1216 1650 -1176
rect 1490 -1286 1650 -1216
rect 1490 -1326 1540 -1286
rect 1510 -1346 1540 -1326
rect 1600 -1326 1650 -1286
rect 1600 -1346 1630 -1326
rect 1710 -1386 1770 -1126
rect 1370 -1396 1450 -1386
rect 1370 -1456 1380 -1396
rect 1440 -1406 1450 -1396
rect 1690 -1396 1770 -1386
rect 1690 -1406 1700 -1396
rect 1440 -1456 1700 -1406
rect 1760 -1456 1770 -1396
rect 1370 -1466 1770 -1456
rect 1826 -1046 2226 -1036
rect 1826 -1106 1836 -1046
rect 1896 -1096 2156 -1046
rect 1896 -1106 1906 -1096
rect 1826 -1116 1906 -1106
rect 2146 -1106 2156 -1096
rect 2216 -1106 2226 -1046
rect 2146 -1116 2226 -1106
rect 1826 -1386 1886 -1116
rect 2156 -1126 2226 -1116
rect 1966 -1176 1996 -1156
rect 1946 -1216 1996 -1176
rect 2056 -1176 2086 -1156
rect 2056 -1216 2106 -1176
rect 1946 -1286 2106 -1216
rect 1946 -1326 1996 -1286
rect 1966 -1346 1996 -1326
rect 2056 -1326 2106 -1286
rect 2056 -1346 2086 -1326
rect 2166 -1386 2226 -1126
rect 1826 -1396 1906 -1386
rect 1826 -1456 1836 -1396
rect 1896 -1406 1906 -1396
rect 2146 -1396 2226 -1386
rect 2146 -1406 2156 -1396
rect 1896 -1456 2156 -1406
rect 2216 -1456 2226 -1396
rect 1826 -1466 2226 -1456
rect 2282 -1046 2682 -1036
rect 2282 -1106 2292 -1046
rect 2352 -1096 2612 -1046
rect 2352 -1106 2362 -1096
rect 2282 -1116 2362 -1106
rect 2602 -1106 2612 -1096
rect 2672 -1106 2682 -1046
rect 2602 -1116 2682 -1106
rect 2282 -1386 2342 -1116
rect 2612 -1126 2682 -1116
rect 2422 -1176 2452 -1156
rect 2402 -1216 2452 -1176
rect 2512 -1176 2542 -1156
rect 2512 -1216 2562 -1176
rect 2402 -1286 2562 -1216
rect 2402 -1326 2452 -1286
rect 2422 -1346 2452 -1326
rect 2512 -1326 2562 -1286
rect 2512 -1346 2542 -1326
rect 2622 -1386 2682 -1126
rect 2282 -1396 2362 -1386
rect 2282 -1456 2292 -1396
rect 2352 -1406 2362 -1396
rect 2602 -1396 2682 -1386
rect 2602 -1406 2612 -1396
rect 2352 -1456 2612 -1406
rect 2672 -1456 2682 -1396
rect 2282 -1466 2682 -1456
rect 2740 -1046 3140 -1036
rect 2740 -1106 2750 -1046
rect 2810 -1096 3070 -1046
rect 2810 -1106 2820 -1096
rect 2740 -1116 2820 -1106
rect 3060 -1106 3070 -1096
rect 3130 -1106 3140 -1046
rect 3060 -1116 3140 -1106
rect 2740 -1386 2800 -1116
rect 3070 -1126 3140 -1116
rect 2880 -1176 2910 -1156
rect 2860 -1216 2910 -1176
rect 2970 -1176 3000 -1156
rect 2970 -1216 3020 -1176
rect 2860 -1286 3020 -1216
rect 2860 -1326 2910 -1286
rect 2880 -1346 2910 -1326
rect 2970 -1326 3020 -1286
rect 2970 -1346 3000 -1326
rect 3080 -1386 3140 -1126
rect 2740 -1396 2820 -1386
rect 2740 -1456 2750 -1396
rect 2810 -1406 2820 -1396
rect 3060 -1396 3140 -1386
rect 3060 -1406 3070 -1396
rect 2810 -1456 3070 -1406
rect 3130 -1456 3140 -1396
rect 2740 -1466 3140 -1456
rect 3196 -1046 3596 -1036
rect 3196 -1106 3206 -1046
rect 3266 -1096 3526 -1046
rect 3266 -1106 3276 -1096
rect 3196 -1116 3276 -1106
rect 3516 -1106 3526 -1096
rect 3586 -1106 3596 -1046
rect 3516 -1116 3596 -1106
rect 3196 -1386 3256 -1116
rect 3526 -1126 3596 -1116
rect 3336 -1176 3366 -1156
rect 3316 -1216 3366 -1176
rect 3426 -1176 3456 -1156
rect 3426 -1216 3476 -1176
rect 3316 -1286 3476 -1216
rect 3316 -1326 3366 -1286
rect 3336 -1346 3366 -1326
rect 3426 -1326 3476 -1286
rect 3426 -1346 3456 -1326
rect 3536 -1386 3596 -1126
rect 3196 -1396 3276 -1386
rect 3196 -1456 3206 -1396
rect 3266 -1406 3276 -1396
rect 3516 -1396 3596 -1386
rect 3516 -1406 3526 -1396
rect 3266 -1456 3526 -1406
rect 3586 -1456 3596 -1396
rect 3196 -1466 3596 -1456
rect 3652 -1046 4052 -1036
rect 3652 -1106 3662 -1046
rect 3722 -1096 3982 -1046
rect 3722 -1106 3732 -1096
rect 3652 -1116 3732 -1106
rect 3972 -1106 3982 -1096
rect 4042 -1106 4052 -1046
rect 3972 -1116 4052 -1106
rect 3652 -1386 3712 -1116
rect 3982 -1126 4052 -1116
rect 3792 -1176 3822 -1156
rect 3772 -1216 3822 -1176
rect 3882 -1176 3912 -1156
rect 3882 -1216 3932 -1176
rect 3772 -1286 3932 -1216
rect 3772 -1326 3822 -1286
rect 3792 -1346 3822 -1326
rect 3882 -1326 3932 -1286
rect 3882 -1346 3912 -1326
rect 3992 -1386 4052 -1126
rect 3652 -1396 3732 -1386
rect 3652 -1456 3662 -1396
rect 3722 -1406 3732 -1396
rect 3972 -1396 4052 -1386
rect 3972 -1406 3982 -1396
rect 3722 -1456 3982 -1406
rect 4042 -1456 4052 -1396
rect 3652 -1466 4052 -1456
rect 4110 -1046 4510 -1036
rect 4110 -1106 4120 -1046
rect 4180 -1096 4440 -1046
rect 4180 -1106 4190 -1096
rect 4110 -1116 4190 -1106
rect 4430 -1106 4440 -1096
rect 4500 -1106 4510 -1046
rect 4430 -1116 4510 -1106
rect 4110 -1386 4170 -1116
rect 4440 -1126 4510 -1116
rect 4250 -1176 4280 -1156
rect 4230 -1216 4280 -1176
rect 4340 -1176 4370 -1156
rect 4340 -1216 4390 -1176
rect 4230 -1286 4390 -1216
rect 4230 -1326 4280 -1286
rect 4250 -1346 4280 -1326
rect 4340 -1326 4390 -1286
rect 4340 -1346 4370 -1326
rect 4450 -1386 4510 -1126
rect 4110 -1396 4190 -1386
rect 4110 -1456 4120 -1396
rect 4180 -1406 4190 -1396
rect 4430 -1396 4510 -1386
rect 4430 -1406 4440 -1396
rect 4180 -1456 4440 -1406
rect 4500 -1456 4510 -1396
rect 4110 -1466 4510 -1456
rect 4566 -1046 4966 -1036
rect 4566 -1106 4576 -1046
rect 4636 -1096 4896 -1046
rect 4636 -1106 4646 -1096
rect 4566 -1116 4646 -1106
rect 4886 -1106 4896 -1096
rect 4956 -1106 4966 -1046
rect 4886 -1116 4966 -1106
rect 4566 -1386 4626 -1116
rect 4896 -1126 4966 -1116
rect 4706 -1176 4736 -1156
rect 4686 -1216 4736 -1176
rect 4796 -1176 4826 -1156
rect 4796 -1216 4846 -1176
rect 4686 -1286 4846 -1216
rect 4686 -1326 4736 -1286
rect 4706 -1346 4736 -1326
rect 4796 -1326 4846 -1286
rect 4796 -1346 4826 -1326
rect 4906 -1386 4966 -1126
rect 4566 -1396 4646 -1386
rect 4566 -1456 4576 -1396
rect 4636 -1406 4646 -1396
rect 4886 -1396 4966 -1386
rect 4886 -1406 4896 -1396
rect 4636 -1456 4896 -1406
rect 4956 -1456 4966 -1396
rect 4566 -1466 4966 -1456
rect 5022 -1046 5422 -1036
rect 5022 -1106 5032 -1046
rect 5092 -1096 5352 -1046
rect 5092 -1106 5102 -1096
rect 5022 -1116 5102 -1106
rect 5342 -1106 5352 -1096
rect 5412 -1106 5422 -1046
rect 5342 -1116 5422 -1106
rect 5022 -1386 5082 -1116
rect 5352 -1126 5422 -1116
rect 5162 -1176 5192 -1156
rect 5142 -1216 5192 -1176
rect 5252 -1176 5282 -1156
rect 5252 -1216 5302 -1176
rect 5142 -1286 5302 -1216
rect 5142 -1326 5192 -1286
rect 5162 -1346 5192 -1326
rect 5252 -1326 5302 -1286
rect 5252 -1346 5282 -1326
rect 5362 -1386 5422 -1126
rect 5022 -1396 5102 -1386
rect 5022 -1456 5032 -1396
rect 5092 -1406 5102 -1396
rect 5342 -1396 5422 -1386
rect 5342 -1406 5352 -1396
rect 5092 -1456 5352 -1406
rect 5412 -1456 5422 -1396
rect 5022 -1466 5422 -1456
rect 5480 -1046 5880 -1036
rect 5480 -1106 5490 -1046
rect 5550 -1096 5810 -1046
rect 5550 -1106 5560 -1096
rect 5480 -1116 5560 -1106
rect 5800 -1106 5810 -1096
rect 5870 -1106 5880 -1046
rect 5800 -1116 5880 -1106
rect 5480 -1386 5540 -1116
rect 5810 -1126 5880 -1116
rect 5620 -1176 5650 -1156
rect 5600 -1216 5650 -1176
rect 5710 -1176 5740 -1156
rect 5710 -1216 5760 -1176
rect 5600 -1286 5760 -1216
rect 5600 -1326 5650 -1286
rect 5620 -1346 5650 -1326
rect 5710 -1326 5760 -1286
rect 5710 -1346 5740 -1326
rect 5820 -1386 5880 -1126
rect 5480 -1396 5560 -1386
rect 5480 -1456 5490 -1396
rect 5550 -1406 5560 -1396
rect 5800 -1396 5880 -1386
rect 5800 -1406 5810 -1396
rect 5550 -1456 5810 -1406
rect 5870 -1456 5880 -1396
rect 5480 -1466 5880 -1456
rect 5936 -1046 6336 -1036
rect 5936 -1106 5946 -1046
rect 6006 -1096 6266 -1046
rect 6006 -1106 6016 -1096
rect 5936 -1116 6016 -1106
rect 6256 -1106 6266 -1096
rect 6326 -1106 6336 -1046
rect 6256 -1116 6336 -1106
rect 5936 -1386 5996 -1116
rect 6266 -1126 6336 -1116
rect 6076 -1176 6106 -1156
rect 6056 -1216 6106 -1176
rect 6166 -1176 6196 -1156
rect 6166 -1216 6216 -1176
rect 6056 -1286 6216 -1216
rect 6056 -1326 6106 -1286
rect 6076 -1346 6106 -1326
rect 6166 -1326 6216 -1286
rect 6166 -1346 6196 -1326
rect 6276 -1386 6336 -1126
rect 5936 -1396 6016 -1386
rect 5936 -1456 5946 -1396
rect 6006 -1406 6016 -1396
rect 6256 -1396 6336 -1386
rect 6256 -1406 6266 -1396
rect 6006 -1456 6266 -1406
rect 6326 -1456 6336 -1396
rect 5936 -1466 6336 -1456
rect 6392 -1046 6792 -1036
rect 6392 -1106 6402 -1046
rect 6462 -1096 6722 -1046
rect 6462 -1106 6472 -1096
rect 6392 -1116 6472 -1106
rect 6712 -1106 6722 -1096
rect 6782 -1106 6792 -1046
rect 6712 -1116 6792 -1106
rect 6392 -1386 6452 -1116
rect 6722 -1126 6792 -1116
rect 6532 -1176 6562 -1156
rect 6512 -1216 6562 -1176
rect 6622 -1176 6652 -1156
rect 6622 -1216 6672 -1176
rect 6512 -1286 6672 -1216
rect 6512 -1326 6562 -1286
rect 6532 -1346 6562 -1326
rect 6622 -1326 6672 -1286
rect 6622 -1346 6652 -1326
rect 6732 -1386 6792 -1126
rect 6392 -1396 6472 -1386
rect 6392 -1456 6402 -1396
rect 6462 -1406 6472 -1396
rect 6712 -1396 6792 -1386
rect 6712 -1406 6722 -1396
rect 6462 -1456 6722 -1406
rect 6782 -1456 6792 -1396
rect 6392 -1466 6792 -1456
rect 6850 -1046 7250 -1036
rect 6850 -1106 6860 -1046
rect 6920 -1096 7180 -1046
rect 6920 -1106 6930 -1096
rect 6850 -1116 6930 -1106
rect 7170 -1106 7180 -1096
rect 7240 -1106 7250 -1046
rect 7170 -1116 7250 -1106
rect 6850 -1386 6910 -1116
rect 7180 -1126 7250 -1116
rect 6990 -1176 7020 -1156
rect 6970 -1216 7020 -1176
rect 7080 -1176 7110 -1156
rect 7080 -1216 7130 -1176
rect 6970 -1286 7130 -1216
rect 6970 -1326 7020 -1286
rect 6990 -1346 7020 -1326
rect 7080 -1326 7130 -1286
rect 7080 -1346 7110 -1326
rect 7190 -1386 7250 -1126
rect 6850 -1396 6930 -1386
rect 6850 -1456 6860 -1396
rect 6920 -1406 6930 -1396
rect 7170 -1396 7250 -1386
rect 7170 -1406 7180 -1396
rect 6920 -1456 7180 -1406
rect 7240 -1456 7250 -1396
rect 6850 -1466 7250 -1456
rect 7306 -1046 7706 -1036
rect 7306 -1106 7316 -1046
rect 7376 -1096 7636 -1046
rect 7376 -1106 7386 -1096
rect 7306 -1116 7386 -1106
rect 7626 -1106 7636 -1096
rect 7696 -1106 7706 -1046
rect 7626 -1116 7706 -1106
rect 7306 -1386 7366 -1116
rect 7636 -1126 7706 -1116
rect 7446 -1176 7476 -1156
rect 7426 -1216 7476 -1176
rect 7536 -1176 7566 -1156
rect 7536 -1216 7586 -1176
rect 7426 -1286 7586 -1216
rect 7426 -1326 7476 -1286
rect 7446 -1346 7476 -1326
rect 7536 -1326 7586 -1286
rect 7536 -1346 7566 -1326
rect 7646 -1386 7706 -1126
rect 7306 -1396 7386 -1386
rect 7306 -1456 7316 -1396
rect 7376 -1406 7386 -1396
rect 7626 -1396 7706 -1386
rect 7626 -1406 7636 -1396
rect 7376 -1456 7636 -1406
rect 7696 -1456 7706 -1396
rect 7306 -1466 7706 -1456
rect 7762 -1046 8162 -1036
rect 7762 -1106 7772 -1046
rect 7832 -1096 8092 -1046
rect 7832 -1106 7842 -1096
rect 7762 -1116 7842 -1106
rect 8082 -1106 8092 -1096
rect 8152 -1106 8162 -1046
rect 8082 -1116 8162 -1106
rect 7762 -1386 7822 -1116
rect 8092 -1126 8162 -1116
rect 7902 -1176 7932 -1156
rect 7882 -1216 7932 -1176
rect 7992 -1176 8022 -1156
rect 7992 -1216 8042 -1176
rect 7882 -1286 8042 -1216
rect 7882 -1326 7932 -1286
rect 7902 -1346 7932 -1326
rect 7992 -1326 8042 -1286
rect 7992 -1346 8022 -1326
rect 8102 -1386 8162 -1126
rect 7762 -1396 7842 -1386
rect 7762 -1456 7772 -1396
rect 7832 -1406 7842 -1396
rect 8082 -1396 8162 -1386
rect 8082 -1406 8092 -1396
rect 7832 -1456 8092 -1406
rect 8152 -1456 8162 -1396
rect 7762 -1466 8162 -1456
rect 8236 -1046 8636 -1036
rect 8236 -1106 8246 -1046
rect 8306 -1096 8566 -1046
rect 8306 -1106 8316 -1096
rect 8236 -1116 8316 -1106
rect 8556 -1106 8566 -1096
rect 8626 -1106 8636 -1046
rect 8556 -1116 8636 -1106
rect 8236 -1386 8296 -1116
rect 8566 -1126 8636 -1116
rect 8376 -1176 8406 -1156
rect 8356 -1216 8406 -1176
rect 8466 -1176 8496 -1156
rect 8466 -1216 8516 -1176
rect 8356 -1286 8516 -1216
rect 8356 -1326 8406 -1286
rect 8376 -1346 8406 -1326
rect 8466 -1326 8516 -1286
rect 8466 -1346 8496 -1326
rect 8576 -1386 8636 -1126
rect 8236 -1396 8316 -1386
rect 8236 -1456 8246 -1396
rect 8306 -1406 8316 -1396
rect 8556 -1396 8636 -1386
rect 8556 -1406 8566 -1396
rect 8306 -1456 8566 -1406
rect 8626 -1456 8636 -1396
rect 8236 -1466 8636 -1456
rect 8692 -1046 9092 -1036
rect 8692 -1106 8702 -1046
rect 8762 -1096 9022 -1046
rect 8762 -1106 8772 -1096
rect 8692 -1116 8772 -1106
rect 9012 -1106 9022 -1096
rect 9082 -1106 9092 -1046
rect 9012 -1116 9092 -1106
rect 8692 -1386 8752 -1116
rect 9022 -1126 9092 -1116
rect 8832 -1176 8862 -1156
rect 8812 -1216 8862 -1176
rect 8922 -1176 8952 -1156
rect 8922 -1216 8972 -1176
rect 8812 -1286 8972 -1216
rect 8812 -1326 8862 -1286
rect 8832 -1346 8862 -1326
rect 8922 -1326 8972 -1286
rect 8922 -1346 8952 -1326
rect 9032 -1386 9092 -1126
rect 8692 -1396 8772 -1386
rect 8692 -1456 8702 -1396
rect 8762 -1406 8772 -1396
rect 9012 -1396 9092 -1386
rect 9012 -1406 9022 -1396
rect 8762 -1456 9022 -1406
rect 9082 -1456 9092 -1396
rect 8692 -1466 9092 -1456
rect 9150 -1046 9550 -1036
rect 9150 -1106 9160 -1046
rect 9220 -1096 9480 -1046
rect 9220 -1106 9230 -1096
rect 9150 -1116 9230 -1106
rect 9470 -1106 9480 -1096
rect 9540 -1106 9550 -1046
rect 9470 -1116 9550 -1106
rect 9150 -1386 9210 -1116
rect 9480 -1126 9550 -1116
rect 9290 -1176 9320 -1156
rect 9270 -1216 9320 -1176
rect 9380 -1176 9410 -1156
rect 9380 -1216 9430 -1176
rect 9270 -1286 9430 -1216
rect 9270 -1326 9320 -1286
rect 9290 -1346 9320 -1326
rect 9380 -1326 9430 -1286
rect 9380 -1346 9410 -1326
rect 9490 -1386 9550 -1126
rect 9150 -1396 9230 -1386
rect 9150 -1456 9160 -1396
rect 9220 -1406 9230 -1396
rect 9470 -1396 9550 -1386
rect 9470 -1406 9480 -1396
rect 9220 -1456 9480 -1406
rect 9540 -1456 9550 -1396
rect 9150 -1466 9550 -1456
rect 9606 -1046 10006 -1036
rect 9606 -1106 9616 -1046
rect 9676 -1096 9936 -1046
rect 9676 -1106 9686 -1096
rect 9606 -1116 9686 -1106
rect 9926 -1106 9936 -1096
rect 9996 -1106 10006 -1046
rect 9926 -1116 10006 -1106
rect 9606 -1386 9666 -1116
rect 9936 -1126 10006 -1116
rect 9746 -1176 9776 -1156
rect 9726 -1216 9776 -1176
rect 9836 -1176 9866 -1156
rect 9836 -1216 9886 -1176
rect 9726 -1286 9886 -1216
rect 9726 -1326 9776 -1286
rect 9746 -1346 9776 -1326
rect 9836 -1326 9886 -1286
rect 9836 -1346 9866 -1326
rect 9946 -1386 10006 -1126
rect 9606 -1396 9686 -1386
rect 9606 -1456 9616 -1396
rect 9676 -1406 9686 -1396
rect 9926 -1396 10006 -1386
rect 9926 -1406 9936 -1396
rect 9676 -1456 9936 -1406
rect 9996 -1456 10006 -1396
rect 9606 -1466 10006 -1456
rect 10062 -1046 10462 -1036
rect 10062 -1106 10072 -1046
rect 10132 -1096 10392 -1046
rect 10132 -1106 10142 -1096
rect 10062 -1116 10142 -1106
rect 10382 -1106 10392 -1096
rect 10452 -1106 10462 -1046
rect 10382 -1116 10462 -1106
rect 10062 -1386 10122 -1116
rect 10392 -1126 10462 -1116
rect 10202 -1176 10232 -1156
rect 10182 -1216 10232 -1176
rect 10292 -1176 10322 -1156
rect 10292 -1216 10342 -1176
rect 10182 -1286 10342 -1216
rect 10182 -1326 10232 -1286
rect 10202 -1346 10232 -1326
rect 10292 -1326 10342 -1286
rect 10292 -1346 10322 -1326
rect 10402 -1386 10462 -1126
rect 10062 -1396 10142 -1386
rect 10062 -1456 10072 -1396
rect 10132 -1406 10142 -1396
rect 10382 -1396 10462 -1386
rect 10382 -1406 10392 -1396
rect 10132 -1456 10392 -1406
rect 10452 -1456 10462 -1396
rect 10062 -1466 10462 -1456
rect 10520 -1046 10920 -1036
rect 10520 -1106 10530 -1046
rect 10590 -1096 10850 -1046
rect 10590 -1106 10600 -1096
rect 10520 -1116 10600 -1106
rect 10840 -1106 10850 -1096
rect 10910 -1106 10920 -1046
rect 10840 -1116 10920 -1106
rect 10520 -1386 10580 -1116
rect 10850 -1126 10920 -1116
rect 10660 -1176 10690 -1156
rect 10640 -1216 10690 -1176
rect 10750 -1176 10780 -1156
rect 10750 -1216 10800 -1176
rect 10640 -1286 10800 -1216
rect 10640 -1326 10690 -1286
rect 10660 -1346 10690 -1326
rect 10750 -1326 10800 -1286
rect 10750 -1346 10780 -1326
rect 10860 -1386 10920 -1126
rect 10520 -1396 10600 -1386
rect 10520 -1456 10530 -1396
rect 10590 -1406 10600 -1396
rect 10840 -1396 10920 -1386
rect 10840 -1406 10850 -1396
rect 10590 -1456 10850 -1406
rect 10910 -1456 10920 -1396
rect 10520 -1466 10920 -1456
rect 10976 -1046 11376 -1036
rect 10976 -1106 10986 -1046
rect 11046 -1096 11306 -1046
rect 11046 -1106 11056 -1096
rect 10976 -1116 11056 -1106
rect 11296 -1106 11306 -1096
rect 11366 -1106 11376 -1046
rect 11296 -1116 11376 -1106
rect 10976 -1386 11036 -1116
rect 11306 -1126 11376 -1116
rect 11116 -1176 11146 -1156
rect 11096 -1216 11146 -1176
rect 11206 -1176 11236 -1156
rect 11206 -1216 11256 -1176
rect 11096 -1286 11256 -1216
rect 11096 -1326 11146 -1286
rect 11116 -1346 11146 -1326
rect 11206 -1326 11256 -1286
rect 11206 -1346 11236 -1326
rect 11316 -1386 11376 -1126
rect 10976 -1396 11056 -1386
rect 10976 -1456 10986 -1396
rect 11046 -1406 11056 -1396
rect 11296 -1396 11376 -1386
rect 11296 -1406 11306 -1396
rect 11046 -1456 11306 -1406
rect 11366 -1456 11376 -1396
rect 10976 -1466 11376 -1456
rect 11432 -1046 11832 -1036
rect 11432 -1106 11442 -1046
rect 11502 -1096 11762 -1046
rect 11502 -1106 11512 -1096
rect 11432 -1116 11512 -1106
rect 11752 -1106 11762 -1096
rect 11822 -1106 11832 -1046
rect 11752 -1116 11832 -1106
rect 11432 -1386 11492 -1116
rect 11762 -1126 11832 -1116
rect 11572 -1176 11602 -1156
rect 11552 -1216 11602 -1176
rect 11662 -1176 11692 -1156
rect 11662 -1216 11712 -1176
rect 11552 -1286 11712 -1216
rect 11552 -1326 11602 -1286
rect 11572 -1346 11602 -1326
rect 11662 -1326 11712 -1286
rect 11662 -1346 11692 -1326
rect 11772 -1386 11832 -1126
rect 11432 -1396 11512 -1386
rect 11432 -1456 11442 -1396
rect 11502 -1406 11512 -1396
rect 11752 -1396 11832 -1386
rect 11752 -1406 11762 -1396
rect 11502 -1456 11762 -1406
rect 11822 -1456 11832 -1396
rect 11432 -1466 11832 -1456
rect 11890 -1046 12290 -1036
rect 11890 -1106 11900 -1046
rect 11960 -1096 12220 -1046
rect 11960 -1106 11970 -1096
rect 11890 -1116 11970 -1106
rect 12210 -1106 12220 -1096
rect 12280 -1106 12290 -1046
rect 12210 -1116 12290 -1106
rect 11890 -1386 11950 -1116
rect 12220 -1126 12290 -1116
rect 12030 -1176 12060 -1156
rect 12010 -1216 12060 -1176
rect 12120 -1176 12150 -1156
rect 12120 -1216 12170 -1176
rect 12010 -1286 12170 -1216
rect 12010 -1326 12060 -1286
rect 12030 -1346 12060 -1326
rect 12120 -1326 12170 -1286
rect 12120 -1346 12150 -1326
rect 12230 -1386 12290 -1126
rect 11890 -1396 11970 -1386
rect 11890 -1456 11900 -1396
rect 11960 -1406 11970 -1396
rect 12210 -1396 12290 -1386
rect 12210 -1406 12220 -1396
rect 11960 -1456 12220 -1406
rect 12280 -1456 12290 -1396
rect 11890 -1466 12290 -1456
rect 12346 -1046 12746 -1036
rect 12346 -1106 12356 -1046
rect 12416 -1096 12676 -1046
rect 12416 -1106 12426 -1096
rect 12346 -1116 12426 -1106
rect 12666 -1106 12676 -1096
rect 12736 -1106 12746 -1046
rect 12666 -1116 12746 -1106
rect 12346 -1386 12406 -1116
rect 12676 -1126 12746 -1116
rect 12486 -1176 12516 -1156
rect 12466 -1216 12516 -1176
rect 12576 -1176 12606 -1156
rect 12576 -1216 12626 -1176
rect 12466 -1286 12626 -1216
rect 12466 -1326 12516 -1286
rect 12486 -1346 12516 -1326
rect 12576 -1326 12626 -1286
rect 12576 -1346 12606 -1326
rect 12686 -1386 12746 -1126
rect 12346 -1396 12426 -1386
rect 12346 -1456 12356 -1396
rect 12416 -1406 12426 -1396
rect 12666 -1396 12746 -1386
rect 12666 -1406 12676 -1396
rect 12416 -1456 12676 -1406
rect 12736 -1456 12746 -1396
rect 12346 -1466 12746 -1456
rect 12802 -1046 13202 -1036
rect 12802 -1106 12812 -1046
rect 12872 -1096 13132 -1046
rect 12872 -1106 12882 -1096
rect 12802 -1116 12882 -1106
rect 13122 -1106 13132 -1096
rect 13192 -1106 13202 -1046
rect 13122 -1116 13202 -1106
rect 12802 -1386 12862 -1116
rect 13132 -1126 13202 -1116
rect 12942 -1176 12972 -1156
rect 12922 -1216 12972 -1176
rect 13032 -1176 13062 -1156
rect 13032 -1216 13082 -1176
rect 12922 -1286 13082 -1216
rect 12922 -1326 12972 -1286
rect 12942 -1346 12972 -1326
rect 13032 -1326 13082 -1286
rect 13032 -1346 13062 -1326
rect 13142 -1386 13202 -1126
rect 12802 -1396 12882 -1386
rect 12802 -1456 12812 -1396
rect 12872 -1406 12882 -1396
rect 13122 -1396 13202 -1386
rect 13122 -1406 13132 -1396
rect 12872 -1456 13132 -1406
rect 13192 -1456 13202 -1396
rect 12802 -1466 13202 -1456
rect 13260 -1046 13660 -1036
rect 13260 -1106 13270 -1046
rect 13330 -1096 13590 -1046
rect 13330 -1106 13340 -1096
rect 13260 -1116 13340 -1106
rect 13580 -1106 13590 -1096
rect 13650 -1106 13660 -1046
rect 13580 -1116 13660 -1106
rect 13260 -1386 13320 -1116
rect 13590 -1126 13660 -1116
rect 13400 -1176 13430 -1156
rect 13380 -1216 13430 -1176
rect 13490 -1176 13520 -1156
rect 13490 -1216 13540 -1176
rect 13380 -1286 13540 -1216
rect 13380 -1326 13430 -1286
rect 13400 -1346 13430 -1326
rect 13490 -1326 13540 -1286
rect 13490 -1346 13520 -1326
rect 13600 -1386 13660 -1126
rect 13260 -1396 13340 -1386
rect 13260 -1456 13270 -1396
rect 13330 -1406 13340 -1396
rect 13580 -1396 13660 -1386
rect 13580 -1406 13590 -1396
rect 13330 -1456 13590 -1406
rect 13650 -1456 13660 -1396
rect 13260 -1466 13660 -1456
rect 13716 -1046 14116 -1036
rect 13716 -1106 13726 -1046
rect 13786 -1096 14046 -1046
rect 13786 -1106 13796 -1096
rect 13716 -1116 13796 -1106
rect 14036 -1106 14046 -1096
rect 14106 -1106 14116 -1046
rect 14036 -1116 14116 -1106
rect 13716 -1386 13776 -1116
rect 14046 -1126 14116 -1116
rect 13856 -1176 13886 -1156
rect 13836 -1216 13886 -1176
rect 13946 -1176 13976 -1156
rect 13946 -1216 13996 -1176
rect 13836 -1286 13996 -1216
rect 13836 -1326 13886 -1286
rect 13856 -1346 13886 -1326
rect 13946 -1326 13996 -1286
rect 13946 -1346 13976 -1326
rect 14056 -1386 14116 -1126
rect 13716 -1396 13796 -1386
rect 13716 -1456 13726 -1396
rect 13786 -1406 13796 -1396
rect 14036 -1396 14116 -1386
rect 14036 -1406 14046 -1396
rect 13786 -1456 14046 -1406
rect 14106 -1456 14116 -1396
rect 13716 -1466 14116 -1456
rect 14172 -1046 14572 -1036
rect 14172 -1106 14182 -1046
rect 14242 -1096 14502 -1046
rect 14242 -1106 14252 -1096
rect 14172 -1116 14252 -1106
rect 14492 -1106 14502 -1096
rect 14562 -1106 14572 -1046
rect 14492 -1116 14572 -1106
rect 14172 -1386 14232 -1116
rect 14502 -1126 14572 -1116
rect 14312 -1176 14342 -1156
rect 14292 -1216 14342 -1176
rect 14402 -1176 14432 -1156
rect 14402 -1216 14452 -1176
rect 14292 -1286 14452 -1216
rect 14292 -1326 14342 -1286
rect 14312 -1346 14342 -1326
rect 14402 -1326 14452 -1286
rect 14402 -1346 14432 -1326
rect 14512 -1386 14572 -1126
rect 14172 -1396 14252 -1386
rect 14172 -1456 14182 -1396
rect 14242 -1406 14252 -1396
rect 14492 -1396 14572 -1386
rect 14492 -1406 14502 -1396
rect 14242 -1456 14502 -1406
rect 14562 -1456 14572 -1396
rect 14172 -1466 14572 -1456
rect 14630 -1046 15030 -1036
rect 14630 -1106 14640 -1046
rect 14700 -1096 14960 -1046
rect 14700 -1106 14710 -1096
rect 14630 -1116 14710 -1106
rect 14950 -1106 14960 -1096
rect 15020 -1106 15030 -1046
rect 14950 -1116 15030 -1106
rect 14630 -1386 14690 -1116
rect 14960 -1126 15030 -1116
rect 14770 -1176 14800 -1156
rect 14750 -1216 14800 -1176
rect 14860 -1176 14890 -1156
rect 14860 -1216 14910 -1176
rect 14750 -1286 14910 -1216
rect 14750 -1326 14800 -1286
rect 14770 -1346 14800 -1326
rect 14860 -1326 14910 -1286
rect 14860 -1346 14890 -1326
rect 14970 -1386 15030 -1126
rect 14630 -1396 14710 -1386
rect 14630 -1456 14640 -1396
rect 14700 -1406 14710 -1396
rect 14950 -1396 15030 -1386
rect 14950 -1406 14960 -1396
rect 14700 -1456 14960 -1406
rect 15020 -1456 15030 -1396
rect 14630 -1466 15030 -1456
rect 15086 -1046 15486 -1036
rect 15086 -1106 15096 -1046
rect 15156 -1096 15416 -1046
rect 15156 -1106 15166 -1096
rect 15086 -1116 15166 -1106
rect 15406 -1106 15416 -1096
rect 15476 -1106 15486 -1046
rect 15406 -1116 15486 -1106
rect 15086 -1386 15146 -1116
rect 15416 -1126 15486 -1116
rect 15226 -1176 15256 -1156
rect 15206 -1216 15256 -1176
rect 15316 -1176 15346 -1156
rect 15316 -1216 15366 -1176
rect 15206 -1286 15366 -1216
rect 15206 -1326 15256 -1286
rect 15226 -1346 15256 -1326
rect 15316 -1326 15366 -1286
rect 15316 -1346 15346 -1326
rect 15426 -1386 15486 -1126
rect 15086 -1396 15166 -1386
rect 15086 -1456 15096 -1396
rect 15156 -1406 15166 -1396
rect 15406 -1396 15486 -1386
rect 15406 -1406 15416 -1396
rect 15156 -1456 15416 -1406
rect 15476 -1456 15486 -1396
rect 15086 -1466 15486 -1456
rect 0 -1562 400 -1552
rect 0 -1622 10 -1562
rect 70 -1612 330 -1562
rect 70 -1622 80 -1612
rect 0 -1632 80 -1622
rect 320 -1622 330 -1612
rect 390 -1622 400 -1562
rect 320 -1632 400 -1622
rect 0 -1902 60 -1632
rect 330 -1642 400 -1632
rect 140 -1692 170 -1672
rect 120 -1732 170 -1692
rect 230 -1692 260 -1672
rect 230 -1732 280 -1692
rect 120 -1802 280 -1732
rect 120 -1842 170 -1802
rect 140 -1862 170 -1842
rect 230 -1842 280 -1802
rect 230 -1862 260 -1842
rect 340 -1902 400 -1642
rect 0 -1912 80 -1902
rect 0 -1972 10 -1912
rect 70 -1922 80 -1912
rect 320 -1912 400 -1902
rect 320 -1922 330 -1912
rect 70 -1972 330 -1922
rect 390 -1972 400 -1912
rect 0 -1982 400 -1972
rect 456 -1562 856 -1552
rect 456 -1622 466 -1562
rect 526 -1612 786 -1562
rect 526 -1622 536 -1612
rect 456 -1632 536 -1622
rect 776 -1622 786 -1612
rect 846 -1622 856 -1562
rect 776 -1632 856 -1622
rect 456 -1902 516 -1632
rect 786 -1642 856 -1632
rect 596 -1692 626 -1672
rect 576 -1732 626 -1692
rect 686 -1692 716 -1672
rect 686 -1732 736 -1692
rect 576 -1802 736 -1732
rect 576 -1842 626 -1802
rect 596 -1862 626 -1842
rect 686 -1842 736 -1802
rect 686 -1862 716 -1842
rect 796 -1902 856 -1642
rect 456 -1912 536 -1902
rect 456 -1972 466 -1912
rect 526 -1922 536 -1912
rect 776 -1912 856 -1902
rect 776 -1922 786 -1912
rect 526 -1972 786 -1922
rect 846 -1972 856 -1912
rect 456 -1982 856 -1972
rect 912 -1562 1312 -1552
rect 912 -1622 922 -1562
rect 982 -1612 1242 -1562
rect 982 -1622 992 -1612
rect 912 -1632 992 -1622
rect 1232 -1622 1242 -1612
rect 1302 -1622 1312 -1562
rect 1232 -1632 1312 -1622
rect 912 -1902 972 -1632
rect 1242 -1642 1312 -1632
rect 1052 -1692 1082 -1672
rect 1032 -1732 1082 -1692
rect 1142 -1692 1172 -1672
rect 1142 -1732 1192 -1692
rect 1032 -1802 1192 -1732
rect 1032 -1842 1082 -1802
rect 1052 -1862 1082 -1842
rect 1142 -1842 1192 -1802
rect 1142 -1862 1172 -1842
rect 1252 -1902 1312 -1642
rect 912 -1912 992 -1902
rect 912 -1972 922 -1912
rect 982 -1922 992 -1912
rect 1232 -1912 1312 -1902
rect 1232 -1922 1242 -1912
rect 982 -1972 1242 -1922
rect 1302 -1972 1312 -1912
rect 912 -1982 1312 -1972
rect 1370 -1562 1770 -1552
rect 1370 -1622 1380 -1562
rect 1440 -1612 1700 -1562
rect 1440 -1622 1450 -1612
rect 1370 -1632 1450 -1622
rect 1690 -1622 1700 -1612
rect 1760 -1622 1770 -1562
rect 1690 -1632 1770 -1622
rect 1370 -1902 1430 -1632
rect 1700 -1642 1770 -1632
rect 1510 -1692 1540 -1672
rect 1490 -1732 1540 -1692
rect 1600 -1692 1630 -1672
rect 1600 -1732 1650 -1692
rect 1490 -1802 1650 -1732
rect 1490 -1842 1540 -1802
rect 1510 -1862 1540 -1842
rect 1600 -1842 1650 -1802
rect 1600 -1862 1630 -1842
rect 1710 -1902 1770 -1642
rect 1370 -1912 1450 -1902
rect 1370 -1972 1380 -1912
rect 1440 -1922 1450 -1912
rect 1690 -1912 1770 -1902
rect 1690 -1922 1700 -1912
rect 1440 -1972 1700 -1922
rect 1760 -1972 1770 -1912
rect 1370 -1982 1770 -1972
rect 1826 -1562 2226 -1552
rect 1826 -1622 1836 -1562
rect 1896 -1612 2156 -1562
rect 1896 -1622 1906 -1612
rect 1826 -1632 1906 -1622
rect 2146 -1622 2156 -1612
rect 2216 -1622 2226 -1562
rect 2146 -1632 2226 -1622
rect 1826 -1902 1886 -1632
rect 2156 -1642 2226 -1632
rect 1966 -1692 1996 -1672
rect 1946 -1732 1996 -1692
rect 2056 -1692 2086 -1672
rect 2056 -1732 2106 -1692
rect 1946 -1802 2106 -1732
rect 1946 -1842 1996 -1802
rect 1966 -1862 1996 -1842
rect 2056 -1842 2106 -1802
rect 2056 -1862 2086 -1842
rect 2166 -1902 2226 -1642
rect 1826 -1912 1906 -1902
rect 1826 -1972 1836 -1912
rect 1896 -1922 1906 -1912
rect 2146 -1912 2226 -1902
rect 2146 -1922 2156 -1912
rect 1896 -1972 2156 -1922
rect 2216 -1972 2226 -1912
rect 1826 -1982 2226 -1972
rect 2282 -1562 2682 -1552
rect 2282 -1622 2292 -1562
rect 2352 -1612 2612 -1562
rect 2352 -1622 2362 -1612
rect 2282 -1632 2362 -1622
rect 2602 -1622 2612 -1612
rect 2672 -1622 2682 -1562
rect 2602 -1632 2682 -1622
rect 2282 -1902 2342 -1632
rect 2612 -1642 2682 -1632
rect 2422 -1692 2452 -1672
rect 2402 -1732 2452 -1692
rect 2512 -1692 2542 -1672
rect 2512 -1732 2562 -1692
rect 2402 -1802 2562 -1732
rect 2402 -1842 2452 -1802
rect 2422 -1862 2452 -1842
rect 2512 -1842 2562 -1802
rect 2512 -1862 2542 -1842
rect 2622 -1902 2682 -1642
rect 2282 -1912 2362 -1902
rect 2282 -1972 2292 -1912
rect 2352 -1922 2362 -1912
rect 2602 -1912 2682 -1902
rect 2602 -1922 2612 -1912
rect 2352 -1972 2612 -1922
rect 2672 -1972 2682 -1912
rect 2282 -1982 2682 -1972
rect 2740 -1562 3140 -1552
rect 2740 -1622 2750 -1562
rect 2810 -1612 3070 -1562
rect 2810 -1622 2820 -1612
rect 2740 -1632 2820 -1622
rect 3060 -1622 3070 -1612
rect 3130 -1622 3140 -1562
rect 3060 -1632 3140 -1622
rect 2740 -1902 2800 -1632
rect 3070 -1642 3140 -1632
rect 2880 -1692 2910 -1672
rect 2860 -1732 2910 -1692
rect 2970 -1692 3000 -1672
rect 2970 -1732 3020 -1692
rect 2860 -1802 3020 -1732
rect 2860 -1842 2910 -1802
rect 2880 -1862 2910 -1842
rect 2970 -1842 3020 -1802
rect 2970 -1862 3000 -1842
rect 3080 -1902 3140 -1642
rect 2740 -1912 2820 -1902
rect 2740 -1972 2750 -1912
rect 2810 -1922 2820 -1912
rect 3060 -1912 3140 -1902
rect 3060 -1922 3070 -1912
rect 2810 -1972 3070 -1922
rect 3130 -1972 3140 -1912
rect 2740 -1982 3140 -1972
rect 3196 -1562 3596 -1552
rect 3196 -1622 3206 -1562
rect 3266 -1612 3526 -1562
rect 3266 -1622 3276 -1612
rect 3196 -1632 3276 -1622
rect 3516 -1622 3526 -1612
rect 3586 -1622 3596 -1562
rect 3516 -1632 3596 -1622
rect 3196 -1902 3256 -1632
rect 3526 -1642 3596 -1632
rect 3336 -1692 3366 -1672
rect 3316 -1732 3366 -1692
rect 3426 -1692 3456 -1672
rect 3426 -1732 3476 -1692
rect 3316 -1802 3476 -1732
rect 3316 -1842 3366 -1802
rect 3336 -1862 3366 -1842
rect 3426 -1842 3476 -1802
rect 3426 -1862 3456 -1842
rect 3536 -1902 3596 -1642
rect 3196 -1912 3276 -1902
rect 3196 -1972 3206 -1912
rect 3266 -1922 3276 -1912
rect 3516 -1912 3596 -1902
rect 3516 -1922 3526 -1912
rect 3266 -1972 3526 -1922
rect 3586 -1972 3596 -1912
rect 3196 -1982 3596 -1972
rect 3652 -1562 4052 -1552
rect 3652 -1622 3662 -1562
rect 3722 -1612 3982 -1562
rect 3722 -1622 3732 -1612
rect 3652 -1632 3732 -1622
rect 3972 -1622 3982 -1612
rect 4042 -1622 4052 -1562
rect 3972 -1632 4052 -1622
rect 3652 -1902 3712 -1632
rect 3982 -1642 4052 -1632
rect 3792 -1692 3822 -1672
rect 3772 -1732 3822 -1692
rect 3882 -1692 3912 -1672
rect 3882 -1732 3932 -1692
rect 3772 -1802 3932 -1732
rect 3772 -1842 3822 -1802
rect 3792 -1862 3822 -1842
rect 3882 -1842 3932 -1802
rect 3882 -1862 3912 -1842
rect 3992 -1902 4052 -1642
rect 3652 -1912 3732 -1902
rect 3652 -1972 3662 -1912
rect 3722 -1922 3732 -1912
rect 3972 -1912 4052 -1902
rect 3972 -1922 3982 -1912
rect 3722 -1972 3982 -1922
rect 4042 -1972 4052 -1912
rect 3652 -1982 4052 -1972
rect 4110 -1562 4510 -1552
rect 4110 -1622 4120 -1562
rect 4180 -1612 4440 -1562
rect 4180 -1622 4190 -1612
rect 4110 -1632 4190 -1622
rect 4430 -1622 4440 -1612
rect 4500 -1622 4510 -1562
rect 4430 -1632 4510 -1622
rect 4110 -1902 4170 -1632
rect 4440 -1642 4510 -1632
rect 4250 -1692 4280 -1672
rect 4230 -1732 4280 -1692
rect 4340 -1692 4370 -1672
rect 4340 -1732 4390 -1692
rect 4230 -1802 4390 -1732
rect 4230 -1842 4280 -1802
rect 4250 -1862 4280 -1842
rect 4340 -1842 4390 -1802
rect 4340 -1862 4370 -1842
rect 4450 -1902 4510 -1642
rect 4110 -1912 4190 -1902
rect 4110 -1972 4120 -1912
rect 4180 -1922 4190 -1912
rect 4430 -1912 4510 -1902
rect 4430 -1922 4440 -1912
rect 4180 -1972 4440 -1922
rect 4500 -1972 4510 -1912
rect 4110 -1982 4510 -1972
rect 4566 -1562 4966 -1552
rect 4566 -1622 4576 -1562
rect 4636 -1612 4896 -1562
rect 4636 -1622 4646 -1612
rect 4566 -1632 4646 -1622
rect 4886 -1622 4896 -1612
rect 4956 -1622 4966 -1562
rect 4886 -1632 4966 -1622
rect 4566 -1902 4626 -1632
rect 4896 -1642 4966 -1632
rect 4706 -1692 4736 -1672
rect 4686 -1732 4736 -1692
rect 4796 -1692 4826 -1672
rect 4796 -1732 4846 -1692
rect 4686 -1802 4846 -1732
rect 4686 -1842 4736 -1802
rect 4706 -1862 4736 -1842
rect 4796 -1842 4846 -1802
rect 4796 -1862 4826 -1842
rect 4906 -1902 4966 -1642
rect 4566 -1912 4646 -1902
rect 4566 -1972 4576 -1912
rect 4636 -1922 4646 -1912
rect 4886 -1912 4966 -1902
rect 4886 -1922 4896 -1912
rect 4636 -1972 4896 -1922
rect 4956 -1972 4966 -1912
rect 4566 -1982 4966 -1972
rect 5022 -1562 5422 -1552
rect 5022 -1622 5032 -1562
rect 5092 -1612 5352 -1562
rect 5092 -1622 5102 -1612
rect 5022 -1632 5102 -1622
rect 5342 -1622 5352 -1612
rect 5412 -1622 5422 -1562
rect 5342 -1632 5422 -1622
rect 5022 -1902 5082 -1632
rect 5352 -1642 5422 -1632
rect 5162 -1692 5192 -1672
rect 5142 -1732 5192 -1692
rect 5252 -1692 5282 -1672
rect 5252 -1732 5302 -1692
rect 5142 -1802 5302 -1732
rect 5142 -1842 5192 -1802
rect 5162 -1862 5192 -1842
rect 5252 -1842 5302 -1802
rect 5252 -1862 5282 -1842
rect 5362 -1902 5422 -1642
rect 5022 -1912 5102 -1902
rect 5022 -1972 5032 -1912
rect 5092 -1922 5102 -1912
rect 5342 -1912 5422 -1902
rect 5342 -1922 5352 -1912
rect 5092 -1972 5352 -1922
rect 5412 -1972 5422 -1912
rect 5022 -1982 5422 -1972
rect 5480 -1562 5880 -1552
rect 5480 -1622 5490 -1562
rect 5550 -1612 5810 -1562
rect 5550 -1622 5560 -1612
rect 5480 -1632 5560 -1622
rect 5800 -1622 5810 -1612
rect 5870 -1622 5880 -1562
rect 5800 -1632 5880 -1622
rect 5480 -1902 5540 -1632
rect 5810 -1642 5880 -1632
rect 5620 -1692 5650 -1672
rect 5600 -1732 5650 -1692
rect 5710 -1692 5740 -1672
rect 5710 -1732 5760 -1692
rect 5600 -1802 5760 -1732
rect 5600 -1842 5650 -1802
rect 5620 -1862 5650 -1842
rect 5710 -1842 5760 -1802
rect 5710 -1862 5740 -1842
rect 5820 -1902 5880 -1642
rect 5480 -1912 5560 -1902
rect 5480 -1972 5490 -1912
rect 5550 -1922 5560 -1912
rect 5800 -1912 5880 -1902
rect 5800 -1922 5810 -1912
rect 5550 -1972 5810 -1922
rect 5870 -1972 5880 -1912
rect 5480 -1982 5880 -1972
rect 5936 -1562 6336 -1552
rect 5936 -1622 5946 -1562
rect 6006 -1612 6266 -1562
rect 6006 -1622 6016 -1612
rect 5936 -1632 6016 -1622
rect 6256 -1622 6266 -1612
rect 6326 -1622 6336 -1562
rect 6256 -1632 6336 -1622
rect 5936 -1902 5996 -1632
rect 6266 -1642 6336 -1632
rect 6076 -1692 6106 -1672
rect 6056 -1732 6106 -1692
rect 6166 -1692 6196 -1672
rect 6166 -1732 6216 -1692
rect 6056 -1802 6216 -1732
rect 6056 -1842 6106 -1802
rect 6076 -1862 6106 -1842
rect 6166 -1842 6216 -1802
rect 6166 -1862 6196 -1842
rect 6276 -1902 6336 -1642
rect 5936 -1912 6016 -1902
rect 5936 -1972 5946 -1912
rect 6006 -1922 6016 -1912
rect 6256 -1912 6336 -1902
rect 6256 -1922 6266 -1912
rect 6006 -1972 6266 -1922
rect 6326 -1972 6336 -1912
rect 5936 -1982 6336 -1972
rect 6392 -1562 6792 -1552
rect 6392 -1622 6402 -1562
rect 6462 -1612 6722 -1562
rect 6462 -1622 6472 -1612
rect 6392 -1632 6472 -1622
rect 6712 -1622 6722 -1612
rect 6782 -1622 6792 -1562
rect 6712 -1632 6792 -1622
rect 6392 -1902 6452 -1632
rect 6722 -1642 6792 -1632
rect 6532 -1692 6562 -1672
rect 6512 -1732 6562 -1692
rect 6622 -1692 6652 -1672
rect 6622 -1732 6672 -1692
rect 6512 -1802 6672 -1732
rect 6512 -1842 6562 -1802
rect 6532 -1862 6562 -1842
rect 6622 -1842 6672 -1802
rect 6622 -1862 6652 -1842
rect 6732 -1902 6792 -1642
rect 6392 -1912 6472 -1902
rect 6392 -1972 6402 -1912
rect 6462 -1922 6472 -1912
rect 6712 -1912 6792 -1902
rect 6712 -1922 6722 -1912
rect 6462 -1972 6722 -1922
rect 6782 -1972 6792 -1912
rect 6392 -1982 6792 -1972
rect 6850 -1562 7250 -1552
rect 6850 -1622 6860 -1562
rect 6920 -1612 7180 -1562
rect 6920 -1622 6930 -1612
rect 6850 -1632 6930 -1622
rect 7170 -1622 7180 -1612
rect 7240 -1622 7250 -1562
rect 7170 -1632 7250 -1622
rect 6850 -1902 6910 -1632
rect 7180 -1642 7250 -1632
rect 6990 -1692 7020 -1672
rect 6970 -1732 7020 -1692
rect 7080 -1692 7110 -1672
rect 7080 -1732 7130 -1692
rect 6970 -1802 7130 -1732
rect 6970 -1842 7020 -1802
rect 6990 -1862 7020 -1842
rect 7080 -1842 7130 -1802
rect 7080 -1862 7110 -1842
rect 7190 -1902 7250 -1642
rect 6850 -1912 6930 -1902
rect 6850 -1972 6860 -1912
rect 6920 -1922 6930 -1912
rect 7170 -1912 7250 -1902
rect 7170 -1922 7180 -1912
rect 6920 -1972 7180 -1922
rect 7240 -1972 7250 -1912
rect 6850 -1982 7250 -1972
rect 7306 -1562 7706 -1552
rect 7306 -1622 7316 -1562
rect 7376 -1612 7636 -1562
rect 7376 -1622 7386 -1612
rect 7306 -1632 7386 -1622
rect 7626 -1622 7636 -1612
rect 7696 -1622 7706 -1562
rect 7626 -1632 7706 -1622
rect 7306 -1902 7366 -1632
rect 7636 -1642 7706 -1632
rect 7446 -1692 7476 -1672
rect 7426 -1732 7476 -1692
rect 7536 -1692 7566 -1672
rect 7536 -1732 7586 -1692
rect 7426 -1802 7586 -1732
rect 7426 -1842 7476 -1802
rect 7446 -1862 7476 -1842
rect 7536 -1842 7586 -1802
rect 7536 -1862 7566 -1842
rect 7646 -1902 7706 -1642
rect 7306 -1912 7386 -1902
rect 7306 -1972 7316 -1912
rect 7376 -1922 7386 -1912
rect 7626 -1912 7706 -1902
rect 7626 -1922 7636 -1912
rect 7376 -1972 7636 -1922
rect 7696 -1972 7706 -1912
rect 7306 -1982 7706 -1972
rect 7762 -1562 8162 -1552
rect 7762 -1622 7772 -1562
rect 7832 -1612 8092 -1562
rect 7832 -1622 7842 -1612
rect 7762 -1632 7842 -1622
rect 8082 -1622 8092 -1612
rect 8152 -1622 8162 -1562
rect 8082 -1632 8162 -1622
rect 7762 -1902 7822 -1632
rect 8092 -1642 8162 -1632
rect 7902 -1692 7932 -1672
rect 7882 -1732 7932 -1692
rect 7992 -1692 8022 -1672
rect 7992 -1732 8042 -1692
rect 7882 -1802 8042 -1732
rect 7882 -1842 7932 -1802
rect 7902 -1862 7932 -1842
rect 7992 -1842 8042 -1802
rect 7992 -1862 8022 -1842
rect 8102 -1902 8162 -1642
rect 7762 -1912 7842 -1902
rect 7762 -1972 7772 -1912
rect 7832 -1922 7842 -1912
rect 8082 -1912 8162 -1902
rect 8082 -1922 8092 -1912
rect 7832 -1972 8092 -1922
rect 8152 -1972 8162 -1912
rect 7762 -1982 8162 -1972
rect 8236 -1562 8636 -1552
rect 8236 -1622 8246 -1562
rect 8306 -1612 8566 -1562
rect 8306 -1622 8316 -1612
rect 8236 -1632 8316 -1622
rect 8556 -1622 8566 -1612
rect 8626 -1622 8636 -1562
rect 8556 -1632 8636 -1622
rect 8236 -1902 8296 -1632
rect 8566 -1642 8636 -1632
rect 8376 -1692 8406 -1672
rect 8356 -1732 8406 -1692
rect 8466 -1692 8496 -1672
rect 8466 -1732 8516 -1692
rect 8356 -1802 8516 -1732
rect 8356 -1842 8406 -1802
rect 8376 -1862 8406 -1842
rect 8466 -1842 8516 -1802
rect 8466 -1862 8496 -1842
rect 8576 -1902 8636 -1642
rect 8236 -1912 8316 -1902
rect 8236 -1972 8246 -1912
rect 8306 -1922 8316 -1912
rect 8556 -1912 8636 -1902
rect 8556 -1922 8566 -1912
rect 8306 -1972 8566 -1922
rect 8626 -1972 8636 -1912
rect 8236 -1982 8636 -1972
rect 8692 -1562 9092 -1552
rect 8692 -1622 8702 -1562
rect 8762 -1612 9022 -1562
rect 8762 -1622 8772 -1612
rect 8692 -1632 8772 -1622
rect 9012 -1622 9022 -1612
rect 9082 -1622 9092 -1562
rect 9012 -1632 9092 -1622
rect 8692 -1902 8752 -1632
rect 9022 -1642 9092 -1632
rect 8832 -1692 8862 -1672
rect 8812 -1732 8862 -1692
rect 8922 -1692 8952 -1672
rect 8922 -1732 8972 -1692
rect 8812 -1802 8972 -1732
rect 8812 -1842 8862 -1802
rect 8832 -1862 8862 -1842
rect 8922 -1842 8972 -1802
rect 8922 -1862 8952 -1842
rect 9032 -1902 9092 -1642
rect 8692 -1912 8772 -1902
rect 8692 -1972 8702 -1912
rect 8762 -1922 8772 -1912
rect 9012 -1912 9092 -1902
rect 9012 -1922 9022 -1912
rect 8762 -1972 9022 -1922
rect 9082 -1972 9092 -1912
rect 8692 -1982 9092 -1972
rect 9150 -1562 9550 -1552
rect 9150 -1622 9160 -1562
rect 9220 -1612 9480 -1562
rect 9220 -1622 9230 -1612
rect 9150 -1632 9230 -1622
rect 9470 -1622 9480 -1612
rect 9540 -1622 9550 -1562
rect 9470 -1632 9550 -1622
rect 9150 -1902 9210 -1632
rect 9480 -1642 9550 -1632
rect 9290 -1692 9320 -1672
rect 9270 -1732 9320 -1692
rect 9380 -1692 9410 -1672
rect 9380 -1732 9430 -1692
rect 9270 -1802 9430 -1732
rect 9270 -1842 9320 -1802
rect 9290 -1862 9320 -1842
rect 9380 -1842 9430 -1802
rect 9380 -1862 9410 -1842
rect 9490 -1902 9550 -1642
rect 9150 -1912 9230 -1902
rect 9150 -1972 9160 -1912
rect 9220 -1922 9230 -1912
rect 9470 -1912 9550 -1902
rect 9470 -1922 9480 -1912
rect 9220 -1972 9480 -1922
rect 9540 -1972 9550 -1912
rect 9150 -1982 9550 -1972
rect 9606 -1562 10006 -1552
rect 9606 -1622 9616 -1562
rect 9676 -1612 9936 -1562
rect 9676 -1622 9686 -1612
rect 9606 -1632 9686 -1622
rect 9926 -1622 9936 -1612
rect 9996 -1622 10006 -1562
rect 9926 -1632 10006 -1622
rect 9606 -1902 9666 -1632
rect 9936 -1642 10006 -1632
rect 9746 -1692 9776 -1672
rect 9726 -1732 9776 -1692
rect 9836 -1692 9866 -1672
rect 9836 -1732 9886 -1692
rect 9726 -1802 9886 -1732
rect 9726 -1842 9776 -1802
rect 9746 -1862 9776 -1842
rect 9836 -1842 9886 -1802
rect 9836 -1862 9866 -1842
rect 9946 -1902 10006 -1642
rect 9606 -1912 9686 -1902
rect 9606 -1972 9616 -1912
rect 9676 -1922 9686 -1912
rect 9926 -1912 10006 -1902
rect 9926 -1922 9936 -1912
rect 9676 -1972 9936 -1922
rect 9996 -1972 10006 -1912
rect 9606 -1982 10006 -1972
rect 10062 -1562 10462 -1552
rect 10062 -1622 10072 -1562
rect 10132 -1612 10392 -1562
rect 10132 -1622 10142 -1612
rect 10062 -1632 10142 -1622
rect 10382 -1622 10392 -1612
rect 10452 -1622 10462 -1562
rect 10382 -1632 10462 -1622
rect 10062 -1902 10122 -1632
rect 10392 -1642 10462 -1632
rect 10202 -1692 10232 -1672
rect 10182 -1732 10232 -1692
rect 10292 -1692 10322 -1672
rect 10292 -1732 10342 -1692
rect 10182 -1802 10342 -1732
rect 10182 -1842 10232 -1802
rect 10202 -1862 10232 -1842
rect 10292 -1842 10342 -1802
rect 10292 -1862 10322 -1842
rect 10402 -1902 10462 -1642
rect 10062 -1912 10142 -1902
rect 10062 -1972 10072 -1912
rect 10132 -1922 10142 -1912
rect 10382 -1912 10462 -1902
rect 10382 -1922 10392 -1912
rect 10132 -1972 10392 -1922
rect 10452 -1972 10462 -1912
rect 10062 -1982 10462 -1972
rect 10520 -1562 10920 -1552
rect 10520 -1622 10530 -1562
rect 10590 -1612 10850 -1562
rect 10590 -1622 10600 -1612
rect 10520 -1632 10600 -1622
rect 10840 -1622 10850 -1612
rect 10910 -1622 10920 -1562
rect 10840 -1632 10920 -1622
rect 10520 -1902 10580 -1632
rect 10850 -1642 10920 -1632
rect 10660 -1692 10690 -1672
rect 10640 -1732 10690 -1692
rect 10750 -1692 10780 -1672
rect 10750 -1732 10800 -1692
rect 10640 -1802 10800 -1732
rect 10640 -1842 10690 -1802
rect 10660 -1862 10690 -1842
rect 10750 -1842 10800 -1802
rect 10750 -1862 10780 -1842
rect 10860 -1902 10920 -1642
rect 10520 -1912 10600 -1902
rect 10520 -1972 10530 -1912
rect 10590 -1922 10600 -1912
rect 10840 -1912 10920 -1902
rect 10840 -1922 10850 -1912
rect 10590 -1972 10850 -1922
rect 10910 -1972 10920 -1912
rect 10520 -1982 10920 -1972
rect 10976 -1562 11376 -1552
rect 10976 -1622 10986 -1562
rect 11046 -1612 11306 -1562
rect 11046 -1622 11056 -1612
rect 10976 -1632 11056 -1622
rect 11296 -1622 11306 -1612
rect 11366 -1622 11376 -1562
rect 11296 -1632 11376 -1622
rect 10976 -1902 11036 -1632
rect 11306 -1642 11376 -1632
rect 11116 -1692 11146 -1672
rect 11096 -1732 11146 -1692
rect 11206 -1692 11236 -1672
rect 11206 -1732 11256 -1692
rect 11096 -1802 11256 -1732
rect 11096 -1842 11146 -1802
rect 11116 -1862 11146 -1842
rect 11206 -1842 11256 -1802
rect 11206 -1862 11236 -1842
rect 11316 -1902 11376 -1642
rect 10976 -1912 11056 -1902
rect 10976 -1972 10986 -1912
rect 11046 -1922 11056 -1912
rect 11296 -1912 11376 -1902
rect 11296 -1922 11306 -1912
rect 11046 -1972 11306 -1922
rect 11366 -1972 11376 -1912
rect 10976 -1982 11376 -1972
rect 11432 -1562 11832 -1552
rect 11432 -1622 11442 -1562
rect 11502 -1612 11762 -1562
rect 11502 -1622 11512 -1612
rect 11432 -1632 11512 -1622
rect 11752 -1622 11762 -1612
rect 11822 -1622 11832 -1562
rect 11752 -1632 11832 -1622
rect 11432 -1902 11492 -1632
rect 11762 -1642 11832 -1632
rect 11572 -1692 11602 -1672
rect 11552 -1732 11602 -1692
rect 11662 -1692 11692 -1672
rect 11662 -1732 11712 -1692
rect 11552 -1802 11712 -1732
rect 11552 -1842 11602 -1802
rect 11572 -1862 11602 -1842
rect 11662 -1842 11712 -1802
rect 11662 -1862 11692 -1842
rect 11772 -1902 11832 -1642
rect 11432 -1912 11512 -1902
rect 11432 -1972 11442 -1912
rect 11502 -1922 11512 -1912
rect 11752 -1912 11832 -1902
rect 11752 -1922 11762 -1912
rect 11502 -1972 11762 -1922
rect 11822 -1972 11832 -1912
rect 11432 -1982 11832 -1972
rect 11890 -1562 12290 -1552
rect 11890 -1622 11900 -1562
rect 11960 -1612 12220 -1562
rect 11960 -1622 11970 -1612
rect 11890 -1632 11970 -1622
rect 12210 -1622 12220 -1612
rect 12280 -1622 12290 -1562
rect 12210 -1632 12290 -1622
rect 11890 -1902 11950 -1632
rect 12220 -1642 12290 -1632
rect 12030 -1692 12060 -1672
rect 12010 -1732 12060 -1692
rect 12120 -1692 12150 -1672
rect 12120 -1732 12170 -1692
rect 12010 -1802 12170 -1732
rect 12010 -1842 12060 -1802
rect 12030 -1862 12060 -1842
rect 12120 -1842 12170 -1802
rect 12120 -1862 12150 -1842
rect 12230 -1902 12290 -1642
rect 11890 -1912 11970 -1902
rect 11890 -1972 11900 -1912
rect 11960 -1922 11970 -1912
rect 12210 -1912 12290 -1902
rect 12210 -1922 12220 -1912
rect 11960 -1972 12220 -1922
rect 12280 -1972 12290 -1912
rect 11890 -1982 12290 -1972
rect 12346 -1562 12746 -1552
rect 12346 -1622 12356 -1562
rect 12416 -1612 12676 -1562
rect 12416 -1622 12426 -1612
rect 12346 -1632 12426 -1622
rect 12666 -1622 12676 -1612
rect 12736 -1622 12746 -1562
rect 12666 -1632 12746 -1622
rect 12346 -1902 12406 -1632
rect 12676 -1642 12746 -1632
rect 12486 -1692 12516 -1672
rect 12466 -1732 12516 -1692
rect 12576 -1692 12606 -1672
rect 12576 -1732 12626 -1692
rect 12466 -1802 12626 -1732
rect 12466 -1842 12516 -1802
rect 12486 -1862 12516 -1842
rect 12576 -1842 12626 -1802
rect 12576 -1862 12606 -1842
rect 12686 -1902 12746 -1642
rect 12346 -1912 12426 -1902
rect 12346 -1972 12356 -1912
rect 12416 -1922 12426 -1912
rect 12666 -1912 12746 -1902
rect 12666 -1922 12676 -1912
rect 12416 -1972 12676 -1922
rect 12736 -1972 12746 -1912
rect 12346 -1982 12746 -1972
rect 12802 -1562 13202 -1552
rect 12802 -1622 12812 -1562
rect 12872 -1612 13132 -1562
rect 12872 -1622 12882 -1612
rect 12802 -1632 12882 -1622
rect 13122 -1622 13132 -1612
rect 13192 -1622 13202 -1562
rect 13122 -1632 13202 -1622
rect 12802 -1902 12862 -1632
rect 13132 -1642 13202 -1632
rect 12942 -1692 12972 -1672
rect 12922 -1732 12972 -1692
rect 13032 -1692 13062 -1672
rect 13032 -1732 13082 -1692
rect 12922 -1802 13082 -1732
rect 12922 -1842 12972 -1802
rect 12942 -1862 12972 -1842
rect 13032 -1842 13082 -1802
rect 13032 -1862 13062 -1842
rect 13142 -1902 13202 -1642
rect 12802 -1912 12882 -1902
rect 12802 -1972 12812 -1912
rect 12872 -1922 12882 -1912
rect 13122 -1912 13202 -1902
rect 13122 -1922 13132 -1912
rect 12872 -1972 13132 -1922
rect 13192 -1972 13202 -1912
rect 12802 -1982 13202 -1972
rect 13260 -1562 13660 -1552
rect 13260 -1622 13270 -1562
rect 13330 -1612 13590 -1562
rect 13330 -1622 13340 -1612
rect 13260 -1632 13340 -1622
rect 13580 -1622 13590 -1612
rect 13650 -1622 13660 -1562
rect 13580 -1632 13660 -1622
rect 13260 -1902 13320 -1632
rect 13590 -1642 13660 -1632
rect 13400 -1692 13430 -1672
rect 13380 -1732 13430 -1692
rect 13490 -1692 13520 -1672
rect 13490 -1732 13540 -1692
rect 13380 -1802 13540 -1732
rect 13380 -1842 13430 -1802
rect 13400 -1862 13430 -1842
rect 13490 -1842 13540 -1802
rect 13490 -1862 13520 -1842
rect 13600 -1902 13660 -1642
rect 13260 -1912 13340 -1902
rect 13260 -1972 13270 -1912
rect 13330 -1922 13340 -1912
rect 13580 -1912 13660 -1902
rect 13580 -1922 13590 -1912
rect 13330 -1972 13590 -1922
rect 13650 -1972 13660 -1912
rect 13260 -1982 13660 -1972
rect 13716 -1562 14116 -1552
rect 13716 -1622 13726 -1562
rect 13786 -1612 14046 -1562
rect 13786 -1622 13796 -1612
rect 13716 -1632 13796 -1622
rect 14036 -1622 14046 -1612
rect 14106 -1622 14116 -1562
rect 14036 -1632 14116 -1622
rect 13716 -1902 13776 -1632
rect 14046 -1642 14116 -1632
rect 13856 -1692 13886 -1672
rect 13836 -1732 13886 -1692
rect 13946 -1692 13976 -1672
rect 13946 -1732 13996 -1692
rect 13836 -1802 13996 -1732
rect 13836 -1842 13886 -1802
rect 13856 -1862 13886 -1842
rect 13946 -1842 13996 -1802
rect 13946 -1862 13976 -1842
rect 14056 -1902 14116 -1642
rect 13716 -1912 13796 -1902
rect 13716 -1972 13726 -1912
rect 13786 -1922 13796 -1912
rect 14036 -1912 14116 -1902
rect 14036 -1922 14046 -1912
rect 13786 -1972 14046 -1922
rect 14106 -1972 14116 -1912
rect 13716 -1982 14116 -1972
rect 14172 -1562 14572 -1552
rect 14172 -1622 14182 -1562
rect 14242 -1612 14502 -1562
rect 14242 -1622 14252 -1612
rect 14172 -1632 14252 -1622
rect 14492 -1622 14502 -1612
rect 14562 -1622 14572 -1562
rect 14492 -1632 14572 -1622
rect 14172 -1902 14232 -1632
rect 14502 -1642 14572 -1632
rect 14312 -1692 14342 -1672
rect 14292 -1732 14342 -1692
rect 14402 -1692 14432 -1672
rect 14402 -1732 14452 -1692
rect 14292 -1802 14452 -1732
rect 14292 -1842 14342 -1802
rect 14312 -1862 14342 -1842
rect 14402 -1842 14452 -1802
rect 14402 -1862 14432 -1842
rect 14512 -1902 14572 -1642
rect 14172 -1912 14252 -1902
rect 14172 -1972 14182 -1912
rect 14242 -1922 14252 -1912
rect 14492 -1912 14572 -1902
rect 14492 -1922 14502 -1912
rect 14242 -1972 14502 -1922
rect 14562 -1972 14572 -1912
rect 14172 -1982 14572 -1972
rect 14630 -1562 15030 -1552
rect 14630 -1622 14640 -1562
rect 14700 -1612 14960 -1562
rect 14700 -1622 14710 -1612
rect 14630 -1632 14710 -1622
rect 14950 -1622 14960 -1612
rect 15020 -1622 15030 -1562
rect 14950 -1632 15030 -1622
rect 14630 -1902 14690 -1632
rect 14960 -1642 15030 -1632
rect 14770 -1692 14800 -1672
rect 14750 -1732 14800 -1692
rect 14860 -1692 14890 -1672
rect 14860 -1732 14910 -1692
rect 14750 -1802 14910 -1732
rect 14750 -1842 14800 -1802
rect 14770 -1862 14800 -1842
rect 14860 -1842 14910 -1802
rect 14860 -1862 14890 -1842
rect 14970 -1902 15030 -1642
rect 14630 -1912 14710 -1902
rect 14630 -1972 14640 -1912
rect 14700 -1922 14710 -1912
rect 14950 -1912 15030 -1902
rect 14950 -1922 14960 -1912
rect 14700 -1972 14960 -1922
rect 15020 -1972 15030 -1912
rect 14630 -1982 15030 -1972
rect 15086 -1562 15486 -1552
rect 15086 -1622 15096 -1562
rect 15156 -1612 15416 -1562
rect 15156 -1622 15166 -1612
rect 15086 -1632 15166 -1622
rect 15406 -1622 15416 -1612
rect 15476 -1622 15486 -1562
rect 15406 -1632 15486 -1622
rect 15086 -1902 15146 -1632
rect 15416 -1642 15486 -1632
rect 15226 -1692 15256 -1672
rect 15206 -1732 15256 -1692
rect 15316 -1692 15346 -1672
rect 15316 -1732 15366 -1692
rect 15206 -1802 15366 -1732
rect 15206 -1842 15256 -1802
rect 15226 -1862 15256 -1842
rect 15316 -1842 15366 -1802
rect 15316 -1862 15346 -1842
rect 15426 -1902 15486 -1642
rect 15086 -1912 15166 -1902
rect 15086 -1972 15096 -1912
rect 15156 -1922 15166 -1912
rect 15406 -1912 15486 -1902
rect 15406 -1922 15416 -1912
rect 15156 -1972 15416 -1922
rect 15476 -1972 15486 -1912
rect 15086 -1982 15486 -1972
rect 0 -2064 400 -2054
rect 0 -2124 10 -2064
rect 70 -2114 330 -2064
rect 70 -2124 80 -2114
rect 0 -2134 80 -2124
rect 320 -2124 330 -2114
rect 390 -2124 400 -2064
rect 320 -2134 400 -2124
rect 0 -2404 60 -2134
rect 330 -2144 400 -2134
rect 140 -2194 170 -2174
rect 120 -2234 170 -2194
rect 230 -2194 260 -2174
rect 230 -2234 280 -2194
rect 120 -2304 280 -2234
rect 120 -2344 170 -2304
rect 140 -2364 170 -2344
rect 230 -2344 280 -2304
rect 230 -2364 260 -2344
rect 340 -2404 400 -2144
rect 0 -2414 80 -2404
rect 0 -2474 10 -2414
rect 70 -2424 80 -2414
rect 320 -2414 400 -2404
rect 320 -2424 330 -2414
rect 70 -2474 330 -2424
rect 390 -2474 400 -2414
rect 0 -2484 400 -2474
rect 456 -2064 856 -2054
rect 456 -2124 466 -2064
rect 526 -2114 786 -2064
rect 526 -2124 536 -2114
rect 456 -2134 536 -2124
rect 776 -2124 786 -2114
rect 846 -2124 856 -2064
rect 776 -2134 856 -2124
rect 456 -2404 516 -2134
rect 786 -2144 856 -2134
rect 596 -2194 626 -2174
rect 576 -2234 626 -2194
rect 686 -2194 716 -2174
rect 686 -2234 736 -2194
rect 576 -2304 736 -2234
rect 576 -2344 626 -2304
rect 596 -2364 626 -2344
rect 686 -2344 736 -2304
rect 686 -2364 716 -2344
rect 796 -2404 856 -2144
rect 456 -2414 536 -2404
rect 456 -2474 466 -2414
rect 526 -2424 536 -2414
rect 776 -2414 856 -2404
rect 776 -2424 786 -2414
rect 526 -2474 786 -2424
rect 846 -2474 856 -2414
rect 456 -2484 856 -2474
rect 912 -2064 1312 -2054
rect 912 -2124 922 -2064
rect 982 -2114 1242 -2064
rect 982 -2124 992 -2114
rect 912 -2134 992 -2124
rect 1232 -2124 1242 -2114
rect 1302 -2124 1312 -2064
rect 1232 -2134 1312 -2124
rect 912 -2404 972 -2134
rect 1242 -2144 1312 -2134
rect 1052 -2194 1082 -2174
rect 1032 -2234 1082 -2194
rect 1142 -2194 1172 -2174
rect 1142 -2234 1192 -2194
rect 1032 -2304 1192 -2234
rect 1032 -2344 1082 -2304
rect 1052 -2364 1082 -2344
rect 1142 -2344 1192 -2304
rect 1142 -2364 1172 -2344
rect 1252 -2404 1312 -2144
rect 912 -2414 992 -2404
rect 912 -2474 922 -2414
rect 982 -2424 992 -2414
rect 1232 -2414 1312 -2404
rect 1232 -2424 1242 -2414
rect 982 -2474 1242 -2424
rect 1302 -2474 1312 -2414
rect 912 -2484 1312 -2474
rect 1370 -2064 1770 -2054
rect 1370 -2124 1380 -2064
rect 1440 -2114 1700 -2064
rect 1440 -2124 1450 -2114
rect 1370 -2134 1450 -2124
rect 1690 -2124 1700 -2114
rect 1760 -2124 1770 -2064
rect 1690 -2134 1770 -2124
rect 1370 -2404 1430 -2134
rect 1700 -2144 1770 -2134
rect 1510 -2194 1540 -2174
rect 1490 -2234 1540 -2194
rect 1600 -2194 1630 -2174
rect 1600 -2234 1650 -2194
rect 1490 -2304 1650 -2234
rect 1490 -2344 1540 -2304
rect 1510 -2364 1540 -2344
rect 1600 -2344 1650 -2304
rect 1600 -2364 1630 -2344
rect 1710 -2404 1770 -2144
rect 1370 -2414 1450 -2404
rect 1370 -2474 1380 -2414
rect 1440 -2424 1450 -2414
rect 1690 -2414 1770 -2404
rect 1690 -2424 1700 -2414
rect 1440 -2474 1700 -2424
rect 1760 -2474 1770 -2414
rect 1370 -2484 1770 -2474
rect 1826 -2064 2226 -2054
rect 1826 -2124 1836 -2064
rect 1896 -2114 2156 -2064
rect 1896 -2124 1906 -2114
rect 1826 -2134 1906 -2124
rect 2146 -2124 2156 -2114
rect 2216 -2124 2226 -2064
rect 2146 -2134 2226 -2124
rect 1826 -2404 1886 -2134
rect 2156 -2144 2226 -2134
rect 1966 -2194 1996 -2174
rect 1946 -2234 1996 -2194
rect 2056 -2194 2086 -2174
rect 2056 -2234 2106 -2194
rect 1946 -2304 2106 -2234
rect 1946 -2344 1996 -2304
rect 1966 -2364 1996 -2344
rect 2056 -2344 2106 -2304
rect 2056 -2364 2086 -2344
rect 2166 -2404 2226 -2144
rect 1826 -2414 1906 -2404
rect 1826 -2474 1836 -2414
rect 1896 -2424 1906 -2414
rect 2146 -2414 2226 -2404
rect 2146 -2424 2156 -2414
rect 1896 -2474 2156 -2424
rect 2216 -2474 2226 -2414
rect 1826 -2484 2226 -2474
rect 2282 -2064 2682 -2054
rect 2282 -2124 2292 -2064
rect 2352 -2114 2612 -2064
rect 2352 -2124 2362 -2114
rect 2282 -2134 2362 -2124
rect 2602 -2124 2612 -2114
rect 2672 -2124 2682 -2064
rect 2602 -2134 2682 -2124
rect 2282 -2404 2342 -2134
rect 2612 -2144 2682 -2134
rect 2422 -2194 2452 -2174
rect 2402 -2234 2452 -2194
rect 2512 -2194 2542 -2174
rect 2512 -2234 2562 -2194
rect 2402 -2304 2562 -2234
rect 2402 -2344 2452 -2304
rect 2422 -2364 2452 -2344
rect 2512 -2344 2562 -2304
rect 2512 -2364 2542 -2344
rect 2622 -2404 2682 -2144
rect 2282 -2414 2362 -2404
rect 2282 -2474 2292 -2414
rect 2352 -2424 2362 -2414
rect 2602 -2414 2682 -2404
rect 2602 -2424 2612 -2414
rect 2352 -2474 2612 -2424
rect 2672 -2474 2682 -2414
rect 2282 -2484 2682 -2474
rect 2740 -2064 3140 -2054
rect 2740 -2124 2750 -2064
rect 2810 -2114 3070 -2064
rect 2810 -2124 2820 -2114
rect 2740 -2134 2820 -2124
rect 3060 -2124 3070 -2114
rect 3130 -2124 3140 -2064
rect 3060 -2134 3140 -2124
rect 2740 -2404 2800 -2134
rect 3070 -2144 3140 -2134
rect 2880 -2194 2910 -2174
rect 2860 -2234 2910 -2194
rect 2970 -2194 3000 -2174
rect 2970 -2234 3020 -2194
rect 2860 -2304 3020 -2234
rect 2860 -2344 2910 -2304
rect 2880 -2364 2910 -2344
rect 2970 -2344 3020 -2304
rect 2970 -2364 3000 -2344
rect 3080 -2404 3140 -2144
rect 2740 -2414 2820 -2404
rect 2740 -2474 2750 -2414
rect 2810 -2424 2820 -2414
rect 3060 -2414 3140 -2404
rect 3060 -2424 3070 -2414
rect 2810 -2474 3070 -2424
rect 3130 -2474 3140 -2414
rect 2740 -2484 3140 -2474
rect 3196 -2064 3596 -2054
rect 3196 -2124 3206 -2064
rect 3266 -2114 3526 -2064
rect 3266 -2124 3276 -2114
rect 3196 -2134 3276 -2124
rect 3516 -2124 3526 -2114
rect 3586 -2124 3596 -2064
rect 3516 -2134 3596 -2124
rect 3196 -2404 3256 -2134
rect 3526 -2144 3596 -2134
rect 3336 -2194 3366 -2174
rect 3316 -2234 3366 -2194
rect 3426 -2194 3456 -2174
rect 3426 -2234 3476 -2194
rect 3316 -2304 3476 -2234
rect 3316 -2344 3366 -2304
rect 3336 -2364 3366 -2344
rect 3426 -2344 3476 -2304
rect 3426 -2364 3456 -2344
rect 3536 -2404 3596 -2144
rect 3196 -2414 3276 -2404
rect 3196 -2474 3206 -2414
rect 3266 -2424 3276 -2414
rect 3516 -2414 3596 -2404
rect 3516 -2424 3526 -2414
rect 3266 -2474 3526 -2424
rect 3586 -2474 3596 -2414
rect 3196 -2484 3596 -2474
rect 3652 -2064 4052 -2054
rect 3652 -2124 3662 -2064
rect 3722 -2114 3982 -2064
rect 3722 -2124 3732 -2114
rect 3652 -2134 3732 -2124
rect 3972 -2124 3982 -2114
rect 4042 -2124 4052 -2064
rect 3972 -2134 4052 -2124
rect 3652 -2404 3712 -2134
rect 3982 -2144 4052 -2134
rect 3792 -2194 3822 -2174
rect 3772 -2234 3822 -2194
rect 3882 -2194 3912 -2174
rect 3882 -2234 3932 -2194
rect 3772 -2304 3932 -2234
rect 3772 -2344 3822 -2304
rect 3792 -2364 3822 -2344
rect 3882 -2344 3932 -2304
rect 3882 -2364 3912 -2344
rect 3992 -2404 4052 -2144
rect 3652 -2414 3732 -2404
rect 3652 -2474 3662 -2414
rect 3722 -2424 3732 -2414
rect 3972 -2414 4052 -2404
rect 3972 -2424 3982 -2414
rect 3722 -2474 3982 -2424
rect 4042 -2474 4052 -2414
rect 3652 -2484 4052 -2474
rect 4110 -2064 4510 -2054
rect 4110 -2124 4120 -2064
rect 4180 -2114 4440 -2064
rect 4180 -2124 4190 -2114
rect 4110 -2134 4190 -2124
rect 4430 -2124 4440 -2114
rect 4500 -2124 4510 -2064
rect 4430 -2134 4510 -2124
rect 4110 -2404 4170 -2134
rect 4440 -2144 4510 -2134
rect 4250 -2194 4280 -2174
rect 4230 -2234 4280 -2194
rect 4340 -2194 4370 -2174
rect 4340 -2234 4390 -2194
rect 4230 -2304 4390 -2234
rect 4230 -2344 4280 -2304
rect 4250 -2364 4280 -2344
rect 4340 -2344 4390 -2304
rect 4340 -2364 4370 -2344
rect 4450 -2404 4510 -2144
rect 4110 -2414 4190 -2404
rect 4110 -2474 4120 -2414
rect 4180 -2424 4190 -2414
rect 4430 -2414 4510 -2404
rect 4430 -2424 4440 -2414
rect 4180 -2474 4440 -2424
rect 4500 -2474 4510 -2414
rect 4110 -2484 4510 -2474
rect 4566 -2064 4966 -2054
rect 4566 -2124 4576 -2064
rect 4636 -2114 4896 -2064
rect 4636 -2124 4646 -2114
rect 4566 -2134 4646 -2124
rect 4886 -2124 4896 -2114
rect 4956 -2124 4966 -2064
rect 4886 -2134 4966 -2124
rect 4566 -2404 4626 -2134
rect 4896 -2144 4966 -2134
rect 4706 -2194 4736 -2174
rect 4686 -2234 4736 -2194
rect 4796 -2194 4826 -2174
rect 4796 -2234 4846 -2194
rect 4686 -2304 4846 -2234
rect 4686 -2344 4736 -2304
rect 4706 -2364 4736 -2344
rect 4796 -2344 4846 -2304
rect 4796 -2364 4826 -2344
rect 4906 -2404 4966 -2144
rect 4566 -2414 4646 -2404
rect 4566 -2474 4576 -2414
rect 4636 -2424 4646 -2414
rect 4886 -2414 4966 -2404
rect 4886 -2424 4896 -2414
rect 4636 -2474 4896 -2424
rect 4956 -2474 4966 -2414
rect 4566 -2484 4966 -2474
rect 5022 -2064 5422 -2054
rect 5022 -2124 5032 -2064
rect 5092 -2114 5352 -2064
rect 5092 -2124 5102 -2114
rect 5022 -2134 5102 -2124
rect 5342 -2124 5352 -2114
rect 5412 -2124 5422 -2064
rect 5342 -2134 5422 -2124
rect 5022 -2404 5082 -2134
rect 5352 -2144 5422 -2134
rect 5162 -2194 5192 -2174
rect 5142 -2234 5192 -2194
rect 5252 -2194 5282 -2174
rect 5252 -2234 5302 -2194
rect 5142 -2304 5302 -2234
rect 5142 -2344 5192 -2304
rect 5162 -2364 5192 -2344
rect 5252 -2344 5302 -2304
rect 5252 -2364 5282 -2344
rect 5362 -2404 5422 -2144
rect 5022 -2414 5102 -2404
rect 5022 -2474 5032 -2414
rect 5092 -2424 5102 -2414
rect 5342 -2414 5422 -2404
rect 5342 -2424 5352 -2414
rect 5092 -2474 5352 -2424
rect 5412 -2474 5422 -2414
rect 5022 -2484 5422 -2474
rect 5480 -2064 5880 -2054
rect 5480 -2124 5490 -2064
rect 5550 -2114 5810 -2064
rect 5550 -2124 5560 -2114
rect 5480 -2134 5560 -2124
rect 5800 -2124 5810 -2114
rect 5870 -2124 5880 -2064
rect 5800 -2134 5880 -2124
rect 5480 -2404 5540 -2134
rect 5810 -2144 5880 -2134
rect 5620 -2194 5650 -2174
rect 5600 -2234 5650 -2194
rect 5710 -2194 5740 -2174
rect 5710 -2234 5760 -2194
rect 5600 -2304 5760 -2234
rect 5600 -2344 5650 -2304
rect 5620 -2364 5650 -2344
rect 5710 -2344 5760 -2304
rect 5710 -2364 5740 -2344
rect 5820 -2404 5880 -2144
rect 5480 -2414 5560 -2404
rect 5480 -2474 5490 -2414
rect 5550 -2424 5560 -2414
rect 5800 -2414 5880 -2404
rect 5800 -2424 5810 -2414
rect 5550 -2474 5810 -2424
rect 5870 -2474 5880 -2414
rect 5480 -2484 5880 -2474
rect 5936 -2064 6336 -2054
rect 5936 -2124 5946 -2064
rect 6006 -2114 6266 -2064
rect 6006 -2124 6016 -2114
rect 5936 -2134 6016 -2124
rect 6256 -2124 6266 -2114
rect 6326 -2124 6336 -2064
rect 6256 -2134 6336 -2124
rect 5936 -2404 5996 -2134
rect 6266 -2144 6336 -2134
rect 6076 -2194 6106 -2174
rect 6056 -2234 6106 -2194
rect 6166 -2194 6196 -2174
rect 6166 -2234 6216 -2194
rect 6056 -2304 6216 -2234
rect 6056 -2344 6106 -2304
rect 6076 -2364 6106 -2344
rect 6166 -2344 6216 -2304
rect 6166 -2364 6196 -2344
rect 6276 -2404 6336 -2144
rect 5936 -2414 6016 -2404
rect 5936 -2474 5946 -2414
rect 6006 -2424 6016 -2414
rect 6256 -2414 6336 -2404
rect 6256 -2424 6266 -2414
rect 6006 -2474 6266 -2424
rect 6326 -2474 6336 -2414
rect 5936 -2484 6336 -2474
rect 6392 -2064 6792 -2054
rect 6392 -2124 6402 -2064
rect 6462 -2114 6722 -2064
rect 6462 -2124 6472 -2114
rect 6392 -2134 6472 -2124
rect 6712 -2124 6722 -2114
rect 6782 -2124 6792 -2064
rect 6712 -2134 6792 -2124
rect 6392 -2404 6452 -2134
rect 6722 -2144 6792 -2134
rect 6532 -2194 6562 -2174
rect 6512 -2234 6562 -2194
rect 6622 -2194 6652 -2174
rect 6622 -2234 6672 -2194
rect 6512 -2304 6672 -2234
rect 6512 -2344 6562 -2304
rect 6532 -2364 6562 -2344
rect 6622 -2344 6672 -2304
rect 6622 -2364 6652 -2344
rect 6732 -2404 6792 -2144
rect 6392 -2414 6472 -2404
rect 6392 -2474 6402 -2414
rect 6462 -2424 6472 -2414
rect 6712 -2414 6792 -2404
rect 6712 -2424 6722 -2414
rect 6462 -2474 6722 -2424
rect 6782 -2474 6792 -2414
rect 6392 -2484 6792 -2474
rect 6850 -2064 7250 -2054
rect 6850 -2124 6860 -2064
rect 6920 -2114 7180 -2064
rect 6920 -2124 6930 -2114
rect 6850 -2134 6930 -2124
rect 7170 -2124 7180 -2114
rect 7240 -2124 7250 -2064
rect 7170 -2134 7250 -2124
rect 6850 -2404 6910 -2134
rect 7180 -2144 7250 -2134
rect 6990 -2194 7020 -2174
rect 6970 -2234 7020 -2194
rect 7080 -2194 7110 -2174
rect 7080 -2234 7130 -2194
rect 6970 -2304 7130 -2234
rect 6970 -2344 7020 -2304
rect 6990 -2364 7020 -2344
rect 7080 -2344 7130 -2304
rect 7080 -2364 7110 -2344
rect 7190 -2404 7250 -2144
rect 6850 -2414 6930 -2404
rect 6850 -2474 6860 -2414
rect 6920 -2424 6930 -2414
rect 7170 -2414 7250 -2404
rect 7170 -2424 7180 -2414
rect 6920 -2474 7180 -2424
rect 7240 -2474 7250 -2414
rect 6850 -2484 7250 -2474
rect 7306 -2064 7706 -2054
rect 7306 -2124 7316 -2064
rect 7376 -2114 7636 -2064
rect 7376 -2124 7386 -2114
rect 7306 -2134 7386 -2124
rect 7626 -2124 7636 -2114
rect 7696 -2124 7706 -2064
rect 7626 -2134 7706 -2124
rect 7306 -2404 7366 -2134
rect 7636 -2144 7706 -2134
rect 7446 -2194 7476 -2174
rect 7426 -2234 7476 -2194
rect 7536 -2194 7566 -2174
rect 7536 -2234 7586 -2194
rect 7426 -2304 7586 -2234
rect 7426 -2344 7476 -2304
rect 7446 -2364 7476 -2344
rect 7536 -2344 7586 -2304
rect 7536 -2364 7566 -2344
rect 7646 -2404 7706 -2144
rect 7306 -2414 7386 -2404
rect 7306 -2474 7316 -2414
rect 7376 -2424 7386 -2414
rect 7626 -2414 7706 -2404
rect 7626 -2424 7636 -2414
rect 7376 -2474 7636 -2424
rect 7696 -2474 7706 -2414
rect 7306 -2484 7706 -2474
rect 7762 -2064 8162 -2054
rect 7762 -2124 7772 -2064
rect 7832 -2114 8092 -2064
rect 7832 -2124 7842 -2114
rect 7762 -2134 7842 -2124
rect 8082 -2124 8092 -2114
rect 8152 -2124 8162 -2064
rect 8082 -2134 8162 -2124
rect 7762 -2404 7822 -2134
rect 8092 -2144 8162 -2134
rect 7902 -2194 7932 -2174
rect 7882 -2234 7932 -2194
rect 7992 -2194 8022 -2174
rect 7992 -2234 8042 -2194
rect 7882 -2304 8042 -2234
rect 7882 -2344 7932 -2304
rect 7902 -2364 7932 -2344
rect 7992 -2344 8042 -2304
rect 7992 -2364 8022 -2344
rect 8102 -2404 8162 -2144
rect 7762 -2414 7842 -2404
rect 7762 -2474 7772 -2414
rect 7832 -2424 7842 -2414
rect 8082 -2414 8162 -2404
rect 8082 -2424 8092 -2414
rect 7832 -2474 8092 -2424
rect 8152 -2474 8162 -2414
rect 7762 -2484 8162 -2474
rect 8236 -2064 8636 -2054
rect 8236 -2124 8246 -2064
rect 8306 -2114 8566 -2064
rect 8306 -2124 8316 -2114
rect 8236 -2134 8316 -2124
rect 8556 -2124 8566 -2114
rect 8626 -2124 8636 -2064
rect 8556 -2134 8636 -2124
rect 8236 -2404 8296 -2134
rect 8566 -2144 8636 -2134
rect 8376 -2194 8406 -2174
rect 8356 -2234 8406 -2194
rect 8466 -2194 8496 -2174
rect 8466 -2234 8516 -2194
rect 8356 -2304 8516 -2234
rect 8356 -2344 8406 -2304
rect 8376 -2364 8406 -2344
rect 8466 -2344 8516 -2304
rect 8466 -2364 8496 -2344
rect 8576 -2404 8636 -2144
rect 8236 -2414 8316 -2404
rect 8236 -2474 8246 -2414
rect 8306 -2424 8316 -2414
rect 8556 -2414 8636 -2404
rect 8556 -2424 8566 -2414
rect 8306 -2474 8566 -2424
rect 8626 -2474 8636 -2414
rect 8236 -2484 8636 -2474
rect 8692 -2064 9092 -2054
rect 8692 -2124 8702 -2064
rect 8762 -2114 9022 -2064
rect 8762 -2124 8772 -2114
rect 8692 -2134 8772 -2124
rect 9012 -2124 9022 -2114
rect 9082 -2124 9092 -2064
rect 9012 -2134 9092 -2124
rect 8692 -2404 8752 -2134
rect 9022 -2144 9092 -2134
rect 8832 -2194 8862 -2174
rect 8812 -2234 8862 -2194
rect 8922 -2194 8952 -2174
rect 8922 -2234 8972 -2194
rect 8812 -2304 8972 -2234
rect 8812 -2344 8862 -2304
rect 8832 -2364 8862 -2344
rect 8922 -2344 8972 -2304
rect 8922 -2364 8952 -2344
rect 9032 -2404 9092 -2144
rect 8692 -2414 8772 -2404
rect 8692 -2474 8702 -2414
rect 8762 -2424 8772 -2414
rect 9012 -2414 9092 -2404
rect 9012 -2424 9022 -2414
rect 8762 -2474 9022 -2424
rect 9082 -2474 9092 -2414
rect 8692 -2484 9092 -2474
rect 9150 -2064 9550 -2054
rect 9150 -2124 9160 -2064
rect 9220 -2114 9480 -2064
rect 9220 -2124 9230 -2114
rect 9150 -2134 9230 -2124
rect 9470 -2124 9480 -2114
rect 9540 -2124 9550 -2064
rect 9470 -2134 9550 -2124
rect 9150 -2404 9210 -2134
rect 9480 -2144 9550 -2134
rect 9290 -2194 9320 -2174
rect 9270 -2234 9320 -2194
rect 9380 -2194 9410 -2174
rect 9380 -2234 9430 -2194
rect 9270 -2304 9430 -2234
rect 9270 -2344 9320 -2304
rect 9290 -2364 9320 -2344
rect 9380 -2344 9430 -2304
rect 9380 -2364 9410 -2344
rect 9490 -2404 9550 -2144
rect 9150 -2414 9230 -2404
rect 9150 -2474 9160 -2414
rect 9220 -2424 9230 -2414
rect 9470 -2414 9550 -2404
rect 9470 -2424 9480 -2414
rect 9220 -2474 9480 -2424
rect 9540 -2474 9550 -2414
rect 9150 -2484 9550 -2474
rect 9606 -2064 10006 -2054
rect 9606 -2124 9616 -2064
rect 9676 -2114 9936 -2064
rect 9676 -2124 9686 -2114
rect 9606 -2134 9686 -2124
rect 9926 -2124 9936 -2114
rect 9996 -2124 10006 -2064
rect 9926 -2134 10006 -2124
rect 9606 -2404 9666 -2134
rect 9936 -2144 10006 -2134
rect 9746 -2194 9776 -2174
rect 9726 -2234 9776 -2194
rect 9836 -2194 9866 -2174
rect 9836 -2234 9886 -2194
rect 9726 -2304 9886 -2234
rect 9726 -2344 9776 -2304
rect 9746 -2364 9776 -2344
rect 9836 -2344 9886 -2304
rect 9836 -2364 9866 -2344
rect 9946 -2404 10006 -2144
rect 9606 -2414 9686 -2404
rect 9606 -2474 9616 -2414
rect 9676 -2424 9686 -2414
rect 9926 -2414 10006 -2404
rect 9926 -2424 9936 -2414
rect 9676 -2474 9936 -2424
rect 9996 -2474 10006 -2414
rect 9606 -2484 10006 -2474
rect 10062 -2064 10462 -2054
rect 10062 -2124 10072 -2064
rect 10132 -2114 10392 -2064
rect 10132 -2124 10142 -2114
rect 10062 -2134 10142 -2124
rect 10382 -2124 10392 -2114
rect 10452 -2124 10462 -2064
rect 10382 -2134 10462 -2124
rect 10062 -2404 10122 -2134
rect 10392 -2144 10462 -2134
rect 10202 -2194 10232 -2174
rect 10182 -2234 10232 -2194
rect 10292 -2194 10322 -2174
rect 10292 -2234 10342 -2194
rect 10182 -2304 10342 -2234
rect 10182 -2344 10232 -2304
rect 10202 -2364 10232 -2344
rect 10292 -2344 10342 -2304
rect 10292 -2364 10322 -2344
rect 10402 -2404 10462 -2144
rect 10062 -2414 10142 -2404
rect 10062 -2474 10072 -2414
rect 10132 -2424 10142 -2414
rect 10382 -2414 10462 -2404
rect 10382 -2424 10392 -2414
rect 10132 -2474 10392 -2424
rect 10452 -2474 10462 -2414
rect 10062 -2484 10462 -2474
rect 10520 -2064 10920 -2054
rect 10520 -2124 10530 -2064
rect 10590 -2114 10850 -2064
rect 10590 -2124 10600 -2114
rect 10520 -2134 10600 -2124
rect 10840 -2124 10850 -2114
rect 10910 -2124 10920 -2064
rect 10840 -2134 10920 -2124
rect 10520 -2404 10580 -2134
rect 10850 -2144 10920 -2134
rect 10660 -2194 10690 -2174
rect 10640 -2234 10690 -2194
rect 10750 -2194 10780 -2174
rect 10750 -2234 10800 -2194
rect 10640 -2304 10800 -2234
rect 10640 -2344 10690 -2304
rect 10660 -2364 10690 -2344
rect 10750 -2344 10800 -2304
rect 10750 -2364 10780 -2344
rect 10860 -2404 10920 -2144
rect 10520 -2414 10600 -2404
rect 10520 -2474 10530 -2414
rect 10590 -2424 10600 -2414
rect 10840 -2414 10920 -2404
rect 10840 -2424 10850 -2414
rect 10590 -2474 10850 -2424
rect 10910 -2474 10920 -2414
rect 10520 -2484 10920 -2474
rect 10976 -2064 11376 -2054
rect 10976 -2124 10986 -2064
rect 11046 -2114 11306 -2064
rect 11046 -2124 11056 -2114
rect 10976 -2134 11056 -2124
rect 11296 -2124 11306 -2114
rect 11366 -2124 11376 -2064
rect 11296 -2134 11376 -2124
rect 10976 -2404 11036 -2134
rect 11306 -2144 11376 -2134
rect 11116 -2194 11146 -2174
rect 11096 -2234 11146 -2194
rect 11206 -2194 11236 -2174
rect 11206 -2234 11256 -2194
rect 11096 -2304 11256 -2234
rect 11096 -2344 11146 -2304
rect 11116 -2364 11146 -2344
rect 11206 -2344 11256 -2304
rect 11206 -2364 11236 -2344
rect 11316 -2404 11376 -2144
rect 10976 -2414 11056 -2404
rect 10976 -2474 10986 -2414
rect 11046 -2424 11056 -2414
rect 11296 -2414 11376 -2404
rect 11296 -2424 11306 -2414
rect 11046 -2474 11306 -2424
rect 11366 -2474 11376 -2414
rect 10976 -2484 11376 -2474
rect 11432 -2064 11832 -2054
rect 11432 -2124 11442 -2064
rect 11502 -2114 11762 -2064
rect 11502 -2124 11512 -2114
rect 11432 -2134 11512 -2124
rect 11752 -2124 11762 -2114
rect 11822 -2124 11832 -2064
rect 11752 -2134 11832 -2124
rect 11432 -2404 11492 -2134
rect 11762 -2144 11832 -2134
rect 11572 -2194 11602 -2174
rect 11552 -2234 11602 -2194
rect 11662 -2194 11692 -2174
rect 11662 -2234 11712 -2194
rect 11552 -2304 11712 -2234
rect 11552 -2344 11602 -2304
rect 11572 -2364 11602 -2344
rect 11662 -2344 11712 -2304
rect 11662 -2364 11692 -2344
rect 11772 -2404 11832 -2144
rect 11432 -2414 11512 -2404
rect 11432 -2474 11442 -2414
rect 11502 -2424 11512 -2414
rect 11752 -2414 11832 -2404
rect 11752 -2424 11762 -2414
rect 11502 -2474 11762 -2424
rect 11822 -2474 11832 -2414
rect 11432 -2484 11832 -2474
rect 11890 -2064 12290 -2054
rect 11890 -2124 11900 -2064
rect 11960 -2114 12220 -2064
rect 11960 -2124 11970 -2114
rect 11890 -2134 11970 -2124
rect 12210 -2124 12220 -2114
rect 12280 -2124 12290 -2064
rect 12210 -2134 12290 -2124
rect 11890 -2404 11950 -2134
rect 12220 -2144 12290 -2134
rect 12030 -2194 12060 -2174
rect 12010 -2234 12060 -2194
rect 12120 -2194 12150 -2174
rect 12120 -2234 12170 -2194
rect 12010 -2304 12170 -2234
rect 12010 -2344 12060 -2304
rect 12030 -2364 12060 -2344
rect 12120 -2344 12170 -2304
rect 12120 -2364 12150 -2344
rect 12230 -2404 12290 -2144
rect 11890 -2414 11970 -2404
rect 11890 -2474 11900 -2414
rect 11960 -2424 11970 -2414
rect 12210 -2414 12290 -2404
rect 12210 -2424 12220 -2414
rect 11960 -2474 12220 -2424
rect 12280 -2474 12290 -2414
rect 11890 -2484 12290 -2474
rect 12346 -2064 12746 -2054
rect 12346 -2124 12356 -2064
rect 12416 -2114 12676 -2064
rect 12416 -2124 12426 -2114
rect 12346 -2134 12426 -2124
rect 12666 -2124 12676 -2114
rect 12736 -2124 12746 -2064
rect 12666 -2134 12746 -2124
rect 12346 -2404 12406 -2134
rect 12676 -2144 12746 -2134
rect 12486 -2194 12516 -2174
rect 12466 -2234 12516 -2194
rect 12576 -2194 12606 -2174
rect 12576 -2234 12626 -2194
rect 12466 -2304 12626 -2234
rect 12466 -2344 12516 -2304
rect 12486 -2364 12516 -2344
rect 12576 -2344 12626 -2304
rect 12576 -2364 12606 -2344
rect 12686 -2404 12746 -2144
rect 12346 -2414 12426 -2404
rect 12346 -2474 12356 -2414
rect 12416 -2424 12426 -2414
rect 12666 -2414 12746 -2404
rect 12666 -2424 12676 -2414
rect 12416 -2474 12676 -2424
rect 12736 -2474 12746 -2414
rect 12346 -2484 12746 -2474
rect 12802 -2064 13202 -2054
rect 12802 -2124 12812 -2064
rect 12872 -2114 13132 -2064
rect 12872 -2124 12882 -2114
rect 12802 -2134 12882 -2124
rect 13122 -2124 13132 -2114
rect 13192 -2124 13202 -2064
rect 13122 -2134 13202 -2124
rect 12802 -2404 12862 -2134
rect 13132 -2144 13202 -2134
rect 12942 -2194 12972 -2174
rect 12922 -2234 12972 -2194
rect 13032 -2194 13062 -2174
rect 13032 -2234 13082 -2194
rect 12922 -2304 13082 -2234
rect 12922 -2344 12972 -2304
rect 12942 -2364 12972 -2344
rect 13032 -2344 13082 -2304
rect 13032 -2364 13062 -2344
rect 13142 -2404 13202 -2144
rect 12802 -2414 12882 -2404
rect 12802 -2474 12812 -2414
rect 12872 -2424 12882 -2414
rect 13122 -2414 13202 -2404
rect 13122 -2424 13132 -2414
rect 12872 -2474 13132 -2424
rect 13192 -2474 13202 -2414
rect 12802 -2484 13202 -2474
rect 13260 -2064 13660 -2054
rect 13260 -2124 13270 -2064
rect 13330 -2114 13590 -2064
rect 13330 -2124 13340 -2114
rect 13260 -2134 13340 -2124
rect 13580 -2124 13590 -2114
rect 13650 -2124 13660 -2064
rect 13580 -2134 13660 -2124
rect 13260 -2404 13320 -2134
rect 13590 -2144 13660 -2134
rect 13400 -2194 13430 -2174
rect 13380 -2234 13430 -2194
rect 13490 -2194 13520 -2174
rect 13490 -2234 13540 -2194
rect 13380 -2304 13540 -2234
rect 13380 -2344 13430 -2304
rect 13400 -2364 13430 -2344
rect 13490 -2344 13540 -2304
rect 13490 -2364 13520 -2344
rect 13600 -2404 13660 -2144
rect 13260 -2414 13340 -2404
rect 13260 -2474 13270 -2414
rect 13330 -2424 13340 -2414
rect 13580 -2414 13660 -2404
rect 13580 -2424 13590 -2414
rect 13330 -2474 13590 -2424
rect 13650 -2474 13660 -2414
rect 13260 -2484 13660 -2474
rect 13716 -2064 14116 -2054
rect 13716 -2124 13726 -2064
rect 13786 -2114 14046 -2064
rect 13786 -2124 13796 -2114
rect 13716 -2134 13796 -2124
rect 14036 -2124 14046 -2114
rect 14106 -2124 14116 -2064
rect 14036 -2134 14116 -2124
rect 13716 -2404 13776 -2134
rect 14046 -2144 14116 -2134
rect 13856 -2194 13886 -2174
rect 13836 -2234 13886 -2194
rect 13946 -2194 13976 -2174
rect 13946 -2234 13996 -2194
rect 13836 -2304 13996 -2234
rect 13836 -2344 13886 -2304
rect 13856 -2364 13886 -2344
rect 13946 -2344 13996 -2304
rect 13946 -2364 13976 -2344
rect 14056 -2404 14116 -2144
rect 13716 -2414 13796 -2404
rect 13716 -2474 13726 -2414
rect 13786 -2424 13796 -2414
rect 14036 -2414 14116 -2404
rect 14036 -2424 14046 -2414
rect 13786 -2474 14046 -2424
rect 14106 -2474 14116 -2414
rect 13716 -2484 14116 -2474
rect 14172 -2064 14572 -2054
rect 14172 -2124 14182 -2064
rect 14242 -2114 14502 -2064
rect 14242 -2124 14252 -2114
rect 14172 -2134 14252 -2124
rect 14492 -2124 14502 -2114
rect 14562 -2124 14572 -2064
rect 14492 -2134 14572 -2124
rect 14172 -2404 14232 -2134
rect 14502 -2144 14572 -2134
rect 14312 -2194 14342 -2174
rect 14292 -2234 14342 -2194
rect 14402 -2194 14432 -2174
rect 14402 -2234 14452 -2194
rect 14292 -2304 14452 -2234
rect 14292 -2344 14342 -2304
rect 14312 -2364 14342 -2344
rect 14402 -2344 14452 -2304
rect 14402 -2364 14432 -2344
rect 14512 -2404 14572 -2144
rect 14172 -2414 14252 -2404
rect 14172 -2474 14182 -2414
rect 14242 -2424 14252 -2414
rect 14492 -2414 14572 -2404
rect 14492 -2424 14502 -2414
rect 14242 -2474 14502 -2424
rect 14562 -2474 14572 -2414
rect 14172 -2484 14572 -2474
rect 14630 -2064 15030 -2054
rect 14630 -2124 14640 -2064
rect 14700 -2114 14960 -2064
rect 14700 -2124 14710 -2114
rect 14630 -2134 14710 -2124
rect 14950 -2124 14960 -2114
rect 15020 -2124 15030 -2064
rect 14950 -2134 15030 -2124
rect 14630 -2404 14690 -2134
rect 14960 -2144 15030 -2134
rect 14770 -2194 14800 -2174
rect 14750 -2234 14800 -2194
rect 14860 -2194 14890 -2174
rect 14860 -2234 14910 -2194
rect 14750 -2304 14910 -2234
rect 14750 -2344 14800 -2304
rect 14770 -2364 14800 -2344
rect 14860 -2344 14910 -2304
rect 14860 -2364 14890 -2344
rect 14970 -2404 15030 -2144
rect 14630 -2414 14710 -2404
rect 14630 -2474 14640 -2414
rect 14700 -2424 14710 -2414
rect 14950 -2414 15030 -2404
rect 14950 -2424 14960 -2414
rect 14700 -2474 14960 -2424
rect 15020 -2474 15030 -2414
rect 14630 -2484 15030 -2474
rect 15086 -2064 15486 -2054
rect 15086 -2124 15096 -2064
rect 15156 -2114 15416 -2064
rect 15156 -2124 15166 -2114
rect 15086 -2134 15166 -2124
rect 15406 -2124 15416 -2114
rect 15476 -2124 15486 -2064
rect 15406 -2134 15486 -2124
rect 15086 -2404 15146 -2134
rect 15416 -2144 15486 -2134
rect 15226 -2194 15256 -2174
rect 15206 -2234 15256 -2194
rect 15316 -2194 15346 -2174
rect 15316 -2234 15366 -2194
rect 15206 -2304 15366 -2234
rect 15206 -2344 15256 -2304
rect 15226 -2364 15256 -2344
rect 15316 -2344 15366 -2304
rect 15316 -2364 15346 -2344
rect 15426 -2404 15486 -2144
rect 15086 -2414 15166 -2404
rect 15086 -2474 15096 -2414
rect 15156 -2424 15166 -2414
rect 15406 -2414 15486 -2404
rect 15406 -2424 15416 -2414
rect 15156 -2474 15416 -2424
rect 15476 -2474 15486 -2414
rect 15086 -2484 15486 -2474
rect 0 -2556 400 -2546
rect 0 -2616 10 -2556
rect 70 -2606 330 -2556
rect 70 -2616 80 -2606
rect 0 -2626 80 -2616
rect 320 -2616 330 -2606
rect 390 -2616 400 -2556
rect 320 -2626 400 -2616
rect 0 -2896 60 -2626
rect 330 -2636 400 -2626
rect 140 -2686 170 -2666
rect 120 -2726 170 -2686
rect 230 -2686 260 -2666
rect 230 -2726 280 -2686
rect 120 -2796 280 -2726
rect 120 -2836 170 -2796
rect 140 -2856 170 -2836
rect 230 -2836 280 -2796
rect 230 -2856 260 -2836
rect 340 -2896 400 -2636
rect 0 -2906 80 -2896
rect 0 -2966 10 -2906
rect 70 -2916 80 -2906
rect 320 -2906 400 -2896
rect 320 -2916 330 -2906
rect 70 -2966 330 -2916
rect 390 -2966 400 -2906
rect 0 -2976 400 -2966
rect 456 -2556 856 -2546
rect 456 -2616 466 -2556
rect 526 -2606 786 -2556
rect 526 -2616 536 -2606
rect 456 -2626 536 -2616
rect 776 -2616 786 -2606
rect 846 -2616 856 -2556
rect 776 -2626 856 -2616
rect 456 -2896 516 -2626
rect 786 -2636 856 -2626
rect 596 -2686 626 -2666
rect 576 -2726 626 -2686
rect 686 -2686 716 -2666
rect 686 -2726 736 -2686
rect 576 -2796 736 -2726
rect 576 -2836 626 -2796
rect 596 -2856 626 -2836
rect 686 -2836 736 -2796
rect 686 -2856 716 -2836
rect 796 -2896 856 -2636
rect 456 -2906 536 -2896
rect 456 -2966 466 -2906
rect 526 -2916 536 -2906
rect 776 -2906 856 -2896
rect 776 -2916 786 -2906
rect 526 -2966 786 -2916
rect 846 -2966 856 -2906
rect 456 -2976 856 -2966
rect 912 -2556 1312 -2546
rect 912 -2616 922 -2556
rect 982 -2606 1242 -2556
rect 982 -2616 992 -2606
rect 912 -2626 992 -2616
rect 1232 -2616 1242 -2606
rect 1302 -2616 1312 -2556
rect 1232 -2626 1312 -2616
rect 912 -2896 972 -2626
rect 1242 -2636 1312 -2626
rect 1052 -2686 1082 -2666
rect 1032 -2726 1082 -2686
rect 1142 -2686 1172 -2666
rect 1142 -2726 1192 -2686
rect 1032 -2796 1192 -2726
rect 1032 -2836 1082 -2796
rect 1052 -2856 1082 -2836
rect 1142 -2836 1192 -2796
rect 1142 -2856 1172 -2836
rect 1252 -2896 1312 -2636
rect 912 -2906 992 -2896
rect 912 -2966 922 -2906
rect 982 -2916 992 -2906
rect 1232 -2906 1312 -2896
rect 1232 -2916 1242 -2906
rect 982 -2966 1242 -2916
rect 1302 -2966 1312 -2906
rect 912 -2976 1312 -2966
rect 1370 -2556 1770 -2546
rect 1370 -2616 1380 -2556
rect 1440 -2606 1700 -2556
rect 1440 -2616 1450 -2606
rect 1370 -2626 1450 -2616
rect 1690 -2616 1700 -2606
rect 1760 -2616 1770 -2556
rect 1690 -2626 1770 -2616
rect 1370 -2896 1430 -2626
rect 1700 -2636 1770 -2626
rect 1510 -2686 1540 -2666
rect 1490 -2726 1540 -2686
rect 1600 -2686 1630 -2666
rect 1600 -2726 1650 -2686
rect 1490 -2796 1650 -2726
rect 1490 -2836 1540 -2796
rect 1510 -2856 1540 -2836
rect 1600 -2836 1650 -2796
rect 1600 -2856 1630 -2836
rect 1710 -2896 1770 -2636
rect 1370 -2906 1450 -2896
rect 1370 -2966 1380 -2906
rect 1440 -2916 1450 -2906
rect 1690 -2906 1770 -2896
rect 1690 -2916 1700 -2906
rect 1440 -2966 1700 -2916
rect 1760 -2966 1770 -2906
rect 1370 -2976 1770 -2966
rect 1826 -2556 2226 -2546
rect 1826 -2616 1836 -2556
rect 1896 -2606 2156 -2556
rect 1896 -2616 1906 -2606
rect 1826 -2626 1906 -2616
rect 2146 -2616 2156 -2606
rect 2216 -2616 2226 -2556
rect 2146 -2626 2226 -2616
rect 1826 -2896 1886 -2626
rect 2156 -2636 2226 -2626
rect 1966 -2686 1996 -2666
rect 1946 -2726 1996 -2686
rect 2056 -2686 2086 -2666
rect 2056 -2726 2106 -2686
rect 1946 -2796 2106 -2726
rect 1946 -2836 1996 -2796
rect 1966 -2856 1996 -2836
rect 2056 -2836 2106 -2796
rect 2056 -2856 2086 -2836
rect 2166 -2896 2226 -2636
rect 1826 -2906 1906 -2896
rect 1826 -2966 1836 -2906
rect 1896 -2916 1906 -2906
rect 2146 -2906 2226 -2896
rect 2146 -2916 2156 -2906
rect 1896 -2966 2156 -2916
rect 2216 -2966 2226 -2906
rect 1826 -2976 2226 -2966
rect 2282 -2556 2682 -2546
rect 2282 -2616 2292 -2556
rect 2352 -2606 2612 -2556
rect 2352 -2616 2362 -2606
rect 2282 -2626 2362 -2616
rect 2602 -2616 2612 -2606
rect 2672 -2616 2682 -2556
rect 2602 -2626 2682 -2616
rect 2282 -2896 2342 -2626
rect 2612 -2636 2682 -2626
rect 2422 -2686 2452 -2666
rect 2402 -2726 2452 -2686
rect 2512 -2686 2542 -2666
rect 2512 -2726 2562 -2686
rect 2402 -2796 2562 -2726
rect 2402 -2836 2452 -2796
rect 2422 -2856 2452 -2836
rect 2512 -2836 2562 -2796
rect 2512 -2856 2542 -2836
rect 2622 -2896 2682 -2636
rect 2282 -2906 2362 -2896
rect 2282 -2966 2292 -2906
rect 2352 -2916 2362 -2906
rect 2602 -2906 2682 -2896
rect 2602 -2916 2612 -2906
rect 2352 -2966 2612 -2916
rect 2672 -2966 2682 -2906
rect 2282 -2976 2682 -2966
rect 2740 -2556 3140 -2546
rect 2740 -2616 2750 -2556
rect 2810 -2606 3070 -2556
rect 2810 -2616 2820 -2606
rect 2740 -2626 2820 -2616
rect 3060 -2616 3070 -2606
rect 3130 -2616 3140 -2556
rect 3060 -2626 3140 -2616
rect 2740 -2896 2800 -2626
rect 3070 -2636 3140 -2626
rect 2880 -2686 2910 -2666
rect 2860 -2726 2910 -2686
rect 2970 -2686 3000 -2666
rect 2970 -2726 3020 -2686
rect 2860 -2796 3020 -2726
rect 2860 -2836 2910 -2796
rect 2880 -2856 2910 -2836
rect 2970 -2836 3020 -2796
rect 2970 -2856 3000 -2836
rect 3080 -2896 3140 -2636
rect 2740 -2906 2820 -2896
rect 2740 -2966 2750 -2906
rect 2810 -2916 2820 -2906
rect 3060 -2906 3140 -2896
rect 3060 -2916 3070 -2906
rect 2810 -2966 3070 -2916
rect 3130 -2966 3140 -2906
rect 2740 -2976 3140 -2966
rect 3196 -2556 3596 -2546
rect 3196 -2616 3206 -2556
rect 3266 -2606 3526 -2556
rect 3266 -2616 3276 -2606
rect 3196 -2626 3276 -2616
rect 3516 -2616 3526 -2606
rect 3586 -2616 3596 -2556
rect 3516 -2626 3596 -2616
rect 3196 -2896 3256 -2626
rect 3526 -2636 3596 -2626
rect 3336 -2686 3366 -2666
rect 3316 -2726 3366 -2686
rect 3426 -2686 3456 -2666
rect 3426 -2726 3476 -2686
rect 3316 -2796 3476 -2726
rect 3316 -2836 3366 -2796
rect 3336 -2856 3366 -2836
rect 3426 -2836 3476 -2796
rect 3426 -2856 3456 -2836
rect 3536 -2896 3596 -2636
rect 3196 -2906 3276 -2896
rect 3196 -2966 3206 -2906
rect 3266 -2916 3276 -2906
rect 3516 -2906 3596 -2896
rect 3516 -2916 3526 -2906
rect 3266 -2966 3526 -2916
rect 3586 -2966 3596 -2906
rect 3196 -2976 3596 -2966
rect 3652 -2556 4052 -2546
rect 3652 -2616 3662 -2556
rect 3722 -2606 3982 -2556
rect 3722 -2616 3732 -2606
rect 3652 -2626 3732 -2616
rect 3972 -2616 3982 -2606
rect 4042 -2616 4052 -2556
rect 3972 -2626 4052 -2616
rect 3652 -2896 3712 -2626
rect 3982 -2636 4052 -2626
rect 3792 -2686 3822 -2666
rect 3772 -2726 3822 -2686
rect 3882 -2686 3912 -2666
rect 3882 -2726 3932 -2686
rect 3772 -2796 3932 -2726
rect 3772 -2836 3822 -2796
rect 3792 -2856 3822 -2836
rect 3882 -2836 3932 -2796
rect 3882 -2856 3912 -2836
rect 3992 -2896 4052 -2636
rect 3652 -2906 3732 -2896
rect 3652 -2966 3662 -2906
rect 3722 -2916 3732 -2906
rect 3972 -2906 4052 -2896
rect 3972 -2916 3982 -2906
rect 3722 -2966 3982 -2916
rect 4042 -2966 4052 -2906
rect 3652 -2976 4052 -2966
rect 4110 -2556 4510 -2546
rect 4110 -2616 4120 -2556
rect 4180 -2606 4440 -2556
rect 4180 -2616 4190 -2606
rect 4110 -2626 4190 -2616
rect 4430 -2616 4440 -2606
rect 4500 -2616 4510 -2556
rect 4430 -2626 4510 -2616
rect 4110 -2896 4170 -2626
rect 4440 -2636 4510 -2626
rect 4250 -2686 4280 -2666
rect 4230 -2726 4280 -2686
rect 4340 -2686 4370 -2666
rect 4340 -2726 4390 -2686
rect 4230 -2796 4390 -2726
rect 4230 -2836 4280 -2796
rect 4250 -2856 4280 -2836
rect 4340 -2836 4390 -2796
rect 4340 -2856 4370 -2836
rect 4450 -2896 4510 -2636
rect 4110 -2906 4190 -2896
rect 4110 -2966 4120 -2906
rect 4180 -2916 4190 -2906
rect 4430 -2906 4510 -2896
rect 4430 -2916 4440 -2906
rect 4180 -2966 4440 -2916
rect 4500 -2966 4510 -2906
rect 4110 -2976 4510 -2966
rect 4566 -2556 4966 -2546
rect 4566 -2616 4576 -2556
rect 4636 -2606 4896 -2556
rect 4636 -2616 4646 -2606
rect 4566 -2626 4646 -2616
rect 4886 -2616 4896 -2606
rect 4956 -2616 4966 -2556
rect 4886 -2626 4966 -2616
rect 4566 -2896 4626 -2626
rect 4896 -2636 4966 -2626
rect 4706 -2686 4736 -2666
rect 4686 -2726 4736 -2686
rect 4796 -2686 4826 -2666
rect 4796 -2726 4846 -2686
rect 4686 -2796 4846 -2726
rect 4686 -2836 4736 -2796
rect 4706 -2856 4736 -2836
rect 4796 -2836 4846 -2796
rect 4796 -2856 4826 -2836
rect 4906 -2896 4966 -2636
rect 4566 -2906 4646 -2896
rect 4566 -2966 4576 -2906
rect 4636 -2916 4646 -2906
rect 4886 -2906 4966 -2896
rect 4886 -2916 4896 -2906
rect 4636 -2966 4896 -2916
rect 4956 -2966 4966 -2906
rect 4566 -2976 4966 -2966
rect 5022 -2556 5422 -2546
rect 5022 -2616 5032 -2556
rect 5092 -2606 5352 -2556
rect 5092 -2616 5102 -2606
rect 5022 -2626 5102 -2616
rect 5342 -2616 5352 -2606
rect 5412 -2616 5422 -2556
rect 5342 -2626 5422 -2616
rect 5022 -2896 5082 -2626
rect 5352 -2636 5422 -2626
rect 5162 -2686 5192 -2666
rect 5142 -2726 5192 -2686
rect 5252 -2686 5282 -2666
rect 5252 -2726 5302 -2686
rect 5142 -2796 5302 -2726
rect 5142 -2836 5192 -2796
rect 5162 -2856 5192 -2836
rect 5252 -2836 5302 -2796
rect 5252 -2856 5282 -2836
rect 5362 -2896 5422 -2636
rect 5022 -2906 5102 -2896
rect 5022 -2966 5032 -2906
rect 5092 -2916 5102 -2906
rect 5342 -2906 5422 -2896
rect 5342 -2916 5352 -2906
rect 5092 -2966 5352 -2916
rect 5412 -2966 5422 -2906
rect 5022 -2976 5422 -2966
rect 5480 -2556 5880 -2546
rect 5480 -2616 5490 -2556
rect 5550 -2606 5810 -2556
rect 5550 -2616 5560 -2606
rect 5480 -2626 5560 -2616
rect 5800 -2616 5810 -2606
rect 5870 -2616 5880 -2556
rect 5800 -2626 5880 -2616
rect 5480 -2896 5540 -2626
rect 5810 -2636 5880 -2626
rect 5620 -2686 5650 -2666
rect 5600 -2726 5650 -2686
rect 5710 -2686 5740 -2666
rect 5710 -2726 5760 -2686
rect 5600 -2796 5760 -2726
rect 5600 -2836 5650 -2796
rect 5620 -2856 5650 -2836
rect 5710 -2836 5760 -2796
rect 5710 -2856 5740 -2836
rect 5820 -2896 5880 -2636
rect 5480 -2906 5560 -2896
rect 5480 -2966 5490 -2906
rect 5550 -2916 5560 -2906
rect 5800 -2906 5880 -2896
rect 5800 -2916 5810 -2906
rect 5550 -2966 5810 -2916
rect 5870 -2966 5880 -2906
rect 5480 -2976 5880 -2966
rect 5936 -2556 6336 -2546
rect 5936 -2616 5946 -2556
rect 6006 -2606 6266 -2556
rect 6006 -2616 6016 -2606
rect 5936 -2626 6016 -2616
rect 6256 -2616 6266 -2606
rect 6326 -2616 6336 -2556
rect 6256 -2626 6336 -2616
rect 5936 -2896 5996 -2626
rect 6266 -2636 6336 -2626
rect 6076 -2686 6106 -2666
rect 6056 -2726 6106 -2686
rect 6166 -2686 6196 -2666
rect 6166 -2726 6216 -2686
rect 6056 -2796 6216 -2726
rect 6056 -2836 6106 -2796
rect 6076 -2856 6106 -2836
rect 6166 -2836 6216 -2796
rect 6166 -2856 6196 -2836
rect 6276 -2896 6336 -2636
rect 5936 -2906 6016 -2896
rect 5936 -2966 5946 -2906
rect 6006 -2916 6016 -2906
rect 6256 -2906 6336 -2896
rect 6256 -2916 6266 -2906
rect 6006 -2966 6266 -2916
rect 6326 -2966 6336 -2906
rect 5936 -2976 6336 -2966
rect 6392 -2556 6792 -2546
rect 6392 -2616 6402 -2556
rect 6462 -2606 6722 -2556
rect 6462 -2616 6472 -2606
rect 6392 -2626 6472 -2616
rect 6712 -2616 6722 -2606
rect 6782 -2616 6792 -2556
rect 6712 -2626 6792 -2616
rect 6392 -2896 6452 -2626
rect 6722 -2636 6792 -2626
rect 6532 -2686 6562 -2666
rect 6512 -2726 6562 -2686
rect 6622 -2686 6652 -2666
rect 6622 -2726 6672 -2686
rect 6512 -2796 6672 -2726
rect 6512 -2836 6562 -2796
rect 6532 -2856 6562 -2836
rect 6622 -2836 6672 -2796
rect 6622 -2856 6652 -2836
rect 6732 -2896 6792 -2636
rect 6392 -2906 6472 -2896
rect 6392 -2966 6402 -2906
rect 6462 -2916 6472 -2906
rect 6712 -2906 6792 -2896
rect 6712 -2916 6722 -2906
rect 6462 -2966 6722 -2916
rect 6782 -2966 6792 -2906
rect 6392 -2976 6792 -2966
rect 6850 -2556 7250 -2546
rect 6850 -2616 6860 -2556
rect 6920 -2606 7180 -2556
rect 6920 -2616 6930 -2606
rect 6850 -2626 6930 -2616
rect 7170 -2616 7180 -2606
rect 7240 -2616 7250 -2556
rect 7170 -2626 7250 -2616
rect 6850 -2896 6910 -2626
rect 7180 -2636 7250 -2626
rect 6990 -2686 7020 -2666
rect 6970 -2726 7020 -2686
rect 7080 -2686 7110 -2666
rect 7080 -2726 7130 -2686
rect 6970 -2796 7130 -2726
rect 6970 -2836 7020 -2796
rect 6990 -2856 7020 -2836
rect 7080 -2836 7130 -2796
rect 7080 -2856 7110 -2836
rect 7190 -2896 7250 -2636
rect 6850 -2906 6930 -2896
rect 6850 -2966 6860 -2906
rect 6920 -2916 6930 -2906
rect 7170 -2906 7250 -2896
rect 7170 -2916 7180 -2906
rect 6920 -2966 7180 -2916
rect 7240 -2966 7250 -2906
rect 6850 -2976 7250 -2966
rect 7306 -2556 7706 -2546
rect 7306 -2616 7316 -2556
rect 7376 -2606 7636 -2556
rect 7376 -2616 7386 -2606
rect 7306 -2626 7386 -2616
rect 7626 -2616 7636 -2606
rect 7696 -2616 7706 -2556
rect 7626 -2626 7706 -2616
rect 7306 -2896 7366 -2626
rect 7636 -2636 7706 -2626
rect 7446 -2686 7476 -2666
rect 7426 -2726 7476 -2686
rect 7536 -2686 7566 -2666
rect 7536 -2726 7586 -2686
rect 7426 -2796 7586 -2726
rect 7426 -2836 7476 -2796
rect 7446 -2856 7476 -2836
rect 7536 -2836 7586 -2796
rect 7536 -2856 7566 -2836
rect 7646 -2896 7706 -2636
rect 7306 -2906 7386 -2896
rect 7306 -2966 7316 -2906
rect 7376 -2916 7386 -2906
rect 7626 -2906 7706 -2896
rect 7626 -2916 7636 -2906
rect 7376 -2966 7636 -2916
rect 7696 -2966 7706 -2906
rect 7306 -2976 7706 -2966
rect 7762 -2556 8162 -2546
rect 7762 -2616 7772 -2556
rect 7832 -2606 8092 -2556
rect 7832 -2616 7842 -2606
rect 7762 -2626 7842 -2616
rect 8082 -2616 8092 -2606
rect 8152 -2616 8162 -2556
rect 8082 -2626 8162 -2616
rect 7762 -2896 7822 -2626
rect 8092 -2636 8162 -2626
rect 7902 -2686 7932 -2666
rect 7882 -2726 7932 -2686
rect 7992 -2686 8022 -2666
rect 7992 -2726 8042 -2686
rect 7882 -2796 8042 -2726
rect 7882 -2836 7932 -2796
rect 7902 -2856 7932 -2836
rect 7992 -2836 8042 -2796
rect 7992 -2856 8022 -2836
rect 8102 -2896 8162 -2636
rect 7762 -2906 7842 -2896
rect 7762 -2966 7772 -2906
rect 7832 -2916 7842 -2906
rect 8082 -2906 8162 -2896
rect 8082 -2916 8092 -2906
rect 7832 -2966 8092 -2916
rect 8152 -2966 8162 -2906
rect 7762 -2976 8162 -2966
rect 8236 -2556 8636 -2546
rect 8236 -2616 8246 -2556
rect 8306 -2606 8566 -2556
rect 8306 -2616 8316 -2606
rect 8236 -2626 8316 -2616
rect 8556 -2616 8566 -2606
rect 8626 -2616 8636 -2556
rect 8556 -2626 8636 -2616
rect 8236 -2896 8296 -2626
rect 8566 -2636 8636 -2626
rect 8376 -2686 8406 -2666
rect 8356 -2726 8406 -2686
rect 8466 -2686 8496 -2666
rect 8466 -2726 8516 -2686
rect 8356 -2796 8516 -2726
rect 8356 -2836 8406 -2796
rect 8376 -2856 8406 -2836
rect 8466 -2836 8516 -2796
rect 8466 -2856 8496 -2836
rect 8576 -2896 8636 -2636
rect 8236 -2906 8316 -2896
rect 8236 -2966 8246 -2906
rect 8306 -2916 8316 -2906
rect 8556 -2906 8636 -2896
rect 8556 -2916 8566 -2906
rect 8306 -2966 8566 -2916
rect 8626 -2966 8636 -2906
rect 8236 -2976 8636 -2966
rect 8692 -2556 9092 -2546
rect 8692 -2616 8702 -2556
rect 8762 -2606 9022 -2556
rect 8762 -2616 8772 -2606
rect 8692 -2626 8772 -2616
rect 9012 -2616 9022 -2606
rect 9082 -2616 9092 -2556
rect 9012 -2626 9092 -2616
rect 8692 -2896 8752 -2626
rect 9022 -2636 9092 -2626
rect 8832 -2686 8862 -2666
rect 8812 -2726 8862 -2686
rect 8922 -2686 8952 -2666
rect 8922 -2726 8972 -2686
rect 8812 -2796 8972 -2726
rect 8812 -2836 8862 -2796
rect 8832 -2856 8862 -2836
rect 8922 -2836 8972 -2796
rect 8922 -2856 8952 -2836
rect 9032 -2896 9092 -2636
rect 8692 -2906 8772 -2896
rect 8692 -2966 8702 -2906
rect 8762 -2916 8772 -2906
rect 9012 -2906 9092 -2896
rect 9012 -2916 9022 -2906
rect 8762 -2966 9022 -2916
rect 9082 -2966 9092 -2906
rect 8692 -2976 9092 -2966
rect 9150 -2556 9550 -2546
rect 9150 -2616 9160 -2556
rect 9220 -2606 9480 -2556
rect 9220 -2616 9230 -2606
rect 9150 -2626 9230 -2616
rect 9470 -2616 9480 -2606
rect 9540 -2616 9550 -2556
rect 9470 -2626 9550 -2616
rect 9150 -2896 9210 -2626
rect 9480 -2636 9550 -2626
rect 9290 -2686 9320 -2666
rect 9270 -2726 9320 -2686
rect 9380 -2686 9410 -2666
rect 9380 -2726 9430 -2686
rect 9270 -2796 9430 -2726
rect 9270 -2836 9320 -2796
rect 9290 -2856 9320 -2836
rect 9380 -2836 9430 -2796
rect 9380 -2856 9410 -2836
rect 9490 -2896 9550 -2636
rect 9150 -2906 9230 -2896
rect 9150 -2966 9160 -2906
rect 9220 -2916 9230 -2906
rect 9470 -2906 9550 -2896
rect 9470 -2916 9480 -2906
rect 9220 -2966 9480 -2916
rect 9540 -2966 9550 -2906
rect 9150 -2976 9550 -2966
rect 9606 -2556 10006 -2546
rect 9606 -2616 9616 -2556
rect 9676 -2606 9936 -2556
rect 9676 -2616 9686 -2606
rect 9606 -2626 9686 -2616
rect 9926 -2616 9936 -2606
rect 9996 -2616 10006 -2556
rect 9926 -2626 10006 -2616
rect 9606 -2896 9666 -2626
rect 9936 -2636 10006 -2626
rect 9746 -2686 9776 -2666
rect 9726 -2726 9776 -2686
rect 9836 -2686 9866 -2666
rect 9836 -2726 9886 -2686
rect 9726 -2796 9886 -2726
rect 9726 -2836 9776 -2796
rect 9746 -2856 9776 -2836
rect 9836 -2836 9886 -2796
rect 9836 -2856 9866 -2836
rect 9946 -2896 10006 -2636
rect 9606 -2906 9686 -2896
rect 9606 -2966 9616 -2906
rect 9676 -2916 9686 -2906
rect 9926 -2906 10006 -2896
rect 9926 -2916 9936 -2906
rect 9676 -2966 9936 -2916
rect 9996 -2966 10006 -2906
rect 9606 -2976 10006 -2966
rect 10062 -2556 10462 -2546
rect 10062 -2616 10072 -2556
rect 10132 -2606 10392 -2556
rect 10132 -2616 10142 -2606
rect 10062 -2626 10142 -2616
rect 10382 -2616 10392 -2606
rect 10452 -2616 10462 -2556
rect 10382 -2626 10462 -2616
rect 10062 -2896 10122 -2626
rect 10392 -2636 10462 -2626
rect 10202 -2686 10232 -2666
rect 10182 -2726 10232 -2686
rect 10292 -2686 10322 -2666
rect 10292 -2726 10342 -2686
rect 10182 -2796 10342 -2726
rect 10182 -2836 10232 -2796
rect 10202 -2856 10232 -2836
rect 10292 -2836 10342 -2796
rect 10292 -2856 10322 -2836
rect 10402 -2896 10462 -2636
rect 10062 -2906 10142 -2896
rect 10062 -2966 10072 -2906
rect 10132 -2916 10142 -2906
rect 10382 -2906 10462 -2896
rect 10382 -2916 10392 -2906
rect 10132 -2966 10392 -2916
rect 10452 -2966 10462 -2906
rect 10062 -2976 10462 -2966
rect 10520 -2556 10920 -2546
rect 10520 -2616 10530 -2556
rect 10590 -2606 10850 -2556
rect 10590 -2616 10600 -2606
rect 10520 -2626 10600 -2616
rect 10840 -2616 10850 -2606
rect 10910 -2616 10920 -2556
rect 10840 -2626 10920 -2616
rect 10520 -2896 10580 -2626
rect 10850 -2636 10920 -2626
rect 10660 -2686 10690 -2666
rect 10640 -2726 10690 -2686
rect 10750 -2686 10780 -2666
rect 10750 -2726 10800 -2686
rect 10640 -2796 10800 -2726
rect 10640 -2836 10690 -2796
rect 10660 -2856 10690 -2836
rect 10750 -2836 10800 -2796
rect 10750 -2856 10780 -2836
rect 10860 -2896 10920 -2636
rect 10520 -2906 10600 -2896
rect 10520 -2966 10530 -2906
rect 10590 -2916 10600 -2906
rect 10840 -2906 10920 -2896
rect 10840 -2916 10850 -2906
rect 10590 -2966 10850 -2916
rect 10910 -2966 10920 -2906
rect 10520 -2976 10920 -2966
rect 10976 -2556 11376 -2546
rect 10976 -2616 10986 -2556
rect 11046 -2606 11306 -2556
rect 11046 -2616 11056 -2606
rect 10976 -2626 11056 -2616
rect 11296 -2616 11306 -2606
rect 11366 -2616 11376 -2556
rect 11296 -2626 11376 -2616
rect 10976 -2896 11036 -2626
rect 11306 -2636 11376 -2626
rect 11116 -2686 11146 -2666
rect 11096 -2726 11146 -2686
rect 11206 -2686 11236 -2666
rect 11206 -2726 11256 -2686
rect 11096 -2796 11256 -2726
rect 11096 -2836 11146 -2796
rect 11116 -2856 11146 -2836
rect 11206 -2836 11256 -2796
rect 11206 -2856 11236 -2836
rect 11316 -2896 11376 -2636
rect 10976 -2906 11056 -2896
rect 10976 -2966 10986 -2906
rect 11046 -2916 11056 -2906
rect 11296 -2906 11376 -2896
rect 11296 -2916 11306 -2906
rect 11046 -2966 11306 -2916
rect 11366 -2966 11376 -2906
rect 10976 -2976 11376 -2966
rect 11432 -2556 11832 -2546
rect 11432 -2616 11442 -2556
rect 11502 -2606 11762 -2556
rect 11502 -2616 11512 -2606
rect 11432 -2626 11512 -2616
rect 11752 -2616 11762 -2606
rect 11822 -2616 11832 -2556
rect 11752 -2626 11832 -2616
rect 11432 -2896 11492 -2626
rect 11762 -2636 11832 -2626
rect 11572 -2686 11602 -2666
rect 11552 -2726 11602 -2686
rect 11662 -2686 11692 -2666
rect 11662 -2726 11712 -2686
rect 11552 -2796 11712 -2726
rect 11552 -2836 11602 -2796
rect 11572 -2856 11602 -2836
rect 11662 -2836 11712 -2796
rect 11662 -2856 11692 -2836
rect 11772 -2896 11832 -2636
rect 11432 -2906 11512 -2896
rect 11432 -2966 11442 -2906
rect 11502 -2916 11512 -2906
rect 11752 -2906 11832 -2896
rect 11752 -2916 11762 -2906
rect 11502 -2966 11762 -2916
rect 11822 -2966 11832 -2906
rect 11432 -2976 11832 -2966
rect 11890 -2556 12290 -2546
rect 11890 -2616 11900 -2556
rect 11960 -2606 12220 -2556
rect 11960 -2616 11970 -2606
rect 11890 -2626 11970 -2616
rect 12210 -2616 12220 -2606
rect 12280 -2616 12290 -2556
rect 12210 -2626 12290 -2616
rect 11890 -2896 11950 -2626
rect 12220 -2636 12290 -2626
rect 12030 -2686 12060 -2666
rect 12010 -2726 12060 -2686
rect 12120 -2686 12150 -2666
rect 12120 -2726 12170 -2686
rect 12010 -2796 12170 -2726
rect 12010 -2836 12060 -2796
rect 12030 -2856 12060 -2836
rect 12120 -2836 12170 -2796
rect 12120 -2856 12150 -2836
rect 12230 -2896 12290 -2636
rect 11890 -2906 11970 -2896
rect 11890 -2966 11900 -2906
rect 11960 -2916 11970 -2906
rect 12210 -2906 12290 -2896
rect 12210 -2916 12220 -2906
rect 11960 -2966 12220 -2916
rect 12280 -2966 12290 -2906
rect 11890 -2976 12290 -2966
rect 12346 -2556 12746 -2546
rect 12346 -2616 12356 -2556
rect 12416 -2606 12676 -2556
rect 12416 -2616 12426 -2606
rect 12346 -2626 12426 -2616
rect 12666 -2616 12676 -2606
rect 12736 -2616 12746 -2556
rect 12666 -2626 12746 -2616
rect 12346 -2896 12406 -2626
rect 12676 -2636 12746 -2626
rect 12486 -2686 12516 -2666
rect 12466 -2726 12516 -2686
rect 12576 -2686 12606 -2666
rect 12576 -2726 12626 -2686
rect 12466 -2796 12626 -2726
rect 12466 -2836 12516 -2796
rect 12486 -2856 12516 -2836
rect 12576 -2836 12626 -2796
rect 12576 -2856 12606 -2836
rect 12686 -2896 12746 -2636
rect 12346 -2906 12426 -2896
rect 12346 -2966 12356 -2906
rect 12416 -2916 12426 -2906
rect 12666 -2906 12746 -2896
rect 12666 -2916 12676 -2906
rect 12416 -2966 12676 -2916
rect 12736 -2966 12746 -2906
rect 12346 -2976 12746 -2966
rect 12802 -2556 13202 -2546
rect 12802 -2616 12812 -2556
rect 12872 -2606 13132 -2556
rect 12872 -2616 12882 -2606
rect 12802 -2626 12882 -2616
rect 13122 -2616 13132 -2606
rect 13192 -2616 13202 -2556
rect 13122 -2626 13202 -2616
rect 12802 -2896 12862 -2626
rect 13132 -2636 13202 -2626
rect 12942 -2686 12972 -2666
rect 12922 -2726 12972 -2686
rect 13032 -2686 13062 -2666
rect 13032 -2726 13082 -2686
rect 12922 -2796 13082 -2726
rect 12922 -2836 12972 -2796
rect 12942 -2856 12972 -2836
rect 13032 -2836 13082 -2796
rect 13032 -2856 13062 -2836
rect 13142 -2896 13202 -2636
rect 12802 -2906 12882 -2896
rect 12802 -2966 12812 -2906
rect 12872 -2916 12882 -2906
rect 13122 -2906 13202 -2896
rect 13122 -2916 13132 -2906
rect 12872 -2966 13132 -2916
rect 13192 -2966 13202 -2906
rect 12802 -2976 13202 -2966
rect 13260 -2556 13660 -2546
rect 13260 -2616 13270 -2556
rect 13330 -2606 13590 -2556
rect 13330 -2616 13340 -2606
rect 13260 -2626 13340 -2616
rect 13580 -2616 13590 -2606
rect 13650 -2616 13660 -2556
rect 13580 -2626 13660 -2616
rect 13260 -2896 13320 -2626
rect 13590 -2636 13660 -2626
rect 13400 -2686 13430 -2666
rect 13380 -2726 13430 -2686
rect 13490 -2686 13520 -2666
rect 13490 -2726 13540 -2686
rect 13380 -2796 13540 -2726
rect 13380 -2836 13430 -2796
rect 13400 -2856 13430 -2836
rect 13490 -2836 13540 -2796
rect 13490 -2856 13520 -2836
rect 13600 -2896 13660 -2636
rect 13260 -2906 13340 -2896
rect 13260 -2966 13270 -2906
rect 13330 -2916 13340 -2906
rect 13580 -2906 13660 -2896
rect 13580 -2916 13590 -2906
rect 13330 -2966 13590 -2916
rect 13650 -2966 13660 -2906
rect 13260 -2976 13660 -2966
rect 13716 -2556 14116 -2546
rect 13716 -2616 13726 -2556
rect 13786 -2606 14046 -2556
rect 13786 -2616 13796 -2606
rect 13716 -2626 13796 -2616
rect 14036 -2616 14046 -2606
rect 14106 -2616 14116 -2556
rect 14036 -2626 14116 -2616
rect 13716 -2896 13776 -2626
rect 14046 -2636 14116 -2626
rect 13856 -2686 13886 -2666
rect 13836 -2726 13886 -2686
rect 13946 -2686 13976 -2666
rect 13946 -2726 13996 -2686
rect 13836 -2796 13996 -2726
rect 13836 -2836 13886 -2796
rect 13856 -2856 13886 -2836
rect 13946 -2836 13996 -2796
rect 13946 -2856 13976 -2836
rect 14056 -2896 14116 -2636
rect 13716 -2906 13796 -2896
rect 13716 -2966 13726 -2906
rect 13786 -2916 13796 -2906
rect 14036 -2906 14116 -2896
rect 14036 -2916 14046 -2906
rect 13786 -2966 14046 -2916
rect 14106 -2966 14116 -2906
rect 13716 -2976 14116 -2966
rect 14172 -2556 14572 -2546
rect 14172 -2616 14182 -2556
rect 14242 -2606 14502 -2556
rect 14242 -2616 14252 -2606
rect 14172 -2626 14252 -2616
rect 14492 -2616 14502 -2606
rect 14562 -2616 14572 -2556
rect 14492 -2626 14572 -2616
rect 14172 -2896 14232 -2626
rect 14502 -2636 14572 -2626
rect 14312 -2686 14342 -2666
rect 14292 -2726 14342 -2686
rect 14402 -2686 14432 -2666
rect 14402 -2726 14452 -2686
rect 14292 -2796 14452 -2726
rect 14292 -2836 14342 -2796
rect 14312 -2856 14342 -2836
rect 14402 -2836 14452 -2796
rect 14402 -2856 14432 -2836
rect 14512 -2896 14572 -2636
rect 14172 -2906 14252 -2896
rect 14172 -2966 14182 -2906
rect 14242 -2916 14252 -2906
rect 14492 -2906 14572 -2896
rect 14492 -2916 14502 -2906
rect 14242 -2966 14502 -2916
rect 14562 -2966 14572 -2906
rect 14172 -2976 14572 -2966
rect 14630 -2556 15030 -2546
rect 14630 -2616 14640 -2556
rect 14700 -2606 14960 -2556
rect 14700 -2616 14710 -2606
rect 14630 -2626 14710 -2616
rect 14950 -2616 14960 -2606
rect 15020 -2616 15030 -2556
rect 14950 -2626 15030 -2616
rect 14630 -2896 14690 -2626
rect 14960 -2636 15030 -2626
rect 14770 -2686 14800 -2666
rect 14750 -2726 14800 -2686
rect 14860 -2686 14890 -2666
rect 14860 -2726 14910 -2686
rect 14750 -2796 14910 -2726
rect 14750 -2836 14800 -2796
rect 14770 -2856 14800 -2836
rect 14860 -2836 14910 -2796
rect 14860 -2856 14890 -2836
rect 14970 -2896 15030 -2636
rect 14630 -2906 14710 -2896
rect 14630 -2966 14640 -2906
rect 14700 -2916 14710 -2906
rect 14950 -2906 15030 -2896
rect 14950 -2916 14960 -2906
rect 14700 -2966 14960 -2916
rect 15020 -2966 15030 -2906
rect 14630 -2976 15030 -2966
rect 15086 -2556 15486 -2546
rect 15086 -2616 15096 -2556
rect 15156 -2606 15416 -2556
rect 15156 -2616 15166 -2606
rect 15086 -2626 15166 -2616
rect 15406 -2616 15416 -2606
rect 15476 -2616 15486 -2556
rect 15406 -2626 15486 -2616
rect 15086 -2896 15146 -2626
rect 15416 -2636 15486 -2626
rect 15226 -2686 15256 -2666
rect 15206 -2726 15256 -2686
rect 15316 -2686 15346 -2666
rect 15316 -2726 15366 -2686
rect 15206 -2796 15366 -2726
rect 15206 -2836 15256 -2796
rect 15226 -2856 15256 -2836
rect 15316 -2836 15366 -2796
rect 15316 -2856 15346 -2836
rect 15426 -2896 15486 -2636
rect 15086 -2906 15166 -2896
rect 15086 -2966 15096 -2906
rect 15156 -2916 15166 -2906
rect 15406 -2906 15486 -2896
rect 15406 -2916 15416 -2906
rect 15156 -2966 15416 -2916
rect 15476 -2966 15486 -2906
rect 15086 -2976 15486 -2966
rect 0 -3552 400 -3542
rect 0 -3612 10 -3552
rect 70 -3602 330 -3552
rect 70 -3612 80 -3602
rect 0 -3622 80 -3612
rect 320 -3612 330 -3602
rect 390 -3612 400 -3552
rect 320 -3622 400 -3612
rect 0 -3892 60 -3622
rect 330 -3632 400 -3622
rect 140 -3682 170 -3662
rect 120 -3722 170 -3682
rect 230 -3682 260 -3662
rect 230 -3722 280 -3682
rect 120 -3792 280 -3722
rect 120 -3832 170 -3792
rect 140 -3852 170 -3832
rect 230 -3832 280 -3792
rect 230 -3852 260 -3832
rect 340 -3892 400 -3632
rect 0 -3902 80 -3892
rect 0 -3962 10 -3902
rect 70 -3912 80 -3902
rect 320 -3902 400 -3892
rect 320 -3912 330 -3902
rect 70 -3962 330 -3912
rect 390 -3962 400 -3902
rect 0 -3972 400 -3962
rect 456 -3552 856 -3542
rect 456 -3612 466 -3552
rect 526 -3602 786 -3552
rect 526 -3612 536 -3602
rect 456 -3622 536 -3612
rect 776 -3612 786 -3602
rect 846 -3612 856 -3552
rect 776 -3622 856 -3612
rect 456 -3892 516 -3622
rect 786 -3632 856 -3622
rect 596 -3682 626 -3662
rect 576 -3722 626 -3682
rect 686 -3682 716 -3662
rect 686 -3722 736 -3682
rect 576 -3792 736 -3722
rect 576 -3832 626 -3792
rect 596 -3852 626 -3832
rect 686 -3832 736 -3792
rect 686 -3852 716 -3832
rect 796 -3892 856 -3632
rect 456 -3902 536 -3892
rect 456 -3962 466 -3902
rect 526 -3912 536 -3902
rect 776 -3902 856 -3892
rect 776 -3912 786 -3902
rect 526 -3962 786 -3912
rect 846 -3962 856 -3902
rect 456 -3972 856 -3962
rect 912 -3552 1312 -3542
rect 912 -3612 922 -3552
rect 982 -3602 1242 -3552
rect 982 -3612 992 -3602
rect 912 -3622 992 -3612
rect 1232 -3612 1242 -3602
rect 1302 -3612 1312 -3552
rect 1232 -3622 1312 -3612
rect 912 -3892 972 -3622
rect 1242 -3632 1312 -3622
rect 1052 -3682 1082 -3662
rect 1032 -3722 1082 -3682
rect 1142 -3682 1172 -3662
rect 1142 -3722 1192 -3682
rect 1032 -3792 1192 -3722
rect 1032 -3832 1082 -3792
rect 1052 -3852 1082 -3832
rect 1142 -3832 1192 -3792
rect 1142 -3852 1172 -3832
rect 1252 -3892 1312 -3632
rect 912 -3902 992 -3892
rect 912 -3962 922 -3902
rect 982 -3912 992 -3902
rect 1232 -3902 1312 -3892
rect 1232 -3912 1242 -3902
rect 982 -3962 1242 -3912
rect 1302 -3962 1312 -3902
rect 912 -3972 1312 -3962
rect 1370 -3552 1770 -3542
rect 1370 -3612 1380 -3552
rect 1440 -3602 1700 -3552
rect 1440 -3612 1450 -3602
rect 1370 -3622 1450 -3612
rect 1690 -3612 1700 -3602
rect 1760 -3612 1770 -3552
rect 1690 -3622 1770 -3612
rect 1370 -3892 1430 -3622
rect 1700 -3632 1770 -3622
rect 1510 -3682 1540 -3662
rect 1490 -3722 1540 -3682
rect 1600 -3682 1630 -3662
rect 1600 -3722 1650 -3682
rect 1490 -3792 1650 -3722
rect 1490 -3832 1540 -3792
rect 1510 -3852 1540 -3832
rect 1600 -3832 1650 -3792
rect 1600 -3852 1630 -3832
rect 1710 -3892 1770 -3632
rect 1370 -3902 1450 -3892
rect 1370 -3962 1380 -3902
rect 1440 -3912 1450 -3902
rect 1690 -3902 1770 -3892
rect 1690 -3912 1700 -3902
rect 1440 -3962 1700 -3912
rect 1760 -3962 1770 -3902
rect 1370 -3972 1770 -3962
rect 1826 -3552 2226 -3542
rect 1826 -3612 1836 -3552
rect 1896 -3602 2156 -3552
rect 1896 -3612 1906 -3602
rect 1826 -3622 1906 -3612
rect 2146 -3612 2156 -3602
rect 2216 -3612 2226 -3552
rect 2146 -3622 2226 -3612
rect 1826 -3892 1886 -3622
rect 2156 -3632 2226 -3622
rect 1966 -3682 1996 -3662
rect 1946 -3722 1996 -3682
rect 2056 -3682 2086 -3662
rect 2056 -3722 2106 -3682
rect 1946 -3792 2106 -3722
rect 1946 -3832 1996 -3792
rect 1966 -3852 1996 -3832
rect 2056 -3832 2106 -3792
rect 2056 -3852 2086 -3832
rect 2166 -3892 2226 -3632
rect 1826 -3902 1906 -3892
rect 1826 -3962 1836 -3902
rect 1896 -3912 1906 -3902
rect 2146 -3902 2226 -3892
rect 2146 -3912 2156 -3902
rect 1896 -3962 2156 -3912
rect 2216 -3962 2226 -3902
rect 1826 -3972 2226 -3962
rect 2282 -3552 2682 -3542
rect 2282 -3612 2292 -3552
rect 2352 -3602 2612 -3552
rect 2352 -3612 2362 -3602
rect 2282 -3622 2362 -3612
rect 2602 -3612 2612 -3602
rect 2672 -3612 2682 -3552
rect 2602 -3622 2682 -3612
rect 2282 -3892 2342 -3622
rect 2612 -3632 2682 -3622
rect 2422 -3682 2452 -3662
rect 2402 -3722 2452 -3682
rect 2512 -3682 2542 -3662
rect 2512 -3722 2562 -3682
rect 2402 -3792 2562 -3722
rect 2402 -3832 2452 -3792
rect 2422 -3852 2452 -3832
rect 2512 -3832 2562 -3792
rect 2512 -3852 2542 -3832
rect 2622 -3892 2682 -3632
rect 2282 -3902 2362 -3892
rect 2282 -3962 2292 -3902
rect 2352 -3912 2362 -3902
rect 2602 -3902 2682 -3892
rect 2602 -3912 2612 -3902
rect 2352 -3962 2612 -3912
rect 2672 -3962 2682 -3902
rect 2282 -3972 2682 -3962
rect 2740 -3552 3140 -3542
rect 2740 -3612 2750 -3552
rect 2810 -3602 3070 -3552
rect 2810 -3612 2820 -3602
rect 2740 -3622 2820 -3612
rect 3060 -3612 3070 -3602
rect 3130 -3612 3140 -3552
rect 3060 -3622 3140 -3612
rect 2740 -3892 2800 -3622
rect 3070 -3632 3140 -3622
rect 2880 -3682 2910 -3662
rect 2860 -3722 2910 -3682
rect 2970 -3682 3000 -3662
rect 2970 -3722 3020 -3682
rect 2860 -3792 3020 -3722
rect 2860 -3832 2910 -3792
rect 2880 -3852 2910 -3832
rect 2970 -3832 3020 -3792
rect 2970 -3852 3000 -3832
rect 3080 -3892 3140 -3632
rect 2740 -3902 2820 -3892
rect 2740 -3962 2750 -3902
rect 2810 -3912 2820 -3902
rect 3060 -3902 3140 -3892
rect 3060 -3912 3070 -3902
rect 2810 -3962 3070 -3912
rect 3130 -3962 3140 -3902
rect 2740 -3972 3140 -3962
rect 3196 -3552 3596 -3542
rect 3196 -3612 3206 -3552
rect 3266 -3602 3526 -3552
rect 3266 -3612 3276 -3602
rect 3196 -3622 3276 -3612
rect 3516 -3612 3526 -3602
rect 3586 -3612 3596 -3552
rect 3516 -3622 3596 -3612
rect 3196 -3892 3256 -3622
rect 3526 -3632 3596 -3622
rect 3336 -3682 3366 -3662
rect 3316 -3722 3366 -3682
rect 3426 -3682 3456 -3662
rect 3426 -3722 3476 -3682
rect 3316 -3792 3476 -3722
rect 3316 -3832 3366 -3792
rect 3336 -3852 3366 -3832
rect 3426 -3832 3476 -3792
rect 3426 -3852 3456 -3832
rect 3536 -3892 3596 -3632
rect 3196 -3902 3276 -3892
rect 3196 -3962 3206 -3902
rect 3266 -3912 3276 -3902
rect 3516 -3902 3596 -3892
rect 3516 -3912 3526 -3902
rect 3266 -3962 3526 -3912
rect 3586 -3962 3596 -3902
rect 3196 -3972 3596 -3962
rect 3652 -3552 4052 -3542
rect 3652 -3612 3662 -3552
rect 3722 -3602 3982 -3552
rect 3722 -3612 3732 -3602
rect 3652 -3622 3732 -3612
rect 3972 -3612 3982 -3602
rect 4042 -3612 4052 -3552
rect 3972 -3622 4052 -3612
rect 3652 -3892 3712 -3622
rect 3982 -3632 4052 -3622
rect 3792 -3682 3822 -3662
rect 3772 -3722 3822 -3682
rect 3882 -3682 3912 -3662
rect 3882 -3722 3932 -3682
rect 3772 -3792 3932 -3722
rect 3772 -3832 3822 -3792
rect 3792 -3852 3822 -3832
rect 3882 -3832 3932 -3792
rect 3882 -3852 3912 -3832
rect 3992 -3892 4052 -3632
rect 3652 -3902 3732 -3892
rect 3652 -3962 3662 -3902
rect 3722 -3912 3732 -3902
rect 3972 -3902 4052 -3892
rect 3972 -3912 3982 -3902
rect 3722 -3962 3982 -3912
rect 4042 -3962 4052 -3902
rect 3652 -3972 4052 -3962
rect 4110 -3552 4510 -3542
rect 4110 -3612 4120 -3552
rect 4180 -3602 4440 -3552
rect 4180 -3612 4190 -3602
rect 4110 -3622 4190 -3612
rect 4430 -3612 4440 -3602
rect 4500 -3612 4510 -3552
rect 4430 -3622 4510 -3612
rect 4110 -3892 4170 -3622
rect 4440 -3632 4510 -3622
rect 4250 -3682 4280 -3662
rect 4230 -3722 4280 -3682
rect 4340 -3682 4370 -3662
rect 4340 -3722 4390 -3682
rect 4230 -3792 4390 -3722
rect 4230 -3832 4280 -3792
rect 4250 -3852 4280 -3832
rect 4340 -3832 4390 -3792
rect 4340 -3852 4370 -3832
rect 4450 -3892 4510 -3632
rect 4110 -3902 4190 -3892
rect 4110 -3962 4120 -3902
rect 4180 -3912 4190 -3902
rect 4430 -3902 4510 -3892
rect 4430 -3912 4440 -3902
rect 4180 -3962 4440 -3912
rect 4500 -3962 4510 -3902
rect 4110 -3972 4510 -3962
rect 4566 -3552 4966 -3542
rect 4566 -3612 4576 -3552
rect 4636 -3602 4896 -3552
rect 4636 -3612 4646 -3602
rect 4566 -3622 4646 -3612
rect 4886 -3612 4896 -3602
rect 4956 -3612 4966 -3552
rect 4886 -3622 4966 -3612
rect 4566 -3892 4626 -3622
rect 4896 -3632 4966 -3622
rect 4706 -3682 4736 -3662
rect 4686 -3722 4736 -3682
rect 4796 -3682 4826 -3662
rect 4796 -3722 4846 -3682
rect 4686 -3792 4846 -3722
rect 4686 -3832 4736 -3792
rect 4706 -3852 4736 -3832
rect 4796 -3832 4846 -3792
rect 4796 -3852 4826 -3832
rect 4906 -3892 4966 -3632
rect 4566 -3902 4646 -3892
rect 4566 -3962 4576 -3902
rect 4636 -3912 4646 -3902
rect 4886 -3902 4966 -3892
rect 4886 -3912 4896 -3902
rect 4636 -3962 4896 -3912
rect 4956 -3962 4966 -3902
rect 4566 -3972 4966 -3962
rect 5022 -3552 5422 -3542
rect 5022 -3612 5032 -3552
rect 5092 -3602 5352 -3552
rect 5092 -3612 5102 -3602
rect 5022 -3622 5102 -3612
rect 5342 -3612 5352 -3602
rect 5412 -3612 5422 -3552
rect 5342 -3622 5422 -3612
rect 5022 -3892 5082 -3622
rect 5352 -3632 5422 -3622
rect 5162 -3682 5192 -3662
rect 5142 -3722 5192 -3682
rect 5252 -3682 5282 -3662
rect 5252 -3722 5302 -3682
rect 5142 -3792 5302 -3722
rect 5142 -3832 5192 -3792
rect 5162 -3852 5192 -3832
rect 5252 -3832 5302 -3792
rect 5252 -3852 5282 -3832
rect 5362 -3892 5422 -3632
rect 5022 -3902 5102 -3892
rect 5022 -3962 5032 -3902
rect 5092 -3912 5102 -3902
rect 5342 -3902 5422 -3892
rect 5342 -3912 5352 -3902
rect 5092 -3962 5352 -3912
rect 5412 -3962 5422 -3902
rect 5022 -3972 5422 -3962
rect 5480 -3552 5880 -3542
rect 5480 -3612 5490 -3552
rect 5550 -3602 5810 -3552
rect 5550 -3612 5560 -3602
rect 5480 -3622 5560 -3612
rect 5800 -3612 5810 -3602
rect 5870 -3612 5880 -3552
rect 5800 -3622 5880 -3612
rect 5480 -3892 5540 -3622
rect 5810 -3632 5880 -3622
rect 5620 -3682 5650 -3662
rect 5600 -3722 5650 -3682
rect 5710 -3682 5740 -3662
rect 5710 -3722 5760 -3682
rect 5600 -3792 5760 -3722
rect 5600 -3832 5650 -3792
rect 5620 -3852 5650 -3832
rect 5710 -3832 5760 -3792
rect 5710 -3852 5740 -3832
rect 5820 -3892 5880 -3632
rect 5480 -3902 5560 -3892
rect 5480 -3962 5490 -3902
rect 5550 -3912 5560 -3902
rect 5800 -3902 5880 -3892
rect 5800 -3912 5810 -3902
rect 5550 -3962 5810 -3912
rect 5870 -3962 5880 -3902
rect 5480 -3972 5880 -3962
rect 5936 -3552 6336 -3542
rect 5936 -3612 5946 -3552
rect 6006 -3602 6266 -3552
rect 6006 -3612 6016 -3602
rect 5936 -3622 6016 -3612
rect 6256 -3612 6266 -3602
rect 6326 -3612 6336 -3552
rect 6256 -3622 6336 -3612
rect 5936 -3892 5996 -3622
rect 6266 -3632 6336 -3622
rect 6076 -3682 6106 -3662
rect 6056 -3722 6106 -3682
rect 6166 -3682 6196 -3662
rect 6166 -3722 6216 -3682
rect 6056 -3792 6216 -3722
rect 6056 -3832 6106 -3792
rect 6076 -3852 6106 -3832
rect 6166 -3832 6216 -3792
rect 6166 -3852 6196 -3832
rect 6276 -3892 6336 -3632
rect 5936 -3902 6016 -3892
rect 5936 -3962 5946 -3902
rect 6006 -3912 6016 -3902
rect 6256 -3902 6336 -3892
rect 6256 -3912 6266 -3902
rect 6006 -3962 6266 -3912
rect 6326 -3962 6336 -3902
rect 5936 -3972 6336 -3962
rect 6392 -3552 6792 -3542
rect 6392 -3612 6402 -3552
rect 6462 -3602 6722 -3552
rect 6462 -3612 6472 -3602
rect 6392 -3622 6472 -3612
rect 6712 -3612 6722 -3602
rect 6782 -3612 6792 -3552
rect 6712 -3622 6792 -3612
rect 6392 -3892 6452 -3622
rect 6722 -3632 6792 -3622
rect 6532 -3682 6562 -3662
rect 6512 -3722 6562 -3682
rect 6622 -3682 6652 -3662
rect 6622 -3722 6672 -3682
rect 6512 -3792 6672 -3722
rect 6512 -3832 6562 -3792
rect 6532 -3852 6562 -3832
rect 6622 -3832 6672 -3792
rect 6622 -3852 6652 -3832
rect 6732 -3892 6792 -3632
rect 6392 -3902 6472 -3892
rect 6392 -3962 6402 -3902
rect 6462 -3912 6472 -3902
rect 6712 -3902 6792 -3892
rect 6712 -3912 6722 -3902
rect 6462 -3962 6722 -3912
rect 6782 -3962 6792 -3902
rect 6392 -3972 6792 -3962
rect 6850 -3552 7250 -3542
rect 6850 -3612 6860 -3552
rect 6920 -3602 7180 -3552
rect 6920 -3612 6930 -3602
rect 6850 -3622 6930 -3612
rect 7170 -3612 7180 -3602
rect 7240 -3612 7250 -3552
rect 7170 -3622 7250 -3612
rect 6850 -3892 6910 -3622
rect 7180 -3632 7250 -3622
rect 6990 -3682 7020 -3662
rect 6970 -3722 7020 -3682
rect 7080 -3682 7110 -3662
rect 7080 -3722 7130 -3682
rect 6970 -3792 7130 -3722
rect 6970 -3832 7020 -3792
rect 6990 -3852 7020 -3832
rect 7080 -3832 7130 -3792
rect 7080 -3852 7110 -3832
rect 7190 -3892 7250 -3632
rect 6850 -3902 6930 -3892
rect 6850 -3962 6860 -3902
rect 6920 -3912 6930 -3902
rect 7170 -3902 7250 -3892
rect 7170 -3912 7180 -3902
rect 6920 -3962 7180 -3912
rect 7240 -3962 7250 -3902
rect 6850 -3972 7250 -3962
rect 7306 -3552 7706 -3542
rect 7306 -3612 7316 -3552
rect 7376 -3602 7636 -3552
rect 7376 -3612 7386 -3602
rect 7306 -3622 7386 -3612
rect 7626 -3612 7636 -3602
rect 7696 -3612 7706 -3552
rect 7626 -3622 7706 -3612
rect 7306 -3892 7366 -3622
rect 7636 -3632 7706 -3622
rect 7446 -3682 7476 -3662
rect 7426 -3722 7476 -3682
rect 7536 -3682 7566 -3662
rect 7536 -3722 7586 -3682
rect 7426 -3792 7586 -3722
rect 7426 -3832 7476 -3792
rect 7446 -3852 7476 -3832
rect 7536 -3832 7586 -3792
rect 7536 -3852 7566 -3832
rect 7646 -3892 7706 -3632
rect 7306 -3902 7386 -3892
rect 7306 -3962 7316 -3902
rect 7376 -3912 7386 -3902
rect 7626 -3902 7706 -3892
rect 7626 -3912 7636 -3902
rect 7376 -3962 7636 -3912
rect 7696 -3962 7706 -3902
rect 7306 -3972 7706 -3962
rect 7762 -3552 8162 -3542
rect 7762 -3612 7772 -3552
rect 7832 -3602 8092 -3552
rect 7832 -3612 7842 -3602
rect 7762 -3622 7842 -3612
rect 8082 -3612 8092 -3602
rect 8152 -3612 8162 -3552
rect 8082 -3622 8162 -3612
rect 7762 -3892 7822 -3622
rect 8092 -3632 8162 -3622
rect 7902 -3682 7932 -3662
rect 7882 -3722 7932 -3682
rect 7992 -3682 8022 -3662
rect 7992 -3722 8042 -3682
rect 7882 -3792 8042 -3722
rect 7882 -3832 7932 -3792
rect 7902 -3852 7932 -3832
rect 7992 -3832 8042 -3792
rect 7992 -3852 8022 -3832
rect 8102 -3892 8162 -3632
rect 7762 -3902 7842 -3892
rect 7762 -3962 7772 -3902
rect 7832 -3912 7842 -3902
rect 8082 -3902 8162 -3892
rect 8082 -3912 8092 -3902
rect 7832 -3962 8092 -3912
rect 8152 -3962 8162 -3902
rect 7762 -3972 8162 -3962
rect 8236 -3552 8636 -3542
rect 8236 -3612 8246 -3552
rect 8306 -3602 8566 -3552
rect 8306 -3612 8316 -3602
rect 8236 -3622 8316 -3612
rect 8556 -3612 8566 -3602
rect 8626 -3612 8636 -3552
rect 8556 -3622 8636 -3612
rect 8236 -3892 8296 -3622
rect 8566 -3632 8636 -3622
rect 8376 -3682 8406 -3662
rect 8356 -3722 8406 -3682
rect 8466 -3682 8496 -3662
rect 8466 -3722 8516 -3682
rect 8356 -3792 8516 -3722
rect 8356 -3832 8406 -3792
rect 8376 -3852 8406 -3832
rect 8466 -3832 8516 -3792
rect 8466 -3852 8496 -3832
rect 8576 -3892 8636 -3632
rect 8236 -3902 8316 -3892
rect 8236 -3962 8246 -3902
rect 8306 -3912 8316 -3902
rect 8556 -3902 8636 -3892
rect 8556 -3912 8566 -3902
rect 8306 -3962 8566 -3912
rect 8626 -3962 8636 -3902
rect 8236 -3972 8636 -3962
rect 8692 -3552 9092 -3542
rect 8692 -3612 8702 -3552
rect 8762 -3602 9022 -3552
rect 8762 -3612 8772 -3602
rect 8692 -3622 8772 -3612
rect 9012 -3612 9022 -3602
rect 9082 -3612 9092 -3552
rect 9012 -3622 9092 -3612
rect 8692 -3892 8752 -3622
rect 9022 -3632 9092 -3622
rect 8832 -3682 8862 -3662
rect 8812 -3722 8862 -3682
rect 8922 -3682 8952 -3662
rect 8922 -3722 8972 -3682
rect 8812 -3792 8972 -3722
rect 8812 -3832 8862 -3792
rect 8832 -3852 8862 -3832
rect 8922 -3832 8972 -3792
rect 8922 -3852 8952 -3832
rect 9032 -3892 9092 -3632
rect 8692 -3902 8772 -3892
rect 8692 -3962 8702 -3902
rect 8762 -3912 8772 -3902
rect 9012 -3902 9092 -3892
rect 9012 -3912 9022 -3902
rect 8762 -3962 9022 -3912
rect 9082 -3962 9092 -3902
rect 8692 -3972 9092 -3962
rect 9150 -3552 9550 -3542
rect 9150 -3612 9160 -3552
rect 9220 -3602 9480 -3552
rect 9220 -3612 9230 -3602
rect 9150 -3622 9230 -3612
rect 9470 -3612 9480 -3602
rect 9540 -3612 9550 -3552
rect 9470 -3622 9550 -3612
rect 9150 -3892 9210 -3622
rect 9480 -3632 9550 -3622
rect 9290 -3682 9320 -3662
rect 9270 -3722 9320 -3682
rect 9380 -3682 9410 -3662
rect 9380 -3722 9430 -3682
rect 9270 -3792 9430 -3722
rect 9270 -3832 9320 -3792
rect 9290 -3852 9320 -3832
rect 9380 -3832 9430 -3792
rect 9380 -3852 9410 -3832
rect 9490 -3892 9550 -3632
rect 9150 -3902 9230 -3892
rect 9150 -3962 9160 -3902
rect 9220 -3912 9230 -3902
rect 9470 -3902 9550 -3892
rect 9470 -3912 9480 -3902
rect 9220 -3962 9480 -3912
rect 9540 -3962 9550 -3902
rect 9150 -3972 9550 -3962
rect 9606 -3552 10006 -3542
rect 9606 -3612 9616 -3552
rect 9676 -3602 9936 -3552
rect 9676 -3612 9686 -3602
rect 9606 -3622 9686 -3612
rect 9926 -3612 9936 -3602
rect 9996 -3612 10006 -3552
rect 9926 -3622 10006 -3612
rect 9606 -3892 9666 -3622
rect 9936 -3632 10006 -3622
rect 9746 -3682 9776 -3662
rect 9726 -3722 9776 -3682
rect 9836 -3682 9866 -3662
rect 9836 -3722 9886 -3682
rect 9726 -3792 9886 -3722
rect 9726 -3832 9776 -3792
rect 9746 -3852 9776 -3832
rect 9836 -3832 9886 -3792
rect 9836 -3852 9866 -3832
rect 9946 -3892 10006 -3632
rect 9606 -3902 9686 -3892
rect 9606 -3962 9616 -3902
rect 9676 -3912 9686 -3902
rect 9926 -3902 10006 -3892
rect 9926 -3912 9936 -3902
rect 9676 -3962 9936 -3912
rect 9996 -3962 10006 -3902
rect 9606 -3972 10006 -3962
rect 10062 -3552 10462 -3542
rect 10062 -3612 10072 -3552
rect 10132 -3602 10392 -3552
rect 10132 -3612 10142 -3602
rect 10062 -3622 10142 -3612
rect 10382 -3612 10392 -3602
rect 10452 -3612 10462 -3552
rect 10382 -3622 10462 -3612
rect 10062 -3892 10122 -3622
rect 10392 -3632 10462 -3622
rect 10202 -3682 10232 -3662
rect 10182 -3722 10232 -3682
rect 10292 -3682 10322 -3662
rect 10292 -3722 10342 -3682
rect 10182 -3792 10342 -3722
rect 10182 -3832 10232 -3792
rect 10202 -3852 10232 -3832
rect 10292 -3832 10342 -3792
rect 10292 -3852 10322 -3832
rect 10402 -3892 10462 -3632
rect 10062 -3902 10142 -3892
rect 10062 -3962 10072 -3902
rect 10132 -3912 10142 -3902
rect 10382 -3902 10462 -3892
rect 10382 -3912 10392 -3902
rect 10132 -3962 10392 -3912
rect 10452 -3962 10462 -3902
rect 10062 -3972 10462 -3962
rect 10520 -3552 10920 -3542
rect 10520 -3612 10530 -3552
rect 10590 -3602 10850 -3552
rect 10590 -3612 10600 -3602
rect 10520 -3622 10600 -3612
rect 10840 -3612 10850 -3602
rect 10910 -3612 10920 -3552
rect 10840 -3622 10920 -3612
rect 10520 -3892 10580 -3622
rect 10850 -3632 10920 -3622
rect 10660 -3682 10690 -3662
rect 10640 -3722 10690 -3682
rect 10750 -3682 10780 -3662
rect 10750 -3722 10800 -3682
rect 10640 -3792 10800 -3722
rect 10640 -3832 10690 -3792
rect 10660 -3852 10690 -3832
rect 10750 -3832 10800 -3792
rect 10750 -3852 10780 -3832
rect 10860 -3892 10920 -3632
rect 10520 -3902 10600 -3892
rect 10520 -3962 10530 -3902
rect 10590 -3912 10600 -3902
rect 10840 -3902 10920 -3892
rect 10840 -3912 10850 -3902
rect 10590 -3962 10850 -3912
rect 10910 -3962 10920 -3902
rect 10520 -3972 10920 -3962
rect 10976 -3552 11376 -3542
rect 10976 -3612 10986 -3552
rect 11046 -3602 11306 -3552
rect 11046 -3612 11056 -3602
rect 10976 -3622 11056 -3612
rect 11296 -3612 11306 -3602
rect 11366 -3612 11376 -3552
rect 11296 -3622 11376 -3612
rect 10976 -3892 11036 -3622
rect 11306 -3632 11376 -3622
rect 11116 -3682 11146 -3662
rect 11096 -3722 11146 -3682
rect 11206 -3682 11236 -3662
rect 11206 -3722 11256 -3682
rect 11096 -3792 11256 -3722
rect 11096 -3832 11146 -3792
rect 11116 -3852 11146 -3832
rect 11206 -3832 11256 -3792
rect 11206 -3852 11236 -3832
rect 11316 -3892 11376 -3632
rect 10976 -3902 11056 -3892
rect 10976 -3962 10986 -3902
rect 11046 -3912 11056 -3902
rect 11296 -3902 11376 -3892
rect 11296 -3912 11306 -3902
rect 11046 -3962 11306 -3912
rect 11366 -3962 11376 -3902
rect 10976 -3972 11376 -3962
rect 11432 -3552 11832 -3542
rect 11432 -3612 11442 -3552
rect 11502 -3602 11762 -3552
rect 11502 -3612 11512 -3602
rect 11432 -3622 11512 -3612
rect 11752 -3612 11762 -3602
rect 11822 -3612 11832 -3552
rect 11752 -3622 11832 -3612
rect 11432 -3892 11492 -3622
rect 11762 -3632 11832 -3622
rect 11572 -3682 11602 -3662
rect 11552 -3722 11602 -3682
rect 11662 -3682 11692 -3662
rect 11662 -3722 11712 -3682
rect 11552 -3792 11712 -3722
rect 11552 -3832 11602 -3792
rect 11572 -3852 11602 -3832
rect 11662 -3832 11712 -3792
rect 11662 -3852 11692 -3832
rect 11772 -3892 11832 -3632
rect 11432 -3902 11512 -3892
rect 11432 -3962 11442 -3902
rect 11502 -3912 11512 -3902
rect 11752 -3902 11832 -3892
rect 11752 -3912 11762 -3902
rect 11502 -3962 11762 -3912
rect 11822 -3962 11832 -3902
rect 11432 -3972 11832 -3962
rect 11890 -3552 12290 -3542
rect 11890 -3612 11900 -3552
rect 11960 -3602 12220 -3552
rect 11960 -3612 11970 -3602
rect 11890 -3622 11970 -3612
rect 12210 -3612 12220 -3602
rect 12280 -3612 12290 -3552
rect 12210 -3622 12290 -3612
rect 11890 -3892 11950 -3622
rect 12220 -3632 12290 -3622
rect 12030 -3682 12060 -3662
rect 12010 -3722 12060 -3682
rect 12120 -3682 12150 -3662
rect 12120 -3722 12170 -3682
rect 12010 -3792 12170 -3722
rect 12010 -3832 12060 -3792
rect 12030 -3852 12060 -3832
rect 12120 -3832 12170 -3792
rect 12120 -3852 12150 -3832
rect 12230 -3892 12290 -3632
rect 11890 -3902 11970 -3892
rect 11890 -3962 11900 -3902
rect 11960 -3912 11970 -3902
rect 12210 -3902 12290 -3892
rect 12210 -3912 12220 -3902
rect 11960 -3962 12220 -3912
rect 12280 -3962 12290 -3902
rect 11890 -3972 12290 -3962
rect 12346 -3552 12746 -3542
rect 12346 -3612 12356 -3552
rect 12416 -3602 12676 -3552
rect 12416 -3612 12426 -3602
rect 12346 -3622 12426 -3612
rect 12666 -3612 12676 -3602
rect 12736 -3612 12746 -3552
rect 12666 -3622 12746 -3612
rect 12346 -3892 12406 -3622
rect 12676 -3632 12746 -3622
rect 12486 -3682 12516 -3662
rect 12466 -3722 12516 -3682
rect 12576 -3682 12606 -3662
rect 12576 -3722 12626 -3682
rect 12466 -3792 12626 -3722
rect 12466 -3832 12516 -3792
rect 12486 -3852 12516 -3832
rect 12576 -3832 12626 -3792
rect 12576 -3852 12606 -3832
rect 12686 -3892 12746 -3632
rect 12346 -3902 12426 -3892
rect 12346 -3962 12356 -3902
rect 12416 -3912 12426 -3902
rect 12666 -3902 12746 -3892
rect 12666 -3912 12676 -3902
rect 12416 -3962 12676 -3912
rect 12736 -3962 12746 -3902
rect 12346 -3972 12746 -3962
rect 12802 -3552 13202 -3542
rect 12802 -3612 12812 -3552
rect 12872 -3602 13132 -3552
rect 12872 -3612 12882 -3602
rect 12802 -3622 12882 -3612
rect 13122 -3612 13132 -3602
rect 13192 -3612 13202 -3552
rect 13122 -3622 13202 -3612
rect 12802 -3892 12862 -3622
rect 13132 -3632 13202 -3622
rect 12942 -3682 12972 -3662
rect 12922 -3722 12972 -3682
rect 13032 -3682 13062 -3662
rect 13032 -3722 13082 -3682
rect 12922 -3792 13082 -3722
rect 12922 -3832 12972 -3792
rect 12942 -3852 12972 -3832
rect 13032 -3832 13082 -3792
rect 13032 -3852 13062 -3832
rect 13142 -3892 13202 -3632
rect 12802 -3902 12882 -3892
rect 12802 -3962 12812 -3902
rect 12872 -3912 12882 -3902
rect 13122 -3902 13202 -3892
rect 13122 -3912 13132 -3902
rect 12872 -3962 13132 -3912
rect 13192 -3962 13202 -3902
rect 12802 -3972 13202 -3962
rect 13260 -3552 13660 -3542
rect 13260 -3612 13270 -3552
rect 13330 -3602 13590 -3552
rect 13330 -3612 13340 -3602
rect 13260 -3622 13340 -3612
rect 13580 -3612 13590 -3602
rect 13650 -3612 13660 -3552
rect 13580 -3622 13660 -3612
rect 13260 -3892 13320 -3622
rect 13590 -3632 13660 -3622
rect 13400 -3682 13430 -3662
rect 13380 -3722 13430 -3682
rect 13490 -3682 13520 -3662
rect 13490 -3722 13540 -3682
rect 13380 -3792 13540 -3722
rect 13380 -3832 13430 -3792
rect 13400 -3852 13430 -3832
rect 13490 -3832 13540 -3792
rect 13490 -3852 13520 -3832
rect 13600 -3892 13660 -3632
rect 13260 -3902 13340 -3892
rect 13260 -3962 13270 -3902
rect 13330 -3912 13340 -3902
rect 13580 -3902 13660 -3892
rect 13580 -3912 13590 -3902
rect 13330 -3962 13590 -3912
rect 13650 -3962 13660 -3902
rect 13260 -3972 13660 -3962
rect 13716 -3552 14116 -3542
rect 13716 -3612 13726 -3552
rect 13786 -3602 14046 -3552
rect 13786 -3612 13796 -3602
rect 13716 -3622 13796 -3612
rect 14036 -3612 14046 -3602
rect 14106 -3612 14116 -3552
rect 14036 -3622 14116 -3612
rect 13716 -3892 13776 -3622
rect 14046 -3632 14116 -3622
rect 13856 -3682 13886 -3662
rect 13836 -3722 13886 -3682
rect 13946 -3682 13976 -3662
rect 13946 -3722 13996 -3682
rect 13836 -3792 13996 -3722
rect 13836 -3832 13886 -3792
rect 13856 -3852 13886 -3832
rect 13946 -3832 13996 -3792
rect 13946 -3852 13976 -3832
rect 14056 -3892 14116 -3632
rect 13716 -3902 13796 -3892
rect 13716 -3962 13726 -3902
rect 13786 -3912 13796 -3902
rect 14036 -3902 14116 -3892
rect 14036 -3912 14046 -3902
rect 13786 -3962 14046 -3912
rect 14106 -3962 14116 -3902
rect 13716 -3972 14116 -3962
rect 14172 -3552 14572 -3542
rect 14172 -3612 14182 -3552
rect 14242 -3602 14502 -3552
rect 14242 -3612 14252 -3602
rect 14172 -3622 14252 -3612
rect 14492 -3612 14502 -3602
rect 14562 -3612 14572 -3552
rect 14492 -3622 14572 -3612
rect 14172 -3892 14232 -3622
rect 14502 -3632 14572 -3622
rect 14312 -3682 14342 -3662
rect 14292 -3722 14342 -3682
rect 14402 -3682 14432 -3662
rect 14402 -3722 14452 -3682
rect 14292 -3792 14452 -3722
rect 14292 -3832 14342 -3792
rect 14312 -3852 14342 -3832
rect 14402 -3832 14452 -3792
rect 14402 -3852 14432 -3832
rect 14512 -3892 14572 -3632
rect 14172 -3902 14252 -3892
rect 14172 -3962 14182 -3902
rect 14242 -3912 14252 -3902
rect 14492 -3902 14572 -3892
rect 14492 -3912 14502 -3902
rect 14242 -3962 14502 -3912
rect 14562 -3962 14572 -3902
rect 14172 -3972 14572 -3962
rect 14630 -3552 15030 -3542
rect 14630 -3612 14640 -3552
rect 14700 -3602 14960 -3552
rect 14700 -3612 14710 -3602
rect 14630 -3622 14710 -3612
rect 14950 -3612 14960 -3602
rect 15020 -3612 15030 -3552
rect 14950 -3622 15030 -3612
rect 14630 -3892 14690 -3622
rect 14960 -3632 15030 -3622
rect 14770 -3682 14800 -3662
rect 14750 -3722 14800 -3682
rect 14860 -3682 14890 -3662
rect 14860 -3722 14910 -3682
rect 14750 -3792 14910 -3722
rect 14750 -3832 14800 -3792
rect 14770 -3852 14800 -3832
rect 14860 -3832 14910 -3792
rect 14860 -3852 14890 -3832
rect 14970 -3892 15030 -3632
rect 14630 -3902 14710 -3892
rect 14630 -3962 14640 -3902
rect 14700 -3912 14710 -3902
rect 14950 -3902 15030 -3892
rect 14950 -3912 14960 -3902
rect 14700 -3962 14960 -3912
rect 15020 -3962 15030 -3902
rect 14630 -3972 15030 -3962
rect 15086 -3552 15486 -3542
rect 15086 -3612 15096 -3552
rect 15156 -3602 15416 -3552
rect 15156 -3612 15166 -3602
rect 15086 -3622 15166 -3612
rect 15406 -3612 15416 -3602
rect 15476 -3612 15486 -3552
rect 15406 -3622 15486 -3612
rect 15086 -3892 15146 -3622
rect 15416 -3632 15486 -3622
rect 15226 -3682 15256 -3662
rect 15206 -3722 15256 -3682
rect 15316 -3682 15346 -3662
rect 15316 -3722 15366 -3682
rect 15206 -3792 15366 -3722
rect 15206 -3832 15256 -3792
rect 15226 -3852 15256 -3832
rect 15316 -3832 15366 -3792
rect 15316 -3852 15346 -3832
rect 15426 -3892 15486 -3632
rect 15086 -3902 15166 -3892
rect 15086 -3962 15096 -3902
rect 15156 -3912 15166 -3902
rect 15406 -3902 15486 -3892
rect 15406 -3912 15416 -3902
rect 15156 -3962 15416 -3912
rect 15476 -3962 15486 -3902
rect 15086 -3972 15486 -3962
rect 0 -4044 400 -4034
rect 0 -4104 10 -4044
rect 70 -4094 330 -4044
rect 70 -4104 80 -4094
rect 0 -4114 80 -4104
rect 320 -4104 330 -4094
rect 390 -4104 400 -4044
rect 320 -4114 400 -4104
rect 0 -4384 60 -4114
rect 330 -4124 400 -4114
rect 140 -4174 170 -4154
rect 120 -4214 170 -4174
rect 230 -4174 260 -4154
rect 230 -4214 280 -4174
rect 120 -4284 280 -4214
rect 120 -4324 170 -4284
rect 140 -4344 170 -4324
rect 230 -4324 280 -4284
rect 230 -4344 260 -4324
rect 340 -4384 400 -4124
rect 0 -4394 80 -4384
rect 0 -4454 10 -4394
rect 70 -4404 80 -4394
rect 320 -4394 400 -4384
rect 320 -4404 330 -4394
rect 70 -4454 330 -4404
rect 390 -4454 400 -4394
rect 0 -4464 400 -4454
rect 456 -4044 856 -4034
rect 456 -4104 466 -4044
rect 526 -4094 786 -4044
rect 526 -4104 536 -4094
rect 456 -4114 536 -4104
rect 776 -4104 786 -4094
rect 846 -4104 856 -4044
rect 776 -4114 856 -4104
rect 456 -4384 516 -4114
rect 786 -4124 856 -4114
rect 596 -4174 626 -4154
rect 576 -4214 626 -4174
rect 686 -4174 716 -4154
rect 686 -4214 736 -4174
rect 576 -4284 736 -4214
rect 576 -4324 626 -4284
rect 596 -4344 626 -4324
rect 686 -4324 736 -4284
rect 686 -4344 716 -4324
rect 796 -4384 856 -4124
rect 456 -4394 536 -4384
rect 456 -4454 466 -4394
rect 526 -4404 536 -4394
rect 776 -4394 856 -4384
rect 776 -4404 786 -4394
rect 526 -4454 786 -4404
rect 846 -4454 856 -4394
rect 456 -4464 856 -4454
rect 912 -4044 1312 -4034
rect 912 -4104 922 -4044
rect 982 -4094 1242 -4044
rect 982 -4104 992 -4094
rect 912 -4114 992 -4104
rect 1232 -4104 1242 -4094
rect 1302 -4104 1312 -4044
rect 1232 -4114 1312 -4104
rect 912 -4384 972 -4114
rect 1242 -4124 1312 -4114
rect 1052 -4174 1082 -4154
rect 1032 -4214 1082 -4174
rect 1142 -4174 1172 -4154
rect 1142 -4214 1192 -4174
rect 1032 -4284 1192 -4214
rect 1032 -4324 1082 -4284
rect 1052 -4344 1082 -4324
rect 1142 -4324 1192 -4284
rect 1142 -4344 1172 -4324
rect 1252 -4384 1312 -4124
rect 912 -4394 992 -4384
rect 912 -4454 922 -4394
rect 982 -4404 992 -4394
rect 1232 -4394 1312 -4384
rect 1232 -4404 1242 -4394
rect 982 -4454 1242 -4404
rect 1302 -4454 1312 -4394
rect 912 -4464 1312 -4454
rect 1370 -4044 1770 -4034
rect 1370 -4104 1380 -4044
rect 1440 -4094 1700 -4044
rect 1440 -4104 1450 -4094
rect 1370 -4114 1450 -4104
rect 1690 -4104 1700 -4094
rect 1760 -4104 1770 -4044
rect 1690 -4114 1770 -4104
rect 1370 -4384 1430 -4114
rect 1700 -4124 1770 -4114
rect 1510 -4174 1540 -4154
rect 1490 -4214 1540 -4174
rect 1600 -4174 1630 -4154
rect 1600 -4214 1650 -4174
rect 1490 -4284 1650 -4214
rect 1490 -4324 1540 -4284
rect 1510 -4344 1540 -4324
rect 1600 -4324 1650 -4284
rect 1600 -4344 1630 -4324
rect 1710 -4384 1770 -4124
rect 1370 -4394 1450 -4384
rect 1370 -4454 1380 -4394
rect 1440 -4404 1450 -4394
rect 1690 -4394 1770 -4384
rect 1690 -4404 1700 -4394
rect 1440 -4454 1700 -4404
rect 1760 -4454 1770 -4394
rect 1370 -4464 1770 -4454
rect 1826 -4044 2226 -4034
rect 1826 -4104 1836 -4044
rect 1896 -4094 2156 -4044
rect 1896 -4104 1906 -4094
rect 1826 -4114 1906 -4104
rect 2146 -4104 2156 -4094
rect 2216 -4104 2226 -4044
rect 2146 -4114 2226 -4104
rect 1826 -4384 1886 -4114
rect 2156 -4124 2226 -4114
rect 1966 -4174 1996 -4154
rect 1946 -4214 1996 -4174
rect 2056 -4174 2086 -4154
rect 2056 -4214 2106 -4174
rect 1946 -4284 2106 -4214
rect 1946 -4324 1996 -4284
rect 1966 -4344 1996 -4324
rect 2056 -4324 2106 -4284
rect 2056 -4344 2086 -4324
rect 2166 -4384 2226 -4124
rect 1826 -4394 1906 -4384
rect 1826 -4454 1836 -4394
rect 1896 -4404 1906 -4394
rect 2146 -4394 2226 -4384
rect 2146 -4404 2156 -4394
rect 1896 -4454 2156 -4404
rect 2216 -4454 2226 -4394
rect 1826 -4464 2226 -4454
rect 2282 -4044 2682 -4034
rect 2282 -4104 2292 -4044
rect 2352 -4094 2612 -4044
rect 2352 -4104 2362 -4094
rect 2282 -4114 2362 -4104
rect 2602 -4104 2612 -4094
rect 2672 -4104 2682 -4044
rect 2602 -4114 2682 -4104
rect 2282 -4384 2342 -4114
rect 2612 -4124 2682 -4114
rect 2422 -4174 2452 -4154
rect 2402 -4214 2452 -4174
rect 2512 -4174 2542 -4154
rect 2512 -4214 2562 -4174
rect 2402 -4284 2562 -4214
rect 2402 -4324 2452 -4284
rect 2422 -4344 2452 -4324
rect 2512 -4324 2562 -4284
rect 2512 -4344 2542 -4324
rect 2622 -4384 2682 -4124
rect 2282 -4394 2362 -4384
rect 2282 -4454 2292 -4394
rect 2352 -4404 2362 -4394
rect 2602 -4394 2682 -4384
rect 2602 -4404 2612 -4394
rect 2352 -4454 2612 -4404
rect 2672 -4454 2682 -4394
rect 2282 -4464 2682 -4454
rect 2740 -4044 3140 -4034
rect 2740 -4104 2750 -4044
rect 2810 -4094 3070 -4044
rect 2810 -4104 2820 -4094
rect 2740 -4114 2820 -4104
rect 3060 -4104 3070 -4094
rect 3130 -4104 3140 -4044
rect 3060 -4114 3140 -4104
rect 2740 -4384 2800 -4114
rect 3070 -4124 3140 -4114
rect 2880 -4174 2910 -4154
rect 2860 -4214 2910 -4174
rect 2970 -4174 3000 -4154
rect 2970 -4214 3020 -4174
rect 2860 -4284 3020 -4214
rect 2860 -4324 2910 -4284
rect 2880 -4344 2910 -4324
rect 2970 -4324 3020 -4284
rect 2970 -4344 3000 -4324
rect 3080 -4384 3140 -4124
rect 2740 -4394 2820 -4384
rect 2740 -4454 2750 -4394
rect 2810 -4404 2820 -4394
rect 3060 -4394 3140 -4384
rect 3060 -4404 3070 -4394
rect 2810 -4454 3070 -4404
rect 3130 -4454 3140 -4394
rect 2740 -4464 3140 -4454
rect 3196 -4044 3596 -4034
rect 3196 -4104 3206 -4044
rect 3266 -4094 3526 -4044
rect 3266 -4104 3276 -4094
rect 3196 -4114 3276 -4104
rect 3516 -4104 3526 -4094
rect 3586 -4104 3596 -4044
rect 3516 -4114 3596 -4104
rect 3196 -4384 3256 -4114
rect 3526 -4124 3596 -4114
rect 3336 -4174 3366 -4154
rect 3316 -4214 3366 -4174
rect 3426 -4174 3456 -4154
rect 3426 -4214 3476 -4174
rect 3316 -4284 3476 -4214
rect 3316 -4324 3366 -4284
rect 3336 -4344 3366 -4324
rect 3426 -4324 3476 -4284
rect 3426 -4344 3456 -4324
rect 3536 -4384 3596 -4124
rect 3196 -4394 3276 -4384
rect 3196 -4454 3206 -4394
rect 3266 -4404 3276 -4394
rect 3516 -4394 3596 -4384
rect 3516 -4404 3526 -4394
rect 3266 -4454 3526 -4404
rect 3586 -4454 3596 -4394
rect 3196 -4464 3596 -4454
rect 3652 -4044 4052 -4034
rect 3652 -4104 3662 -4044
rect 3722 -4094 3982 -4044
rect 3722 -4104 3732 -4094
rect 3652 -4114 3732 -4104
rect 3972 -4104 3982 -4094
rect 4042 -4104 4052 -4044
rect 3972 -4114 4052 -4104
rect 3652 -4384 3712 -4114
rect 3982 -4124 4052 -4114
rect 3792 -4174 3822 -4154
rect 3772 -4214 3822 -4174
rect 3882 -4174 3912 -4154
rect 3882 -4214 3932 -4174
rect 3772 -4284 3932 -4214
rect 3772 -4324 3822 -4284
rect 3792 -4344 3822 -4324
rect 3882 -4324 3932 -4284
rect 3882 -4344 3912 -4324
rect 3992 -4384 4052 -4124
rect 3652 -4394 3732 -4384
rect 3652 -4454 3662 -4394
rect 3722 -4404 3732 -4394
rect 3972 -4394 4052 -4384
rect 3972 -4404 3982 -4394
rect 3722 -4454 3982 -4404
rect 4042 -4454 4052 -4394
rect 3652 -4464 4052 -4454
rect 4110 -4044 4510 -4034
rect 4110 -4104 4120 -4044
rect 4180 -4094 4440 -4044
rect 4180 -4104 4190 -4094
rect 4110 -4114 4190 -4104
rect 4430 -4104 4440 -4094
rect 4500 -4104 4510 -4044
rect 4430 -4114 4510 -4104
rect 4110 -4384 4170 -4114
rect 4440 -4124 4510 -4114
rect 4250 -4174 4280 -4154
rect 4230 -4214 4280 -4174
rect 4340 -4174 4370 -4154
rect 4340 -4214 4390 -4174
rect 4230 -4284 4390 -4214
rect 4230 -4324 4280 -4284
rect 4250 -4344 4280 -4324
rect 4340 -4324 4390 -4284
rect 4340 -4344 4370 -4324
rect 4450 -4384 4510 -4124
rect 4110 -4394 4190 -4384
rect 4110 -4454 4120 -4394
rect 4180 -4404 4190 -4394
rect 4430 -4394 4510 -4384
rect 4430 -4404 4440 -4394
rect 4180 -4454 4440 -4404
rect 4500 -4454 4510 -4394
rect 4110 -4464 4510 -4454
rect 4566 -4044 4966 -4034
rect 4566 -4104 4576 -4044
rect 4636 -4094 4896 -4044
rect 4636 -4104 4646 -4094
rect 4566 -4114 4646 -4104
rect 4886 -4104 4896 -4094
rect 4956 -4104 4966 -4044
rect 4886 -4114 4966 -4104
rect 4566 -4384 4626 -4114
rect 4896 -4124 4966 -4114
rect 4706 -4174 4736 -4154
rect 4686 -4214 4736 -4174
rect 4796 -4174 4826 -4154
rect 4796 -4214 4846 -4174
rect 4686 -4284 4846 -4214
rect 4686 -4324 4736 -4284
rect 4706 -4344 4736 -4324
rect 4796 -4324 4846 -4284
rect 4796 -4344 4826 -4324
rect 4906 -4384 4966 -4124
rect 4566 -4394 4646 -4384
rect 4566 -4454 4576 -4394
rect 4636 -4404 4646 -4394
rect 4886 -4394 4966 -4384
rect 4886 -4404 4896 -4394
rect 4636 -4454 4896 -4404
rect 4956 -4454 4966 -4394
rect 4566 -4464 4966 -4454
rect 5022 -4044 5422 -4034
rect 5022 -4104 5032 -4044
rect 5092 -4094 5352 -4044
rect 5092 -4104 5102 -4094
rect 5022 -4114 5102 -4104
rect 5342 -4104 5352 -4094
rect 5412 -4104 5422 -4044
rect 5342 -4114 5422 -4104
rect 5022 -4384 5082 -4114
rect 5352 -4124 5422 -4114
rect 5162 -4174 5192 -4154
rect 5142 -4214 5192 -4174
rect 5252 -4174 5282 -4154
rect 5252 -4214 5302 -4174
rect 5142 -4284 5302 -4214
rect 5142 -4324 5192 -4284
rect 5162 -4344 5192 -4324
rect 5252 -4324 5302 -4284
rect 5252 -4344 5282 -4324
rect 5362 -4384 5422 -4124
rect 5022 -4394 5102 -4384
rect 5022 -4454 5032 -4394
rect 5092 -4404 5102 -4394
rect 5342 -4394 5422 -4384
rect 5342 -4404 5352 -4394
rect 5092 -4454 5352 -4404
rect 5412 -4454 5422 -4394
rect 5022 -4464 5422 -4454
rect 5480 -4044 5880 -4034
rect 5480 -4104 5490 -4044
rect 5550 -4094 5810 -4044
rect 5550 -4104 5560 -4094
rect 5480 -4114 5560 -4104
rect 5800 -4104 5810 -4094
rect 5870 -4104 5880 -4044
rect 5800 -4114 5880 -4104
rect 5480 -4384 5540 -4114
rect 5810 -4124 5880 -4114
rect 5620 -4174 5650 -4154
rect 5600 -4214 5650 -4174
rect 5710 -4174 5740 -4154
rect 5710 -4214 5760 -4174
rect 5600 -4284 5760 -4214
rect 5600 -4324 5650 -4284
rect 5620 -4344 5650 -4324
rect 5710 -4324 5760 -4284
rect 5710 -4344 5740 -4324
rect 5820 -4384 5880 -4124
rect 5480 -4394 5560 -4384
rect 5480 -4454 5490 -4394
rect 5550 -4404 5560 -4394
rect 5800 -4394 5880 -4384
rect 5800 -4404 5810 -4394
rect 5550 -4454 5810 -4404
rect 5870 -4454 5880 -4394
rect 5480 -4464 5880 -4454
rect 5936 -4044 6336 -4034
rect 5936 -4104 5946 -4044
rect 6006 -4094 6266 -4044
rect 6006 -4104 6016 -4094
rect 5936 -4114 6016 -4104
rect 6256 -4104 6266 -4094
rect 6326 -4104 6336 -4044
rect 6256 -4114 6336 -4104
rect 5936 -4384 5996 -4114
rect 6266 -4124 6336 -4114
rect 6076 -4174 6106 -4154
rect 6056 -4214 6106 -4174
rect 6166 -4174 6196 -4154
rect 6166 -4214 6216 -4174
rect 6056 -4284 6216 -4214
rect 6056 -4324 6106 -4284
rect 6076 -4344 6106 -4324
rect 6166 -4324 6216 -4284
rect 6166 -4344 6196 -4324
rect 6276 -4384 6336 -4124
rect 5936 -4394 6016 -4384
rect 5936 -4454 5946 -4394
rect 6006 -4404 6016 -4394
rect 6256 -4394 6336 -4384
rect 6256 -4404 6266 -4394
rect 6006 -4454 6266 -4404
rect 6326 -4454 6336 -4394
rect 5936 -4464 6336 -4454
rect 6392 -4044 6792 -4034
rect 6392 -4104 6402 -4044
rect 6462 -4094 6722 -4044
rect 6462 -4104 6472 -4094
rect 6392 -4114 6472 -4104
rect 6712 -4104 6722 -4094
rect 6782 -4104 6792 -4044
rect 6712 -4114 6792 -4104
rect 6392 -4384 6452 -4114
rect 6722 -4124 6792 -4114
rect 6532 -4174 6562 -4154
rect 6512 -4214 6562 -4174
rect 6622 -4174 6652 -4154
rect 6622 -4214 6672 -4174
rect 6512 -4284 6672 -4214
rect 6512 -4324 6562 -4284
rect 6532 -4344 6562 -4324
rect 6622 -4324 6672 -4284
rect 6622 -4344 6652 -4324
rect 6732 -4384 6792 -4124
rect 6392 -4394 6472 -4384
rect 6392 -4454 6402 -4394
rect 6462 -4404 6472 -4394
rect 6712 -4394 6792 -4384
rect 6712 -4404 6722 -4394
rect 6462 -4454 6722 -4404
rect 6782 -4454 6792 -4394
rect 6392 -4464 6792 -4454
rect 6850 -4044 7250 -4034
rect 6850 -4104 6860 -4044
rect 6920 -4094 7180 -4044
rect 6920 -4104 6930 -4094
rect 6850 -4114 6930 -4104
rect 7170 -4104 7180 -4094
rect 7240 -4104 7250 -4044
rect 7170 -4114 7250 -4104
rect 6850 -4384 6910 -4114
rect 7180 -4124 7250 -4114
rect 6990 -4174 7020 -4154
rect 6970 -4214 7020 -4174
rect 7080 -4174 7110 -4154
rect 7080 -4214 7130 -4174
rect 6970 -4284 7130 -4214
rect 6970 -4324 7020 -4284
rect 6990 -4344 7020 -4324
rect 7080 -4324 7130 -4284
rect 7080 -4344 7110 -4324
rect 7190 -4384 7250 -4124
rect 6850 -4394 6930 -4384
rect 6850 -4454 6860 -4394
rect 6920 -4404 6930 -4394
rect 7170 -4394 7250 -4384
rect 7170 -4404 7180 -4394
rect 6920 -4454 7180 -4404
rect 7240 -4454 7250 -4394
rect 6850 -4464 7250 -4454
rect 7306 -4044 7706 -4034
rect 7306 -4104 7316 -4044
rect 7376 -4094 7636 -4044
rect 7376 -4104 7386 -4094
rect 7306 -4114 7386 -4104
rect 7626 -4104 7636 -4094
rect 7696 -4104 7706 -4044
rect 7626 -4114 7706 -4104
rect 7306 -4384 7366 -4114
rect 7636 -4124 7706 -4114
rect 7446 -4174 7476 -4154
rect 7426 -4214 7476 -4174
rect 7536 -4174 7566 -4154
rect 7536 -4214 7586 -4174
rect 7426 -4284 7586 -4214
rect 7426 -4324 7476 -4284
rect 7446 -4344 7476 -4324
rect 7536 -4324 7586 -4284
rect 7536 -4344 7566 -4324
rect 7646 -4384 7706 -4124
rect 7306 -4394 7386 -4384
rect 7306 -4454 7316 -4394
rect 7376 -4404 7386 -4394
rect 7626 -4394 7706 -4384
rect 7626 -4404 7636 -4394
rect 7376 -4454 7636 -4404
rect 7696 -4454 7706 -4394
rect 7306 -4464 7706 -4454
rect 7762 -4044 8162 -4034
rect 7762 -4104 7772 -4044
rect 7832 -4094 8092 -4044
rect 7832 -4104 7842 -4094
rect 7762 -4114 7842 -4104
rect 8082 -4104 8092 -4094
rect 8152 -4104 8162 -4044
rect 8082 -4114 8162 -4104
rect 7762 -4384 7822 -4114
rect 8092 -4124 8162 -4114
rect 7902 -4174 7932 -4154
rect 7882 -4214 7932 -4174
rect 7992 -4174 8022 -4154
rect 7992 -4214 8042 -4174
rect 7882 -4284 8042 -4214
rect 7882 -4324 7932 -4284
rect 7902 -4344 7932 -4324
rect 7992 -4324 8042 -4284
rect 7992 -4344 8022 -4324
rect 8102 -4384 8162 -4124
rect 7762 -4394 7842 -4384
rect 7762 -4454 7772 -4394
rect 7832 -4404 7842 -4394
rect 8082 -4394 8162 -4384
rect 8082 -4404 8092 -4394
rect 7832 -4454 8092 -4404
rect 8152 -4454 8162 -4394
rect 7762 -4464 8162 -4454
rect 8236 -4044 8636 -4034
rect 8236 -4104 8246 -4044
rect 8306 -4094 8566 -4044
rect 8306 -4104 8316 -4094
rect 8236 -4114 8316 -4104
rect 8556 -4104 8566 -4094
rect 8626 -4104 8636 -4044
rect 8556 -4114 8636 -4104
rect 8236 -4384 8296 -4114
rect 8566 -4124 8636 -4114
rect 8376 -4174 8406 -4154
rect 8356 -4214 8406 -4174
rect 8466 -4174 8496 -4154
rect 8466 -4214 8516 -4174
rect 8356 -4284 8516 -4214
rect 8356 -4324 8406 -4284
rect 8376 -4344 8406 -4324
rect 8466 -4324 8516 -4284
rect 8466 -4344 8496 -4324
rect 8576 -4384 8636 -4124
rect 8236 -4394 8316 -4384
rect 8236 -4454 8246 -4394
rect 8306 -4404 8316 -4394
rect 8556 -4394 8636 -4384
rect 8556 -4404 8566 -4394
rect 8306 -4454 8566 -4404
rect 8626 -4454 8636 -4394
rect 8236 -4464 8636 -4454
rect 8692 -4044 9092 -4034
rect 8692 -4104 8702 -4044
rect 8762 -4094 9022 -4044
rect 8762 -4104 8772 -4094
rect 8692 -4114 8772 -4104
rect 9012 -4104 9022 -4094
rect 9082 -4104 9092 -4044
rect 9012 -4114 9092 -4104
rect 8692 -4384 8752 -4114
rect 9022 -4124 9092 -4114
rect 8832 -4174 8862 -4154
rect 8812 -4214 8862 -4174
rect 8922 -4174 8952 -4154
rect 8922 -4214 8972 -4174
rect 8812 -4284 8972 -4214
rect 8812 -4324 8862 -4284
rect 8832 -4344 8862 -4324
rect 8922 -4324 8972 -4284
rect 8922 -4344 8952 -4324
rect 9032 -4384 9092 -4124
rect 8692 -4394 8772 -4384
rect 8692 -4454 8702 -4394
rect 8762 -4404 8772 -4394
rect 9012 -4394 9092 -4384
rect 9012 -4404 9022 -4394
rect 8762 -4454 9022 -4404
rect 9082 -4454 9092 -4394
rect 8692 -4464 9092 -4454
rect 9150 -4044 9550 -4034
rect 9150 -4104 9160 -4044
rect 9220 -4094 9480 -4044
rect 9220 -4104 9230 -4094
rect 9150 -4114 9230 -4104
rect 9470 -4104 9480 -4094
rect 9540 -4104 9550 -4044
rect 9470 -4114 9550 -4104
rect 9150 -4384 9210 -4114
rect 9480 -4124 9550 -4114
rect 9290 -4174 9320 -4154
rect 9270 -4214 9320 -4174
rect 9380 -4174 9410 -4154
rect 9380 -4214 9430 -4174
rect 9270 -4284 9430 -4214
rect 9270 -4324 9320 -4284
rect 9290 -4344 9320 -4324
rect 9380 -4324 9430 -4284
rect 9380 -4344 9410 -4324
rect 9490 -4384 9550 -4124
rect 9150 -4394 9230 -4384
rect 9150 -4454 9160 -4394
rect 9220 -4404 9230 -4394
rect 9470 -4394 9550 -4384
rect 9470 -4404 9480 -4394
rect 9220 -4454 9480 -4404
rect 9540 -4454 9550 -4394
rect 9150 -4464 9550 -4454
rect 9606 -4044 10006 -4034
rect 9606 -4104 9616 -4044
rect 9676 -4094 9936 -4044
rect 9676 -4104 9686 -4094
rect 9606 -4114 9686 -4104
rect 9926 -4104 9936 -4094
rect 9996 -4104 10006 -4044
rect 9926 -4114 10006 -4104
rect 9606 -4384 9666 -4114
rect 9936 -4124 10006 -4114
rect 9746 -4174 9776 -4154
rect 9726 -4214 9776 -4174
rect 9836 -4174 9866 -4154
rect 9836 -4214 9886 -4174
rect 9726 -4284 9886 -4214
rect 9726 -4324 9776 -4284
rect 9746 -4344 9776 -4324
rect 9836 -4324 9886 -4284
rect 9836 -4344 9866 -4324
rect 9946 -4384 10006 -4124
rect 9606 -4394 9686 -4384
rect 9606 -4454 9616 -4394
rect 9676 -4404 9686 -4394
rect 9926 -4394 10006 -4384
rect 9926 -4404 9936 -4394
rect 9676 -4454 9936 -4404
rect 9996 -4454 10006 -4394
rect 9606 -4464 10006 -4454
rect 10062 -4044 10462 -4034
rect 10062 -4104 10072 -4044
rect 10132 -4094 10392 -4044
rect 10132 -4104 10142 -4094
rect 10062 -4114 10142 -4104
rect 10382 -4104 10392 -4094
rect 10452 -4104 10462 -4044
rect 10382 -4114 10462 -4104
rect 10062 -4384 10122 -4114
rect 10392 -4124 10462 -4114
rect 10202 -4174 10232 -4154
rect 10182 -4214 10232 -4174
rect 10292 -4174 10322 -4154
rect 10292 -4214 10342 -4174
rect 10182 -4284 10342 -4214
rect 10182 -4324 10232 -4284
rect 10202 -4344 10232 -4324
rect 10292 -4324 10342 -4284
rect 10292 -4344 10322 -4324
rect 10402 -4384 10462 -4124
rect 10062 -4394 10142 -4384
rect 10062 -4454 10072 -4394
rect 10132 -4404 10142 -4394
rect 10382 -4394 10462 -4384
rect 10382 -4404 10392 -4394
rect 10132 -4454 10392 -4404
rect 10452 -4454 10462 -4394
rect 10062 -4464 10462 -4454
rect 10520 -4044 10920 -4034
rect 10520 -4104 10530 -4044
rect 10590 -4094 10850 -4044
rect 10590 -4104 10600 -4094
rect 10520 -4114 10600 -4104
rect 10840 -4104 10850 -4094
rect 10910 -4104 10920 -4044
rect 10840 -4114 10920 -4104
rect 10520 -4384 10580 -4114
rect 10850 -4124 10920 -4114
rect 10660 -4174 10690 -4154
rect 10640 -4214 10690 -4174
rect 10750 -4174 10780 -4154
rect 10750 -4214 10800 -4174
rect 10640 -4284 10800 -4214
rect 10640 -4324 10690 -4284
rect 10660 -4344 10690 -4324
rect 10750 -4324 10800 -4284
rect 10750 -4344 10780 -4324
rect 10860 -4384 10920 -4124
rect 10520 -4394 10600 -4384
rect 10520 -4454 10530 -4394
rect 10590 -4404 10600 -4394
rect 10840 -4394 10920 -4384
rect 10840 -4404 10850 -4394
rect 10590 -4454 10850 -4404
rect 10910 -4454 10920 -4394
rect 10520 -4464 10920 -4454
rect 10976 -4044 11376 -4034
rect 10976 -4104 10986 -4044
rect 11046 -4094 11306 -4044
rect 11046 -4104 11056 -4094
rect 10976 -4114 11056 -4104
rect 11296 -4104 11306 -4094
rect 11366 -4104 11376 -4044
rect 11296 -4114 11376 -4104
rect 10976 -4384 11036 -4114
rect 11306 -4124 11376 -4114
rect 11116 -4174 11146 -4154
rect 11096 -4214 11146 -4174
rect 11206 -4174 11236 -4154
rect 11206 -4214 11256 -4174
rect 11096 -4284 11256 -4214
rect 11096 -4324 11146 -4284
rect 11116 -4344 11146 -4324
rect 11206 -4324 11256 -4284
rect 11206 -4344 11236 -4324
rect 11316 -4384 11376 -4124
rect 10976 -4394 11056 -4384
rect 10976 -4454 10986 -4394
rect 11046 -4404 11056 -4394
rect 11296 -4394 11376 -4384
rect 11296 -4404 11306 -4394
rect 11046 -4454 11306 -4404
rect 11366 -4454 11376 -4394
rect 10976 -4464 11376 -4454
rect 11432 -4044 11832 -4034
rect 11432 -4104 11442 -4044
rect 11502 -4094 11762 -4044
rect 11502 -4104 11512 -4094
rect 11432 -4114 11512 -4104
rect 11752 -4104 11762 -4094
rect 11822 -4104 11832 -4044
rect 11752 -4114 11832 -4104
rect 11432 -4384 11492 -4114
rect 11762 -4124 11832 -4114
rect 11572 -4174 11602 -4154
rect 11552 -4214 11602 -4174
rect 11662 -4174 11692 -4154
rect 11662 -4214 11712 -4174
rect 11552 -4284 11712 -4214
rect 11552 -4324 11602 -4284
rect 11572 -4344 11602 -4324
rect 11662 -4324 11712 -4284
rect 11662 -4344 11692 -4324
rect 11772 -4384 11832 -4124
rect 11432 -4394 11512 -4384
rect 11432 -4454 11442 -4394
rect 11502 -4404 11512 -4394
rect 11752 -4394 11832 -4384
rect 11752 -4404 11762 -4394
rect 11502 -4454 11762 -4404
rect 11822 -4454 11832 -4394
rect 11432 -4464 11832 -4454
rect 11890 -4044 12290 -4034
rect 11890 -4104 11900 -4044
rect 11960 -4094 12220 -4044
rect 11960 -4104 11970 -4094
rect 11890 -4114 11970 -4104
rect 12210 -4104 12220 -4094
rect 12280 -4104 12290 -4044
rect 12210 -4114 12290 -4104
rect 11890 -4384 11950 -4114
rect 12220 -4124 12290 -4114
rect 12030 -4174 12060 -4154
rect 12010 -4214 12060 -4174
rect 12120 -4174 12150 -4154
rect 12120 -4214 12170 -4174
rect 12010 -4284 12170 -4214
rect 12010 -4324 12060 -4284
rect 12030 -4344 12060 -4324
rect 12120 -4324 12170 -4284
rect 12120 -4344 12150 -4324
rect 12230 -4384 12290 -4124
rect 11890 -4394 11970 -4384
rect 11890 -4454 11900 -4394
rect 11960 -4404 11970 -4394
rect 12210 -4394 12290 -4384
rect 12210 -4404 12220 -4394
rect 11960 -4454 12220 -4404
rect 12280 -4454 12290 -4394
rect 11890 -4464 12290 -4454
rect 12346 -4044 12746 -4034
rect 12346 -4104 12356 -4044
rect 12416 -4094 12676 -4044
rect 12416 -4104 12426 -4094
rect 12346 -4114 12426 -4104
rect 12666 -4104 12676 -4094
rect 12736 -4104 12746 -4044
rect 12666 -4114 12746 -4104
rect 12346 -4384 12406 -4114
rect 12676 -4124 12746 -4114
rect 12486 -4174 12516 -4154
rect 12466 -4214 12516 -4174
rect 12576 -4174 12606 -4154
rect 12576 -4214 12626 -4174
rect 12466 -4284 12626 -4214
rect 12466 -4324 12516 -4284
rect 12486 -4344 12516 -4324
rect 12576 -4324 12626 -4284
rect 12576 -4344 12606 -4324
rect 12686 -4384 12746 -4124
rect 12346 -4394 12426 -4384
rect 12346 -4454 12356 -4394
rect 12416 -4404 12426 -4394
rect 12666 -4394 12746 -4384
rect 12666 -4404 12676 -4394
rect 12416 -4454 12676 -4404
rect 12736 -4454 12746 -4394
rect 12346 -4464 12746 -4454
rect 12802 -4044 13202 -4034
rect 12802 -4104 12812 -4044
rect 12872 -4094 13132 -4044
rect 12872 -4104 12882 -4094
rect 12802 -4114 12882 -4104
rect 13122 -4104 13132 -4094
rect 13192 -4104 13202 -4044
rect 13122 -4114 13202 -4104
rect 12802 -4384 12862 -4114
rect 13132 -4124 13202 -4114
rect 12942 -4174 12972 -4154
rect 12922 -4214 12972 -4174
rect 13032 -4174 13062 -4154
rect 13032 -4214 13082 -4174
rect 12922 -4284 13082 -4214
rect 12922 -4324 12972 -4284
rect 12942 -4344 12972 -4324
rect 13032 -4324 13082 -4284
rect 13032 -4344 13062 -4324
rect 13142 -4384 13202 -4124
rect 12802 -4394 12882 -4384
rect 12802 -4454 12812 -4394
rect 12872 -4404 12882 -4394
rect 13122 -4394 13202 -4384
rect 13122 -4404 13132 -4394
rect 12872 -4454 13132 -4404
rect 13192 -4454 13202 -4394
rect 12802 -4464 13202 -4454
rect 13260 -4044 13660 -4034
rect 13260 -4104 13270 -4044
rect 13330 -4094 13590 -4044
rect 13330 -4104 13340 -4094
rect 13260 -4114 13340 -4104
rect 13580 -4104 13590 -4094
rect 13650 -4104 13660 -4044
rect 13580 -4114 13660 -4104
rect 13260 -4384 13320 -4114
rect 13590 -4124 13660 -4114
rect 13400 -4174 13430 -4154
rect 13380 -4214 13430 -4174
rect 13490 -4174 13520 -4154
rect 13490 -4214 13540 -4174
rect 13380 -4284 13540 -4214
rect 13380 -4324 13430 -4284
rect 13400 -4344 13430 -4324
rect 13490 -4324 13540 -4284
rect 13490 -4344 13520 -4324
rect 13600 -4384 13660 -4124
rect 13260 -4394 13340 -4384
rect 13260 -4454 13270 -4394
rect 13330 -4404 13340 -4394
rect 13580 -4394 13660 -4384
rect 13580 -4404 13590 -4394
rect 13330 -4454 13590 -4404
rect 13650 -4454 13660 -4394
rect 13260 -4464 13660 -4454
rect 13716 -4044 14116 -4034
rect 13716 -4104 13726 -4044
rect 13786 -4094 14046 -4044
rect 13786 -4104 13796 -4094
rect 13716 -4114 13796 -4104
rect 14036 -4104 14046 -4094
rect 14106 -4104 14116 -4044
rect 14036 -4114 14116 -4104
rect 13716 -4384 13776 -4114
rect 14046 -4124 14116 -4114
rect 13856 -4174 13886 -4154
rect 13836 -4214 13886 -4174
rect 13946 -4174 13976 -4154
rect 13946 -4214 13996 -4174
rect 13836 -4284 13996 -4214
rect 13836 -4324 13886 -4284
rect 13856 -4344 13886 -4324
rect 13946 -4324 13996 -4284
rect 13946 -4344 13976 -4324
rect 14056 -4384 14116 -4124
rect 13716 -4394 13796 -4384
rect 13716 -4454 13726 -4394
rect 13786 -4404 13796 -4394
rect 14036 -4394 14116 -4384
rect 14036 -4404 14046 -4394
rect 13786 -4454 14046 -4404
rect 14106 -4454 14116 -4394
rect 13716 -4464 14116 -4454
rect 14172 -4044 14572 -4034
rect 14172 -4104 14182 -4044
rect 14242 -4094 14502 -4044
rect 14242 -4104 14252 -4094
rect 14172 -4114 14252 -4104
rect 14492 -4104 14502 -4094
rect 14562 -4104 14572 -4044
rect 14492 -4114 14572 -4104
rect 14172 -4384 14232 -4114
rect 14502 -4124 14572 -4114
rect 14312 -4174 14342 -4154
rect 14292 -4214 14342 -4174
rect 14402 -4174 14432 -4154
rect 14402 -4214 14452 -4174
rect 14292 -4284 14452 -4214
rect 14292 -4324 14342 -4284
rect 14312 -4344 14342 -4324
rect 14402 -4324 14452 -4284
rect 14402 -4344 14432 -4324
rect 14512 -4384 14572 -4124
rect 14172 -4394 14252 -4384
rect 14172 -4454 14182 -4394
rect 14242 -4404 14252 -4394
rect 14492 -4394 14572 -4384
rect 14492 -4404 14502 -4394
rect 14242 -4454 14502 -4404
rect 14562 -4454 14572 -4394
rect 14172 -4464 14572 -4454
rect 14630 -4044 15030 -4034
rect 14630 -4104 14640 -4044
rect 14700 -4094 14960 -4044
rect 14700 -4104 14710 -4094
rect 14630 -4114 14710 -4104
rect 14950 -4104 14960 -4094
rect 15020 -4104 15030 -4044
rect 14950 -4114 15030 -4104
rect 14630 -4384 14690 -4114
rect 14960 -4124 15030 -4114
rect 14770 -4174 14800 -4154
rect 14750 -4214 14800 -4174
rect 14860 -4174 14890 -4154
rect 14860 -4214 14910 -4174
rect 14750 -4284 14910 -4214
rect 14750 -4324 14800 -4284
rect 14770 -4344 14800 -4324
rect 14860 -4324 14910 -4284
rect 14860 -4344 14890 -4324
rect 14970 -4384 15030 -4124
rect 14630 -4394 14710 -4384
rect 14630 -4454 14640 -4394
rect 14700 -4404 14710 -4394
rect 14950 -4394 15030 -4384
rect 14950 -4404 14960 -4394
rect 14700 -4454 14960 -4404
rect 15020 -4454 15030 -4394
rect 14630 -4464 15030 -4454
rect 15086 -4044 15486 -4034
rect 15086 -4104 15096 -4044
rect 15156 -4094 15416 -4044
rect 15156 -4104 15166 -4094
rect 15086 -4114 15166 -4104
rect 15406 -4104 15416 -4094
rect 15476 -4104 15486 -4044
rect 15406 -4114 15486 -4104
rect 15086 -4384 15146 -4114
rect 15416 -4124 15486 -4114
rect 15226 -4174 15256 -4154
rect 15206 -4214 15256 -4174
rect 15316 -4174 15346 -4154
rect 15316 -4214 15366 -4174
rect 15206 -4284 15366 -4214
rect 15206 -4324 15256 -4284
rect 15226 -4344 15256 -4324
rect 15316 -4324 15366 -4284
rect 15316 -4344 15346 -4324
rect 15426 -4384 15486 -4124
rect 15086 -4394 15166 -4384
rect 15086 -4454 15096 -4394
rect 15156 -4404 15166 -4394
rect 15406 -4394 15486 -4384
rect 15406 -4404 15416 -4394
rect 15156 -4454 15416 -4404
rect 15476 -4454 15486 -4394
rect 15086 -4464 15486 -4454
rect 0 -4560 400 -4550
rect 0 -4620 10 -4560
rect 70 -4610 330 -4560
rect 70 -4620 80 -4610
rect 0 -4630 80 -4620
rect 320 -4620 330 -4610
rect 390 -4620 400 -4560
rect 320 -4630 400 -4620
rect 0 -4900 60 -4630
rect 330 -4640 400 -4630
rect 140 -4690 170 -4670
rect 120 -4730 170 -4690
rect 230 -4690 260 -4670
rect 230 -4730 280 -4690
rect 120 -4800 280 -4730
rect 120 -4840 170 -4800
rect 140 -4860 170 -4840
rect 230 -4840 280 -4800
rect 230 -4860 260 -4840
rect 340 -4900 400 -4640
rect 0 -4910 80 -4900
rect 0 -4970 10 -4910
rect 70 -4920 80 -4910
rect 320 -4910 400 -4900
rect 320 -4920 330 -4910
rect 70 -4970 330 -4920
rect 390 -4970 400 -4910
rect 0 -4980 400 -4970
rect 456 -4560 856 -4550
rect 456 -4620 466 -4560
rect 526 -4610 786 -4560
rect 526 -4620 536 -4610
rect 456 -4630 536 -4620
rect 776 -4620 786 -4610
rect 846 -4620 856 -4560
rect 776 -4630 856 -4620
rect 456 -4900 516 -4630
rect 786 -4640 856 -4630
rect 596 -4690 626 -4670
rect 576 -4730 626 -4690
rect 686 -4690 716 -4670
rect 686 -4730 736 -4690
rect 576 -4800 736 -4730
rect 576 -4840 626 -4800
rect 596 -4860 626 -4840
rect 686 -4840 736 -4800
rect 686 -4860 716 -4840
rect 796 -4900 856 -4640
rect 456 -4910 536 -4900
rect 456 -4970 466 -4910
rect 526 -4920 536 -4910
rect 776 -4910 856 -4900
rect 776 -4920 786 -4910
rect 526 -4970 786 -4920
rect 846 -4970 856 -4910
rect 456 -4980 856 -4970
rect 912 -4560 1312 -4550
rect 912 -4620 922 -4560
rect 982 -4610 1242 -4560
rect 982 -4620 992 -4610
rect 912 -4630 992 -4620
rect 1232 -4620 1242 -4610
rect 1302 -4620 1312 -4560
rect 1232 -4630 1312 -4620
rect 912 -4900 972 -4630
rect 1242 -4640 1312 -4630
rect 1052 -4690 1082 -4670
rect 1032 -4730 1082 -4690
rect 1142 -4690 1172 -4670
rect 1142 -4730 1192 -4690
rect 1032 -4800 1192 -4730
rect 1032 -4840 1082 -4800
rect 1052 -4860 1082 -4840
rect 1142 -4840 1192 -4800
rect 1142 -4860 1172 -4840
rect 1252 -4900 1312 -4640
rect 912 -4910 992 -4900
rect 912 -4970 922 -4910
rect 982 -4920 992 -4910
rect 1232 -4910 1312 -4900
rect 1232 -4920 1242 -4910
rect 982 -4970 1242 -4920
rect 1302 -4970 1312 -4910
rect 912 -4980 1312 -4970
rect 1370 -4560 1770 -4550
rect 1370 -4620 1380 -4560
rect 1440 -4610 1700 -4560
rect 1440 -4620 1450 -4610
rect 1370 -4630 1450 -4620
rect 1690 -4620 1700 -4610
rect 1760 -4620 1770 -4560
rect 1690 -4630 1770 -4620
rect 1370 -4900 1430 -4630
rect 1700 -4640 1770 -4630
rect 1510 -4690 1540 -4670
rect 1490 -4730 1540 -4690
rect 1600 -4690 1630 -4670
rect 1600 -4730 1650 -4690
rect 1490 -4800 1650 -4730
rect 1490 -4840 1540 -4800
rect 1510 -4860 1540 -4840
rect 1600 -4840 1650 -4800
rect 1600 -4860 1630 -4840
rect 1710 -4900 1770 -4640
rect 1370 -4910 1450 -4900
rect 1370 -4970 1380 -4910
rect 1440 -4920 1450 -4910
rect 1690 -4910 1770 -4900
rect 1690 -4920 1700 -4910
rect 1440 -4970 1700 -4920
rect 1760 -4970 1770 -4910
rect 1370 -4980 1770 -4970
rect 1826 -4560 2226 -4550
rect 1826 -4620 1836 -4560
rect 1896 -4610 2156 -4560
rect 1896 -4620 1906 -4610
rect 1826 -4630 1906 -4620
rect 2146 -4620 2156 -4610
rect 2216 -4620 2226 -4560
rect 2146 -4630 2226 -4620
rect 1826 -4900 1886 -4630
rect 2156 -4640 2226 -4630
rect 1966 -4690 1996 -4670
rect 1946 -4730 1996 -4690
rect 2056 -4690 2086 -4670
rect 2056 -4730 2106 -4690
rect 1946 -4800 2106 -4730
rect 1946 -4840 1996 -4800
rect 1966 -4860 1996 -4840
rect 2056 -4840 2106 -4800
rect 2056 -4860 2086 -4840
rect 2166 -4900 2226 -4640
rect 1826 -4910 1906 -4900
rect 1826 -4970 1836 -4910
rect 1896 -4920 1906 -4910
rect 2146 -4910 2226 -4900
rect 2146 -4920 2156 -4910
rect 1896 -4970 2156 -4920
rect 2216 -4970 2226 -4910
rect 1826 -4980 2226 -4970
rect 2282 -4560 2682 -4550
rect 2282 -4620 2292 -4560
rect 2352 -4610 2612 -4560
rect 2352 -4620 2362 -4610
rect 2282 -4630 2362 -4620
rect 2602 -4620 2612 -4610
rect 2672 -4620 2682 -4560
rect 2602 -4630 2682 -4620
rect 2282 -4900 2342 -4630
rect 2612 -4640 2682 -4630
rect 2422 -4690 2452 -4670
rect 2402 -4730 2452 -4690
rect 2512 -4690 2542 -4670
rect 2512 -4730 2562 -4690
rect 2402 -4800 2562 -4730
rect 2402 -4840 2452 -4800
rect 2422 -4860 2452 -4840
rect 2512 -4840 2562 -4800
rect 2512 -4860 2542 -4840
rect 2622 -4900 2682 -4640
rect 2282 -4910 2362 -4900
rect 2282 -4970 2292 -4910
rect 2352 -4920 2362 -4910
rect 2602 -4910 2682 -4900
rect 2602 -4920 2612 -4910
rect 2352 -4970 2612 -4920
rect 2672 -4970 2682 -4910
rect 2282 -4980 2682 -4970
rect 2740 -4560 3140 -4550
rect 2740 -4620 2750 -4560
rect 2810 -4610 3070 -4560
rect 2810 -4620 2820 -4610
rect 2740 -4630 2820 -4620
rect 3060 -4620 3070 -4610
rect 3130 -4620 3140 -4560
rect 3060 -4630 3140 -4620
rect 2740 -4900 2800 -4630
rect 3070 -4640 3140 -4630
rect 2880 -4690 2910 -4670
rect 2860 -4730 2910 -4690
rect 2970 -4690 3000 -4670
rect 2970 -4730 3020 -4690
rect 2860 -4800 3020 -4730
rect 2860 -4840 2910 -4800
rect 2880 -4860 2910 -4840
rect 2970 -4840 3020 -4800
rect 2970 -4860 3000 -4840
rect 3080 -4900 3140 -4640
rect 2740 -4910 2820 -4900
rect 2740 -4970 2750 -4910
rect 2810 -4920 2820 -4910
rect 3060 -4910 3140 -4900
rect 3060 -4920 3070 -4910
rect 2810 -4970 3070 -4920
rect 3130 -4970 3140 -4910
rect 2740 -4980 3140 -4970
rect 3196 -4560 3596 -4550
rect 3196 -4620 3206 -4560
rect 3266 -4610 3526 -4560
rect 3266 -4620 3276 -4610
rect 3196 -4630 3276 -4620
rect 3516 -4620 3526 -4610
rect 3586 -4620 3596 -4560
rect 3516 -4630 3596 -4620
rect 3196 -4900 3256 -4630
rect 3526 -4640 3596 -4630
rect 3336 -4690 3366 -4670
rect 3316 -4730 3366 -4690
rect 3426 -4690 3456 -4670
rect 3426 -4730 3476 -4690
rect 3316 -4800 3476 -4730
rect 3316 -4840 3366 -4800
rect 3336 -4860 3366 -4840
rect 3426 -4840 3476 -4800
rect 3426 -4860 3456 -4840
rect 3536 -4900 3596 -4640
rect 3196 -4910 3276 -4900
rect 3196 -4970 3206 -4910
rect 3266 -4920 3276 -4910
rect 3516 -4910 3596 -4900
rect 3516 -4920 3526 -4910
rect 3266 -4970 3526 -4920
rect 3586 -4970 3596 -4910
rect 3196 -4980 3596 -4970
rect 3652 -4560 4052 -4550
rect 3652 -4620 3662 -4560
rect 3722 -4610 3982 -4560
rect 3722 -4620 3732 -4610
rect 3652 -4630 3732 -4620
rect 3972 -4620 3982 -4610
rect 4042 -4620 4052 -4560
rect 3972 -4630 4052 -4620
rect 3652 -4900 3712 -4630
rect 3982 -4640 4052 -4630
rect 3792 -4690 3822 -4670
rect 3772 -4730 3822 -4690
rect 3882 -4690 3912 -4670
rect 3882 -4730 3932 -4690
rect 3772 -4800 3932 -4730
rect 3772 -4840 3822 -4800
rect 3792 -4860 3822 -4840
rect 3882 -4840 3932 -4800
rect 3882 -4860 3912 -4840
rect 3992 -4900 4052 -4640
rect 3652 -4910 3732 -4900
rect 3652 -4970 3662 -4910
rect 3722 -4920 3732 -4910
rect 3972 -4910 4052 -4900
rect 3972 -4920 3982 -4910
rect 3722 -4970 3982 -4920
rect 4042 -4970 4052 -4910
rect 3652 -4980 4052 -4970
rect 4110 -4560 4510 -4550
rect 4110 -4620 4120 -4560
rect 4180 -4610 4440 -4560
rect 4180 -4620 4190 -4610
rect 4110 -4630 4190 -4620
rect 4430 -4620 4440 -4610
rect 4500 -4620 4510 -4560
rect 4430 -4630 4510 -4620
rect 4110 -4900 4170 -4630
rect 4440 -4640 4510 -4630
rect 4250 -4690 4280 -4670
rect 4230 -4730 4280 -4690
rect 4340 -4690 4370 -4670
rect 4340 -4730 4390 -4690
rect 4230 -4800 4390 -4730
rect 4230 -4840 4280 -4800
rect 4250 -4860 4280 -4840
rect 4340 -4840 4390 -4800
rect 4340 -4860 4370 -4840
rect 4450 -4900 4510 -4640
rect 4110 -4910 4190 -4900
rect 4110 -4970 4120 -4910
rect 4180 -4920 4190 -4910
rect 4430 -4910 4510 -4900
rect 4430 -4920 4440 -4910
rect 4180 -4970 4440 -4920
rect 4500 -4970 4510 -4910
rect 4110 -4980 4510 -4970
rect 4566 -4560 4966 -4550
rect 4566 -4620 4576 -4560
rect 4636 -4610 4896 -4560
rect 4636 -4620 4646 -4610
rect 4566 -4630 4646 -4620
rect 4886 -4620 4896 -4610
rect 4956 -4620 4966 -4560
rect 4886 -4630 4966 -4620
rect 4566 -4900 4626 -4630
rect 4896 -4640 4966 -4630
rect 4706 -4690 4736 -4670
rect 4686 -4730 4736 -4690
rect 4796 -4690 4826 -4670
rect 4796 -4730 4846 -4690
rect 4686 -4800 4846 -4730
rect 4686 -4840 4736 -4800
rect 4706 -4860 4736 -4840
rect 4796 -4840 4846 -4800
rect 4796 -4860 4826 -4840
rect 4906 -4900 4966 -4640
rect 4566 -4910 4646 -4900
rect 4566 -4970 4576 -4910
rect 4636 -4920 4646 -4910
rect 4886 -4910 4966 -4900
rect 4886 -4920 4896 -4910
rect 4636 -4970 4896 -4920
rect 4956 -4970 4966 -4910
rect 4566 -4980 4966 -4970
rect 5022 -4560 5422 -4550
rect 5022 -4620 5032 -4560
rect 5092 -4610 5352 -4560
rect 5092 -4620 5102 -4610
rect 5022 -4630 5102 -4620
rect 5342 -4620 5352 -4610
rect 5412 -4620 5422 -4560
rect 5342 -4630 5422 -4620
rect 5022 -4900 5082 -4630
rect 5352 -4640 5422 -4630
rect 5162 -4690 5192 -4670
rect 5142 -4730 5192 -4690
rect 5252 -4690 5282 -4670
rect 5252 -4730 5302 -4690
rect 5142 -4800 5302 -4730
rect 5142 -4840 5192 -4800
rect 5162 -4860 5192 -4840
rect 5252 -4840 5302 -4800
rect 5252 -4860 5282 -4840
rect 5362 -4900 5422 -4640
rect 5022 -4910 5102 -4900
rect 5022 -4970 5032 -4910
rect 5092 -4920 5102 -4910
rect 5342 -4910 5422 -4900
rect 5342 -4920 5352 -4910
rect 5092 -4970 5352 -4920
rect 5412 -4970 5422 -4910
rect 5022 -4980 5422 -4970
rect 5480 -4560 5880 -4550
rect 5480 -4620 5490 -4560
rect 5550 -4610 5810 -4560
rect 5550 -4620 5560 -4610
rect 5480 -4630 5560 -4620
rect 5800 -4620 5810 -4610
rect 5870 -4620 5880 -4560
rect 5800 -4630 5880 -4620
rect 5480 -4900 5540 -4630
rect 5810 -4640 5880 -4630
rect 5620 -4690 5650 -4670
rect 5600 -4730 5650 -4690
rect 5710 -4690 5740 -4670
rect 5710 -4730 5760 -4690
rect 5600 -4800 5760 -4730
rect 5600 -4840 5650 -4800
rect 5620 -4860 5650 -4840
rect 5710 -4840 5760 -4800
rect 5710 -4860 5740 -4840
rect 5820 -4900 5880 -4640
rect 5480 -4910 5560 -4900
rect 5480 -4970 5490 -4910
rect 5550 -4920 5560 -4910
rect 5800 -4910 5880 -4900
rect 5800 -4920 5810 -4910
rect 5550 -4970 5810 -4920
rect 5870 -4970 5880 -4910
rect 5480 -4980 5880 -4970
rect 5936 -4560 6336 -4550
rect 5936 -4620 5946 -4560
rect 6006 -4610 6266 -4560
rect 6006 -4620 6016 -4610
rect 5936 -4630 6016 -4620
rect 6256 -4620 6266 -4610
rect 6326 -4620 6336 -4560
rect 6256 -4630 6336 -4620
rect 5936 -4900 5996 -4630
rect 6266 -4640 6336 -4630
rect 6076 -4690 6106 -4670
rect 6056 -4730 6106 -4690
rect 6166 -4690 6196 -4670
rect 6166 -4730 6216 -4690
rect 6056 -4800 6216 -4730
rect 6056 -4840 6106 -4800
rect 6076 -4860 6106 -4840
rect 6166 -4840 6216 -4800
rect 6166 -4860 6196 -4840
rect 6276 -4900 6336 -4640
rect 5936 -4910 6016 -4900
rect 5936 -4970 5946 -4910
rect 6006 -4920 6016 -4910
rect 6256 -4910 6336 -4900
rect 6256 -4920 6266 -4910
rect 6006 -4970 6266 -4920
rect 6326 -4970 6336 -4910
rect 5936 -4980 6336 -4970
rect 6392 -4560 6792 -4550
rect 6392 -4620 6402 -4560
rect 6462 -4610 6722 -4560
rect 6462 -4620 6472 -4610
rect 6392 -4630 6472 -4620
rect 6712 -4620 6722 -4610
rect 6782 -4620 6792 -4560
rect 6712 -4630 6792 -4620
rect 6392 -4900 6452 -4630
rect 6722 -4640 6792 -4630
rect 6532 -4690 6562 -4670
rect 6512 -4730 6562 -4690
rect 6622 -4690 6652 -4670
rect 6622 -4730 6672 -4690
rect 6512 -4800 6672 -4730
rect 6512 -4840 6562 -4800
rect 6532 -4860 6562 -4840
rect 6622 -4840 6672 -4800
rect 6622 -4860 6652 -4840
rect 6732 -4900 6792 -4640
rect 6392 -4910 6472 -4900
rect 6392 -4970 6402 -4910
rect 6462 -4920 6472 -4910
rect 6712 -4910 6792 -4900
rect 6712 -4920 6722 -4910
rect 6462 -4970 6722 -4920
rect 6782 -4970 6792 -4910
rect 6392 -4980 6792 -4970
rect 6850 -4560 7250 -4550
rect 6850 -4620 6860 -4560
rect 6920 -4610 7180 -4560
rect 6920 -4620 6930 -4610
rect 6850 -4630 6930 -4620
rect 7170 -4620 7180 -4610
rect 7240 -4620 7250 -4560
rect 7170 -4630 7250 -4620
rect 6850 -4900 6910 -4630
rect 7180 -4640 7250 -4630
rect 6990 -4690 7020 -4670
rect 6970 -4730 7020 -4690
rect 7080 -4690 7110 -4670
rect 7080 -4730 7130 -4690
rect 6970 -4800 7130 -4730
rect 6970 -4840 7020 -4800
rect 6990 -4860 7020 -4840
rect 7080 -4840 7130 -4800
rect 7080 -4860 7110 -4840
rect 7190 -4900 7250 -4640
rect 6850 -4910 6930 -4900
rect 6850 -4970 6860 -4910
rect 6920 -4920 6930 -4910
rect 7170 -4910 7250 -4900
rect 7170 -4920 7180 -4910
rect 6920 -4970 7180 -4920
rect 7240 -4970 7250 -4910
rect 6850 -4980 7250 -4970
rect 7306 -4560 7706 -4550
rect 7306 -4620 7316 -4560
rect 7376 -4610 7636 -4560
rect 7376 -4620 7386 -4610
rect 7306 -4630 7386 -4620
rect 7626 -4620 7636 -4610
rect 7696 -4620 7706 -4560
rect 7626 -4630 7706 -4620
rect 7306 -4900 7366 -4630
rect 7636 -4640 7706 -4630
rect 7446 -4690 7476 -4670
rect 7426 -4730 7476 -4690
rect 7536 -4690 7566 -4670
rect 7536 -4730 7586 -4690
rect 7426 -4800 7586 -4730
rect 7426 -4840 7476 -4800
rect 7446 -4860 7476 -4840
rect 7536 -4840 7586 -4800
rect 7536 -4860 7566 -4840
rect 7646 -4900 7706 -4640
rect 7306 -4910 7386 -4900
rect 7306 -4970 7316 -4910
rect 7376 -4920 7386 -4910
rect 7626 -4910 7706 -4900
rect 7626 -4920 7636 -4910
rect 7376 -4970 7636 -4920
rect 7696 -4970 7706 -4910
rect 7306 -4980 7706 -4970
rect 7762 -4560 8162 -4550
rect 7762 -4620 7772 -4560
rect 7832 -4610 8092 -4560
rect 7832 -4620 7842 -4610
rect 7762 -4630 7842 -4620
rect 8082 -4620 8092 -4610
rect 8152 -4620 8162 -4560
rect 8082 -4630 8162 -4620
rect 7762 -4900 7822 -4630
rect 8092 -4640 8162 -4630
rect 7902 -4690 7932 -4670
rect 7882 -4730 7932 -4690
rect 7992 -4690 8022 -4670
rect 7992 -4730 8042 -4690
rect 7882 -4800 8042 -4730
rect 7882 -4840 7932 -4800
rect 7902 -4860 7932 -4840
rect 7992 -4840 8042 -4800
rect 7992 -4860 8022 -4840
rect 8102 -4900 8162 -4640
rect 7762 -4910 7842 -4900
rect 7762 -4970 7772 -4910
rect 7832 -4920 7842 -4910
rect 8082 -4910 8162 -4900
rect 8082 -4920 8092 -4910
rect 7832 -4970 8092 -4920
rect 8152 -4970 8162 -4910
rect 7762 -4980 8162 -4970
rect 8236 -4560 8636 -4550
rect 8236 -4620 8246 -4560
rect 8306 -4610 8566 -4560
rect 8306 -4620 8316 -4610
rect 8236 -4630 8316 -4620
rect 8556 -4620 8566 -4610
rect 8626 -4620 8636 -4560
rect 8556 -4630 8636 -4620
rect 8236 -4900 8296 -4630
rect 8566 -4640 8636 -4630
rect 8376 -4690 8406 -4670
rect 8356 -4730 8406 -4690
rect 8466 -4690 8496 -4670
rect 8466 -4730 8516 -4690
rect 8356 -4800 8516 -4730
rect 8356 -4840 8406 -4800
rect 8376 -4860 8406 -4840
rect 8466 -4840 8516 -4800
rect 8466 -4860 8496 -4840
rect 8576 -4900 8636 -4640
rect 8236 -4910 8316 -4900
rect 8236 -4970 8246 -4910
rect 8306 -4920 8316 -4910
rect 8556 -4910 8636 -4900
rect 8556 -4920 8566 -4910
rect 8306 -4970 8566 -4920
rect 8626 -4970 8636 -4910
rect 8236 -4980 8636 -4970
rect 8692 -4560 9092 -4550
rect 8692 -4620 8702 -4560
rect 8762 -4610 9022 -4560
rect 8762 -4620 8772 -4610
rect 8692 -4630 8772 -4620
rect 9012 -4620 9022 -4610
rect 9082 -4620 9092 -4560
rect 9012 -4630 9092 -4620
rect 8692 -4900 8752 -4630
rect 9022 -4640 9092 -4630
rect 8832 -4690 8862 -4670
rect 8812 -4730 8862 -4690
rect 8922 -4690 8952 -4670
rect 8922 -4730 8972 -4690
rect 8812 -4800 8972 -4730
rect 8812 -4840 8862 -4800
rect 8832 -4860 8862 -4840
rect 8922 -4840 8972 -4800
rect 8922 -4860 8952 -4840
rect 9032 -4900 9092 -4640
rect 8692 -4910 8772 -4900
rect 8692 -4970 8702 -4910
rect 8762 -4920 8772 -4910
rect 9012 -4910 9092 -4900
rect 9012 -4920 9022 -4910
rect 8762 -4970 9022 -4920
rect 9082 -4970 9092 -4910
rect 8692 -4980 9092 -4970
rect 9150 -4560 9550 -4550
rect 9150 -4620 9160 -4560
rect 9220 -4610 9480 -4560
rect 9220 -4620 9230 -4610
rect 9150 -4630 9230 -4620
rect 9470 -4620 9480 -4610
rect 9540 -4620 9550 -4560
rect 9470 -4630 9550 -4620
rect 9150 -4900 9210 -4630
rect 9480 -4640 9550 -4630
rect 9290 -4690 9320 -4670
rect 9270 -4730 9320 -4690
rect 9380 -4690 9410 -4670
rect 9380 -4730 9430 -4690
rect 9270 -4800 9430 -4730
rect 9270 -4840 9320 -4800
rect 9290 -4860 9320 -4840
rect 9380 -4840 9430 -4800
rect 9380 -4860 9410 -4840
rect 9490 -4900 9550 -4640
rect 9150 -4910 9230 -4900
rect 9150 -4970 9160 -4910
rect 9220 -4920 9230 -4910
rect 9470 -4910 9550 -4900
rect 9470 -4920 9480 -4910
rect 9220 -4970 9480 -4920
rect 9540 -4970 9550 -4910
rect 9150 -4980 9550 -4970
rect 9606 -4560 10006 -4550
rect 9606 -4620 9616 -4560
rect 9676 -4610 9936 -4560
rect 9676 -4620 9686 -4610
rect 9606 -4630 9686 -4620
rect 9926 -4620 9936 -4610
rect 9996 -4620 10006 -4560
rect 9926 -4630 10006 -4620
rect 9606 -4900 9666 -4630
rect 9936 -4640 10006 -4630
rect 9746 -4690 9776 -4670
rect 9726 -4730 9776 -4690
rect 9836 -4690 9866 -4670
rect 9836 -4730 9886 -4690
rect 9726 -4800 9886 -4730
rect 9726 -4840 9776 -4800
rect 9746 -4860 9776 -4840
rect 9836 -4840 9886 -4800
rect 9836 -4860 9866 -4840
rect 9946 -4900 10006 -4640
rect 9606 -4910 9686 -4900
rect 9606 -4970 9616 -4910
rect 9676 -4920 9686 -4910
rect 9926 -4910 10006 -4900
rect 9926 -4920 9936 -4910
rect 9676 -4970 9936 -4920
rect 9996 -4970 10006 -4910
rect 9606 -4980 10006 -4970
rect 10062 -4560 10462 -4550
rect 10062 -4620 10072 -4560
rect 10132 -4610 10392 -4560
rect 10132 -4620 10142 -4610
rect 10062 -4630 10142 -4620
rect 10382 -4620 10392 -4610
rect 10452 -4620 10462 -4560
rect 10382 -4630 10462 -4620
rect 10062 -4900 10122 -4630
rect 10392 -4640 10462 -4630
rect 10202 -4690 10232 -4670
rect 10182 -4730 10232 -4690
rect 10292 -4690 10322 -4670
rect 10292 -4730 10342 -4690
rect 10182 -4800 10342 -4730
rect 10182 -4840 10232 -4800
rect 10202 -4860 10232 -4840
rect 10292 -4840 10342 -4800
rect 10292 -4860 10322 -4840
rect 10402 -4900 10462 -4640
rect 10062 -4910 10142 -4900
rect 10062 -4970 10072 -4910
rect 10132 -4920 10142 -4910
rect 10382 -4910 10462 -4900
rect 10382 -4920 10392 -4910
rect 10132 -4970 10392 -4920
rect 10452 -4970 10462 -4910
rect 10062 -4980 10462 -4970
rect 10520 -4560 10920 -4550
rect 10520 -4620 10530 -4560
rect 10590 -4610 10850 -4560
rect 10590 -4620 10600 -4610
rect 10520 -4630 10600 -4620
rect 10840 -4620 10850 -4610
rect 10910 -4620 10920 -4560
rect 10840 -4630 10920 -4620
rect 10520 -4900 10580 -4630
rect 10850 -4640 10920 -4630
rect 10660 -4690 10690 -4670
rect 10640 -4730 10690 -4690
rect 10750 -4690 10780 -4670
rect 10750 -4730 10800 -4690
rect 10640 -4800 10800 -4730
rect 10640 -4840 10690 -4800
rect 10660 -4860 10690 -4840
rect 10750 -4840 10800 -4800
rect 10750 -4860 10780 -4840
rect 10860 -4900 10920 -4640
rect 10520 -4910 10600 -4900
rect 10520 -4970 10530 -4910
rect 10590 -4920 10600 -4910
rect 10840 -4910 10920 -4900
rect 10840 -4920 10850 -4910
rect 10590 -4970 10850 -4920
rect 10910 -4970 10920 -4910
rect 10520 -4980 10920 -4970
rect 10976 -4560 11376 -4550
rect 10976 -4620 10986 -4560
rect 11046 -4610 11306 -4560
rect 11046 -4620 11056 -4610
rect 10976 -4630 11056 -4620
rect 11296 -4620 11306 -4610
rect 11366 -4620 11376 -4560
rect 11296 -4630 11376 -4620
rect 10976 -4900 11036 -4630
rect 11306 -4640 11376 -4630
rect 11116 -4690 11146 -4670
rect 11096 -4730 11146 -4690
rect 11206 -4690 11236 -4670
rect 11206 -4730 11256 -4690
rect 11096 -4800 11256 -4730
rect 11096 -4840 11146 -4800
rect 11116 -4860 11146 -4840
rect 11206 -4840 11256 -4800
rect 11206 -4860 11236 -4840
rect 11316 -4900 11376 -4640
rect 10976 -4910 11056 -4900
rect 10976 -4970 10986 -4910
rect 11046 -4920 11056 -4910
rect 11296 -4910 11376 -4900
rect 11296 -4920 11306 -4910
rect 11046 -4970 11306 -4920
rect 11366 -4970 11376 -4910
rect 10976 -4980 11376 -4970
rect 11432 -4560 11832 -4550
rect 11432 -4620 11442 -4560
rect 11502 -4610 11762 -4560
rect 11502 -4620 11512 -4610
rect 11432 -4630 11512 -4620
rect 11752 -4620 11762 -4610
rect 11822 -4620 11832 -4560
rect 11752 -4630 11832 -4620
rect 11432 -4900 11492 -4630
rect 11762 -4640 11832 -4630
rect 11572 -4690 11602 -4670
rect 11552 -4730 11602 -4690
rect 11662 -4690 11692 -4670
rect 11662 -4730 11712 -4690
rect 11552 -4800 11712 -4730
rect 11552 -4840 11602 -4800
rect 11572 -4860 11602 -4840
rect 11662 -4840 11712 -4800
rect 11662 -4860 11692 -4840
rect 11772 -4900 11832 -4640
rect 11432 -4910 11512 -4900
rect 11432 -4970 11442 -4910
rect 11502 -4920 11512 -4910
rect 11752 -4910 11832 -4900
rect 11752 -4920 11762 -4910
rect 11502 -4970 11762 -4920
rect 11822 -4970 11832 -4910
rect 11432 -4980 11832 -4970
rect 11890 -4560 12290 -4550
rect 11890 -4620 11900 -4560
rect 11960 -4610 12220 -4560
rect 11960 -4620 11970 -4610
rect 11890 -4630 11970 -4620
rect 12210 -4620 12220 -4610
rect 12280 -4620 12290 -4560
rect 12210 -4630 12290 -4620
rect 11890 -4900 11950 -4630
rect 12220 -4640 12290 -4630
rect 12030 -4690 12060 -4670
rect 12010 -4730 12060 -4690
rect 12120 -4690 12150 -4670
rect 12120 -4730 12170 -4690
rect 12010 -4800 12170 -4730
rect 12010 -4840 12060 -4800
rect 12030 -4860 12060 -4840
rect 12120 -4840 12170 -4800
rect 12120 -4860 12150 -4840
rect 12230 -4900 12290 -4640
rect 11890 -4910 11970 -4900
rect 11890 -4970 11900 -4910
rect 11960 -4920 11970 -4910
rect 12210 -4910 12290 -4900
rect 12210 -4920 12220 -4910
rect 11960 -4970 12220 -4920
rect 12280 -4970 12290 -4910
rect 11890 -4980 12290 -4970
rect 12346 -4560 12746 -4550
rect 12346 -4620 12356 -4560
rect 12416 -4610 12676 -4560
rect 12416 -4620 12426 -4610
rect 12346 -4630 12426 -4620
rect 12666 -4620 12676 -4610
rect 12736 -4620 12746 -4560
rect 12666 -4630 12746 -4620
rect 12346 -4900 12406 -4630
rect 12676 -4640 12746 -4630
rect 12486 -4690 12516 -4670
rect 12466 -4730 12516 -4690
rect 12576 -4690 12606 -4670
rect 12576 -4730 12626 -4690
rect 12466 -4800 12626 -4730
rect 12466 -4840 12516 -4800
rect 12486 -4860 12516 -4840
rect 12576 -4840 12626 -4800
rect 12576 -4860 12606 -4840
rect 12686 -4900 12746 -4640
rect 12346 -4910 12426 -4900
rect 12346 -4970 12356 -4910
rect 12416 -4920 12426 -4910
rect 12666 -4910 12746 -4900
rect 12666 -4920 12676 -4910
rect 12416 -4970 12676 -4920
rect 12736 -4970 12746 -4910
rect 12346 -4980 12746 -4970
rect 12802 -4560 13202 -4550
rect 12802 -4620 12812 -4560
rect 12872 -4610 13132 -4560
rect 12872 -4620 12882 -4610
rect 12802 -4630 12882 -4620
rect 13122 -4620 13132 -4610
rect 13192 -4620 13202 -4560
rect 13122 -4630 13202 -4620
rect 12802 -4900 12862 -4630
rect 13132 -4640 13202 -4630
rect 12942 -4690 12972 -4670
rect 12922 -4730 12972 -4690
rect 13032 -4690 13062 -4670
rect 13032 -4730 13082 -4690
rect 12922 -4800 13082 -4730
rect 12922 -4840 12972 -4800
rect 12942 -4860 12972 -4840
rect 13032 -4840 13082 -4800
rect 13032 -4860 13062 -4840
rect 13142 -4900 13202 -4640
rect 12802 -4910 12882 -4900
rect 12802 -4970 12812 -4910
rect 12872 -4920 12882 -4910
rect 13122 -4910 13202 -4900
rect 13122 -4920 13132 -4910
rect 12872 -4970 13132 -4920
rect 13192 -4970 13202 -4910
rect 12802 -4980 13202 -4970
rect 13260 -4560 13660 -4550
rect 13260 -4620 13270 -4560
rect 13330 -4610 13590 -4560
rect 13330 -4620 13340 -4610
rect 13260 -4630 13340 -4620
rect 13580 -4620 13590 -4610
rect 13650 -4620 13660 -4560
rect 13580 -4630 13660 -4620
rect 13260 -4900 13320 -4630
rect 13590 -4640 13660 -4630
rect 13400 -4690 13430 -4670
rect 13380 -4730 13430 -4690
rect 13490 -4690 13520 -4670
rect 13490 -4730 13540 -4690
rect 13380 -4800 13540 -4730
rect 13380 -4840 13430 -4800
rect 13400 -4860 13430 -4840
rect 13490 -4840 13540 -4800
rect 13490 -4860 13520 -4840
rect 13600 -4900 13660 -4640
rect 13260 -4910 13340 -4900
rect 13260 -4970 13270 -4910
rect 13330 -4920 13340 -4910
rect 13580 -4910 13660 -4900
rect 13580 -4920 13590 -4910
rect 13330 -4970 13590 -4920
rect 13650 -4970 13660 -4910
rect 13260 -4980 13660 -4970
rect 13716 -4560 14116 -4550
rect 13716 -4620 13726 -4560
rect 13786 -4610 14046 -4560
rect 13786 -4620 13796 -4610
rect 13716 -4630 13796 -4620
rect 14036 -4620 14046 -4610
rect 14106 -4620 14116 -4560
rect 14036 -4630 14116 -4620
rect 13716 -4900 13776 -4630
rect 14046 -4640 14116 -4630
rect 13856 -4690 13886 -4670
rect 13836 -4730 13886 -4690
rect 13946 -4690 13976 -4670
rect 13946 -4730 13996 -4690
rect 13836 -4800 13996 -4730
rect 13836 -4840 13886 -4800
rect 13856 -4860 13886 -4840
rect 13946 -4840 13996 -4800
rect 13946 -4860 13976 -4840
rect 14056 -4900 14116 -4640
rect 13716 -4910 13796 -4900
rect 13716 -4970 13726 -4910
rect 13786 -4920 13796 -4910
rect 14036 -4910 14116 -4900
rect 14036 -4920 14046 -4910
rect 13786 -4970 14046 -4920
rect 14106 -4970 14116 -4910
rect 13716 -4980 14116 -4970
rect 14172 -4560 14572 -4550
rect 14172 -4620 14182 -4560
rect 14242 -4610 14502 -4560
rect 14242 -4620 14252 -4610
rect 14172 -4630 14252 -4620
rect 14492 -4620 14502 -4610
rect 14562 -4620 14572 -4560
rect 14492 -4630 14572 -4620
rect 14172 -4900 14232 -4630
rect 14502 -4640 14572 -4630
rect 14312 -4690 14342 -4670
rect 14292 -4730 14342 -4690
rect 14402 -4690 14432 -4670
rect 14402 -4730 14452 -4690
rect 14292 -4800 14452 -4730
rect 14292 -4840 14342 -4800
rect 14312 -4860 14342 -4840
rect 14402 -4840 14452 -4800
rect 14402 -4860 14432 -4840
rect 14512 -4900 14572 -4640
rect 14172 -4910 14252 -4900
rect 14172 -4970 14182 -4910
rect 14242 -4920 14252 -4910
rect 14492 -4910 14572 -4900
rect 14492 -4920 14502 -4910
rect 14242 -4970 14502 -4920
rect 14562 -4970 14572 -4910
rect 14172 -4980 14572 -4970
rect 14630 -4560 15030 -4550
rect 14630 -4620 14640 -4560
rect 14700 -4610 14960 -4560
rect 14700 -4620 14710 -4610
rect 14630 -4630 14710 -4620
rect 14950 -4620 14960 -4610
rect 15020 -4620 15030 -4560
rect 14950 -4630 15030 -4620
rect 14630 -4900 14690 -4630
rect 14960 -4640 15030 -4630
rect 14770 -4690 14800 -4670
rect 14750 -4730 14800 -4690
rect 14860 -4690 14890 -4670
rect 14860 -4730 14910 -4690
rect 14750 -4800 14910 -4730
rect 14750 -4840 14800 -4800
rect 14770 -4860 14800 -4840
rect 14860 -4840 14910 -4800
rect 14860 -4860 14890 -4840
rect 14970 -4900 15030 -4640
rect 14630 -4910 14710 -4900
rect 14630 -4970 14640 -4910
rect 14700 -4920 14710 -4910
rect 14950 -4910 15030 -4900
rect 14950 -4920 14960 -4910
rect 14700 -4970 14960 -4920
rect 15020 -4970 15030 -4910
rect 14630 -4980 15030 -4970
rect 15086 -4560 15486 -4550
rect 15086 -4620 15096 -4560
rect 15156 -4610 15416 -4560
rect 15156 -4620 15166 -4610
rect 15086 -4630 15166 -4620
rect 15406 -4620 15416 -4610
rect 15476 -4620 15486 -4560
rect 15406 -4630 15486 -4620
rect 15086 -4900 15146 -4630
rect 15416 -4640 15486 -4630
rect 15226 -4690 15256 -4670
rect 15206 -4730 15256 -4690
rect 15316 -4690 15346 -4670
rect 15316 -4730 15366 -4690
rect 15206 -4800 15366 -4730
rect 15206 -4840 15256 -4800
rect 15226 -4860 15256 -4840
rect 15316 -4840 15366 -4800
rect 15316 -4860 15346 -4840
rect 15426 -4900 15486 -4640
rect 15086 -4910 15166 -4900
rect 15086 -4970 15096 -4910
rect 15156 -4920 15166 -4910
rect 15406 -4910 15486 -4900
rect 15406 -4920 15416 -4910
rect 15156 -4970 15416 -4920
rect 15476 -4970 15486 -4910
rect 15086 -4980 15486 -4970
rect 0 -5062 400 -5052
rect 0 -5122 10 -5062
rect 70 -5112 330 -5062
rect 70 -5122 80 -5112
rect 0 -5132 80 -5122
rect 320 -5122 330 -5112
rect 390 -5122 400 -5062
rect 320 -5132 400 -5122
rect 0 -5402 60 -5132
rect 330 -5142 400 -5132
rect 140 -5192 170 -5172
rect 120 -5232 170 -5192
rect 230 -5192 260 -5172
rect 230 -5232 280 -5192
rect 120 -5302 280 -5232
rect 120 -5342 170 -5302
rect 140 -5362 170 -5342
rect 230 -5342 280 -5302
rect 230 -5362 260 -5342
rect 340 -5402 400 -5142
rect 0 -5412 80 -5402
rect 0 -5472 10 -5412
rect 70 -5422 80 -5412
rect 320 -5412 400 -5402
rect 320 -5422 330 -5412
rect 70 -5472 330 -5422
rect 390 -5472 400 -5412
rect 0 -5482 400 -5472
rect 456 -5062 856 -5052
rect 456 -5122 466 -5062
rect 526 -5112 786 -5062
rect 526 -5122 536 -5112
rect 456 -5132 536 -5122
rect 776 -5122 786 -5112
rect 846 -5122 856 -5062
rect 776 -5132 856 -5122
rect 456 -5402 516 -5132
rect 786 -5142 856 -5132
rect 596 -5192 626 -5172
rect 576 -5232 626 -5192
rect 686 -5192 716 -5172
rect 686 -5232 736 -5192
rect 576 -5302 736 -5232
rect 576 -5342 626 -5302
rect 596 -5362 626 -5342
rect 686 -5342 736 -5302
rect 686 -5362 716 -5342
rect 796 -5402 856 -5142
rect 456 -5412 536 -5402
rect 456 -5472 466 -5412
rect 526 -5422 536 -5412
rect 776 -5412 856 -5402
rect 776 -5422 786 -5412
rect 526 -5472 786 -5422
rect 846 -5472 856 -5412
rect 456 -5482 856 -5472
rect 912 -5062 1312 -5052
rect 912 -5122 922 -5062
rect 982 -5112 1242 -5062
rect 982 -5122 992 -5112
rect 912 -5132 992 -5122
rect 1232 -5122 1242 -5112
rect 1302 -5122 1312 -5062
rect 1232 -5132 1312 -5122
rect 912 -5402 972 -5132
rect 1242 -5142 1312 -5132
rect 1052 -5192 1082 -5172
rect 1032 -5232 1082 -5192
rect 1142 -5192 1172 -5172
rect 1142 -5232 1192 -5192
rect 1032 -5302 1192 -5232
rect 1032 -5342 1082 -5302
rect 1052 -5362 1082 -5342
rect 1142 -5342 1192 -5302
rect 1142 -5362 1172 -5342
rect 1252 -5402 1312 -5142
rect 912 -5412 992 -5402
rect 912 -5472 922 -5412
rect 982 -5422 992 -5412
rect 1232 -5412 1312 -5402
rect 1232 -5422 1242 -5412
rect 982 -5472 1242 -5422
rect 1302 -5472 1312 -5412
rect 912 -5482 1312 -5472
rect 1370 -5062 1770 -5052
rect 1370 -5122 1380 -5062
rect 1440 -5112 1700 -5062
rect 1440 -5122 1450 -5112
rect 1370 -5132 1450 -5122
rect 1690 -5122 1700 -5112
rect 1760 -5122 1770 -5062
rect 1690 -5132 1770 -5122
rect 1370 -5402 1430 -5132
rect 1700 -5142 1770 -5132
rect 1510 -5192 1540 -5172
rect 1490 -5232 1540 -5192
rect 1600 -5192 1630 -5172
rect 1600 -5232 1650 -5192
rect 1490 -5302 1650 -5232
rect 1490 -5342 1540 -5302
rect 1510 -5362 1540 -5342
rect 1600 -5342 1650 -5302
rect 1600 -5362 1630 -5342
rect 1710 -5402 1770 -5142
rect 1370 -5412 1450 -5402
rect 1370 -5472 1380 -5412
rect 1440 -5422 1450 -5412
rect 1690 -5412 1770 -5402
rect 1690 -5422 1700 -5412
rect 1440 -5472 1700 -5422
rect 1760 -5472 1770 -5412
rect 1370 -5482 1770 -5472
rect 1826 -5062 2226 -5052
rect 1826 -5122 1836 -5062
rect 1896 -5112 2156 -5062
rect 1896 -5122 1906 -5112
rect 1826 -5132 1906 -5122
rect 2146 -5122 2156 -5112
rect 2216 -5122 2226 -5062
rect 2146 -5132 2226 -5122
rect 1826 -5402 1886 -5132
rect 2156 -5142 2226 -5132
rect 1966 -5192 1996 -5172
rect 1946 -5232 1996 -5192
rect 2056 -5192 2086 -5172
rect 2056 -5232 2106 -5192
rect 1946 -5302 2106 -5232
rect 1946 -5342 1996 -5302
rect 1966 -5362 1996 -5342
rect 2056 -5342 2106 -5302
rect 2056 -5362 2086 -5342
rect 2166 -5402 2226 -5142
rect 1826 -5412 1906 -5402
rect 1826 -5472 1836 -5412
rect 1896 -5422 1906 -5412
rect 2146 -5412 2226 -5402
rect 2146 -5422 2156 -5412
rect 1896 -5472 2156 -5422
rect 2216 -5472 2226 -5412
rect 1826 -5482 2226 -5472
rect 2282 -5062 2682 -5052
rect 2282 -5122 2292 -5062
rect 2352 -5112 2612 -5062
rect 2352 -5122 2362 -5112
rect 2282 -5132 2362 -5122
rect 2602 -5122 2612 -5112
rect 2672 -5122 2682 -5062
rect 2602 -5132 2682 -5122
rect 2282 -5402 2342 -5132
rect 2612 -5142 2682 -5132
rect 2422 -5192 2452 -5172
rect 2402 -5232 2452 -5192
rect 2512 -5192 2542 -5172
rect 2512 -5232 2562 -5192
rect 2402 -5302 2562 -5232
rect 2402 -5342 2452 -5302
rect 2422 -5362 2452 -5342
rect 2512 -5342 2562 -5302
rect 2512 -5362 2542 -5342
rect 2622 -5402 2682 -5142
rect 2282 -5412 2362 -5402
rect 2282 -5472 2292 -5412
rect 2352 -5422 2362 -5412
rect 2602 -5412 2682 -5402
rect 2602 -5422 2612 -5412
rect 2352 -5472 2612 -5422
rect 2672 -5472 2682 -5412
rect 2282 -5482 2682 -5472
rect 2740 -5062 3140 -5052
rect 2740 -5122 2750 -5062
rect 2810 -5112 3070 -5062
rect 2810 -5122 2820 -5112
rect 2740 -5132 2820 -5122
rect 3060 -5122 3070 -5112
rect 3130 -5122 3140 -5062
rect 3060 -5132 3140 -5122
rect 2740 -5402 2800 -5132
rect 3070 -5142 3140 -5132
rect 2880 -5192 2910 -5172
rect 2860 -5232 2910 -5192
rect 2970 -5192 3000 -5172
rect 2970 -5232 3020 -5192
rect 2860 -5302 3020 -5232
rect 2860 -5342 2910 -5302
rect 2880 -5362 2910 -5342
rect 2970 -5342 3020 -5302
rect 2970 -5362 3000 -5342
rect 3080 -5402 3140 -5142
rect 2740 -5412 2820 -5402
rect 2740 -5472 2750 -5412
rect 2810 -5422 2820 -5412
rect 3060 -5412 3140 -5402
rect 3060 -5422 3070 -5412
rect 2810 -5472 3070 -5422
rect 3130 -5472 3140 -5412
rect 2740 -5482 3140 -5472
rect 3196 -5062 3596 -5052
rect 3196 -5122 3206 -5062
rect 3266 -5112 3526 -5062
rect 3266 -5122 3276 -5112
rect 3196 -5132 3276 -5122
rect 3516 -5122 3526 -5112
rect 3586 -5122 3596 -5062
rect 3516 -5132 3596 -5122
rect 3196 -5402 3256 -5132
rect 3526 -5142 3596 -5132
rect 3336 -5192 3366 -5172
rect 3316 -5232 3366 -5192
rect 3426 -5192 3456 -5172
rect 3426 -5232 3476 -5192
rect 3316 -5302 3476 -5232
rect 3316 -5342 3366 -5302
rect 3336 -5362 3366 -5342
rect 3426 -5342 3476 -5302
rect 3426 -5362 3456 -5342
rect 3536 -5402 3596 -5142
rect 3196 -5412 3276 -5402
rect 3196 -5472 3206 -5412
rect 3266 -5422 3276 -5412
rect 3516 -5412 3596 -5402
rect 3516 -5422 3526 -5412
rect 3266 -5472 3526 -5422
rect 3586 -5472 3596 -5412
rect 3196 -5482 3596 -5472
rect 3652 -5062 4052 -5052
rect 3652 -5122 3662 -5062
rect 3722 -5112 3982 -5062
rect 3722 -5122 3732 -5112
rect 3652 -5132 3732 -5122
rect 3972 -5122 3982 -5112
rect 4042 -5122 4052 -5062
rect 3972 -5132 4052 -5122
rect 3652 -5402 3712 -5132
rect 3982 -5142 4052 -5132
rect 3792 -5192 3822 -5172
rect 3772 -5232 3822 -5192
rect 3882 -5192 3912 -5172
rect 3882 -5232 3932 -5192
rect 3772 -5302 3932 -5232
rect 3772 -5342 3822 -5302
rect 3792 -5362 3822 -5342
rect 3882 -5342 3932 -5302
rect 3882 -5362 3912 -5342
rect 3992 -5402 4052 -5142
rect 3652 -5412 3732 -5402
rect 3652 -5472 3662 -5412
rect 3722 -5422 3732 -5412
rect 3972 -5412 4052 -5402
rect 3972 -5422 3982 -5412
rect 3722 -5472 3982 -5422
rect 4042 -5472 4052 -5412
rect 3652 -5482 4052 -5472
rect 4110 -5062 4510 -5052
rect 4110 -5122 4120 -5062
rect 4180 -5112 4440 -5062
rect 4180 -5122 4190 -5112
rect 4110 -5132 4190 -5122
rect 4430 -5122 4440 -5112
rect 4500 -5122 4510 -5062
rect 4430 -5132 4510 -5122
rect 4110 -5402 4170 -5132
rect 4440 -5142 4510 -5132
rect 4250 -5192 4280 -5172
rect 4230 -5232 4280 -5192
rect 4340 -5192 4370 -5172
rect 4340 -5232 4390 -5192
rect 4230 -5302 4390 -5232
rect 4230 -5342 4280 -5302
rect 4250 -5362 4280 -5342
rect 4340 -5342 4390 -5302
rect 4340 -5362 4370 -5342
rect 4450 -5402 4510 -5142
rect 4110 -5412 4190 -5402
rect 4110 -5472 4120 -5412
rect 4180 -5422 4190 -5412
rect 4430 -5412 4510 -5402
rect 4430 -5422 4440 -5412
rect 4180 -5472 4440 -5422
rect 4500 -5472 4510 -5412
rect 4110 -5482 4510 -5472
rect 4566 -5062 4966 -5052
rect 4566 -5122 4576 -5062
rect 4636 -5112 4896 -5062
rect 4636 -5122 4646 -5112
rect 4566 -5132 4646 -5122
rect 4886 -5122 4896 -5112
rect 4956 -5122 4966 -5062
rect 4886 -5132 4966 -5122
rect 4566 -5402 4626 -5132
rect 4896 -5142 4966 -5132
rect 4706 -5192 4736 -5172
rect 4686 -5232 4736 -5192
rect 4796 -5192 4826 -5172
rect 4796 -5232 4846 -5192
rect 4686 -5302 4846 -5232
rect 4686 -5342 4736 -5302
rect 4706 -5362 4736 -5342
rect 4796 -5342 4846 -5302
rect 4796 -5362 4826 -5342
rect 4906 -5402 4966 -5142
rect 4566 -5412 4646 -5402
rect 4566 -5472 4576 -5412
rect 4636 -5422 4646 -5412
rect 4886 -5412 4966 -5402
rect 4886 -5422 4896 -5412
rect 4636 -5472 4896 -5422
rect 4956 -5472 4966 -5412
rect 4566 -5482 4966 -5472
rect 5022 -5062 5422 -5052
rect 5022 -5122 5032 -5062
rect 5092 -5112 5352 -5062
rect 5092 -5122 5102 -5112
rect 5022 -5132 5102 -5122
rect 5342 -5122 5352 -5112
rect 5412 -5122 5422 -5062
rect 5342 -5132 5422 -5122
rect 5022 -5402 5082 -5132
rect 5352 -5142 5422 -5132
rect 5162 -5192 5192 -5172
rect 5142 -5232 5192 -5192
rect 5252 -5192 5282 -5172
rect 5252 -5232 5302 -5192
rect 5142 -5302 5302 -5232
rect 5142 -5342 5192 -5302
rect 5162 -5362 5192 -5342
rect 5252 -5342 5302 -5302
rect 5252 -5362 5282 -5342
rect 5362 -5402 5422 -5142
rect 5022 -5412 5102 -5402
rect 5022 -5472 5032 -5412
rect 5092 -5422 5102 -5412
rect 5342 -5412 5422 -5402
rect 5342 -5422 5352 -5412
rect 5092 -5472 5352 -5422
rect 5412 -5472 5422 -5412
rect 5022 -5482 5422 -5472
rect 5480 -5062 5880 -5052
rect 5480 -5122 5490 -5062
rect 5550 -5112 5810 -5062
rect 5550 -5122 5560 -5112
rect 5480 -5132 5560 -5122
rect 5800 -5122 5810 -5112
rect 5870 -5122 5880 -5062
rect 5800 -5132 5880 -5122
rect 5480 -5402 5540 -5132
rect 5810 -5142 5880 -5132
rect 5620 -5192 5650 -5172
rect 5600 -5232 5650 -5192
rect 5710 -5192 5740 -5172
rect 5710 -5232 5760 -5192
rect 5600 -5302 5760 -5232
rect 5600 -5342 5650 -5302
rect 5620 -5362 5650 -5342
rect 5710 -5342 5760 -5302
rect 5710 -5362 5740 -5342
rect 5820 -5402 5880 -5142
rect 5480 -5412 5560 -5402
rect 5480 -5472 5490 -5412
rect 5550 -5422 5560 -5412
rect 5800 -5412 5880 -5402
rect 5800 -5422 5810 -5412
rect 5550 -5472 5810 -5422
rect 5870 -5472 5880 -5412
rect 5480 -5482 5880 -5472
rect 5936 -5062 6336 -5052
rect 5936 -5122 5946 -5062
rect 6006 -5112 6266 -5062
rect 6006 -5122 6016 -5112
rect 5936 -5132 6016 -5122
rect 6256 -5122 6266 -5112
rect 6326 -5122 6336 -5062
rect 6256 -5132 6336 -5122
rect 5936 -5402 5996 -5132
rect 6266 -5142 6336 -5132
rect 6076 -5192 6106 -5172
rect 6056 -5232 6106 -5192
rect 6166 -5192 6196 -5172
rect 6166 -5232 6216 -5192
rect 6056 -5302 6216 -5232
rect 6056 -5342 6106 -5302
rect 6076 -5362 6106 -5342
rect 6166 -5342 6216 -5302
rect 6166 -5362 6196 -5342
rect 6276 -5402 6336 -5142
rect 5936 -5412 6016 -5402
rect 5936 -5472 5946 -5412
rect 6006 -5422 6016 -5412
rect 6256 -5412 6336 -5402
rect 6256 -5422 6266 -5412
rect 6006 -5472 6266 -5422
rect 6326 -5472 6336 -5412
rect 5936 -5482 6336 -5472
rect 6392 -5062 6792 -5052
rect 6392 -5122 6402 -5062
rect 6462 -5112 6722 -5062
rect 6462 -5122 6472 -5112
rect 6392 -5132 6472 -5122
rect 6712 -5122 6722 -5112
rect 6782 -5122 6792 -5062
rect 6712 -5132 6792 -5122
rect 6392 -5402 6452 -5132
rect 6722 -5142 6792 -5132
rect 6532 -5192 6562 -5172
rect 6512 -5232 6562 -5192
rect 6622 -5192 6652 -5172
rect 6622 -5232 6672 -5192
rect 6512 -5302 6672 -5232
rect 6512 -5342 6562 -5302
rect 6532 -5362 6562 -5342
rect 6622 -5342 6672 -5302
rect 6622 -5362 6652 -5342
rect 6732 -5402 6792 -5142
rect 6392 -5412 6472 -5402
rect 6392 -5472 6402 -5412
rect 6462 -5422 6472 -5412
rect 6712 -5412 6792 -5402
rect 6712 -5422 6722 -5412
rect 6462 -5472 6722 -5422
rect 6782 -5472 6792 -5412
rect 6392 -5482 6792 -5472
rect 6850 -5062 7250 -5052
rect 6850 -5122 6860 -5062
rect 6920 -5112 7180 -5062
rect 6920 -5122 6930 -5112
rect 6850 -5132 6930 -5122
rect 7170 -5122 7180 -5112
rect 7240 -5122 7250 -5062
rect 7170 -5132 7250 -5122
rect 6850 -5402 6910 -5132
rect 7180 -5142 7250 -5132
rect 6990 -5192 7020 -5172
rect 6970 -5232 7020 -5192
rect 7080 -5192 7110 -5172
rect 7080 -5232 7130 -5192
rect 6970 -5302 7130 -5232
rect 6970 -5342 7020 -5302
rect 6990 -5362 7020 -5342
rect 7080 -5342 7130 -5302
rect 7080 -5362 7110 -5342
rect 7190 -5402 7250 -5142
rect 6850 -5412 6930 -5402
rect 6850 -5472 6860 -5412
rect 6920 -5422 6930 -5412
rect 7170 -5412 7250 -5402
rect 7170 -5422 7180 -5412
rect 6920 -5472 7180 -5422
rect 7240 -5472 7250 -5412
rect 6850 -5482 7250 -5472
rect 7306 -5062 7706 -5052
rect 7306 -5122 7316 -5062
rect 7376 -5112 7636 -5062
rect 7376 -5122 7386 -5112
rect 7306 -5132 7386 -5122
rect 7626 -5122 7636 -5112
rect 7696 -5122 7706 -5062
rect 7626 -5132 7706 -5122
rect 7306 -5402 7366 -5132
rect 7636 -5142 7706 -5132
rect 7446 -5192 7476 -5172
rect 7426 -5232 7476 -5192
rect 7536 -5192 7566 -5172
rect 7536 -5232 7586 -5192
rect 7426 -5302 7586 -5232
rect 7426 -5342 7476 -5302
rect 7446 -5362 7476 -5342
rect 7536 -5342 7586 -5302
rect 7536 -5362 7566 -5342
rect 7646 -5402 7706 -5142
rect 7306 -5412 7386 -5402
rect 7306 -5472 7316 -5412
rect 7376 -5422 7386 -5412
rect 7626 -5412 7706 -5402
rect 7626 -5422 7636 -5412
rect 7376 -5472 7636 -5422
rect 7696 -5472 7706 -5412
rect 7306 -5482 7706 -5472
rect 7762 -5062 8162 -5052
rect 7762 -5122 7772 -5062
rect 7832 -5112 8092 -5062
rect 7832 -5122 7842 -5112
rect 7762 -5132 7842 -5122
rect 8082 -5122 8092 -5112
rect 8152 -5122 8162 -5062
rect 8082 -5132 8162 -5122
rect 7762 -5402 7822 -5132
rect 8092 -5142 8162 -5132
rect 7902 -5192 7932 -5172
rect 7882 -5232 7932 -5192
rect 7992 -5192 8022 -5172
rect 7992 -5232 8042 -5192
rect 7882 -5302 8042 -5232
rect 7882 -5342 7932 -5302
rect 7902 -5362 7932 -5342
rect 7992 -5342 8042 -5302
rect 7992 -5362 8022 -5342
rect 8102 -5402 8162 -5142
rect 7762 -5412 7842 -5402
rect 7762 -5472 7772 -5412
rect 7832 -5422 7842 -5412
rect 8082 -5412 8162 -5402
rect 8082 -5422 8092 -5412
rect 7832 -5472 8092 -5422
rect 8152 -5472 8162 -5412
rect 7762 -5482 8162 -5472
rect 8236 -5062 8636 -5052
rect 8236 -5122 8246 -5062
rect 8306 -5112 8566 -5062
rect 8306 -5122 8316 -5112
rect 8236 -5132 8316 -5122
rect 8556 -5122 8566 -5112
rect 8626 -5122 8636 -5062
rect 8556 -5132 8636 -5122
rect 8236 -5402 8296 -5132
rect 8566 -5142 8636 -5132
rect 8376 -5192 8406 -5172
rect 8356 -5232 8406 -5192
rect 8466 -5192 8496 -5172
rect 8466 -5232 8516 -5192
rect 8356 -5302 8516 -5232
rect 8356 -5342 8406 -5302
rect 8376 -5362 8406 -5342
rect 8466 -5342 8516 -5302
rect 8466 -5362 8496 -5342
rect 8576 -5402 8636 -5142
rect 8236 -5412 8316 -5402
rect 8236 -5472 8246 -5412
rect 8306 -5422 8316 -5412
rect 8556 -5412 8636 -5402
rect 8556 -5422 8566 -5412
rect 8306 -5472 8566 -5422
rect 8626 -5472 8636 -5412
rect 8236 -5482 8636 -5472
rect 8692 -5062 9092 -5052
rect 8692 -5122 8702 -5062
rect 8762 -5112 9022 -5062
rect 8762 -5122 8772 -5112
rect 8692 -5132 8772 -5122
rect 9012 -5122 9022 -5112
rect 9082 -5122 9092 -5062
rect 9012 -5132 9092 -5122
rect 8692 -5402 8752 -5132
rect 9022 -5142 9092 -5132
rect 8832 -5192 8862 -5172
rect 8812 -5232 8862 -5192
rect 8922 -5192 8952 -5172
rect 8922 -5232 8972 -5192
rect 8812 -5302 8972 -5232
rect 8812 -5342 8862 -5302
rect 8832 -5362 8862 -5342
rect 8922 -5342 8972 -5302
rect 8922 -5362 8952 -5342
rect 9032 -5402 9092 -5142
rect 8692 -5412 8772 -5402
rect 8692 -5472 8702 -5412
rect 8762 -5422 8772 -5412
rect 9012 -5412 9092 -5402
rect 9012 -5422 9022 -5412
rect 8762 -5472 9022 -5422
rect 9082 -5472 9092 -5412
rect 8692 -5482 9092 -5472
rect 9150 -5062 9550 -5052
rect 9150 -5122 9160 -5062
rect 9220 -5112 9480 -5062
rect 9220 -5122 9230 -5112
rect 9150 -5132 9230 -5122
rect 9470 -5122 9480 -5112
rect 9540 -5122 9550 -5062
rect 9470 -5132 9550 -5122
rect 9150 -5402 9210 -5132
rect 9480 -5142 9550 -5132
rect 9290 -5192 9320 -5172
rect 9270 -5232 9320 -5192
rect 9380 -5192 9410 -5172
rect 9380 -5232 9430 -5192
rect 9270 -5302 9430 -5232
rect 9270 -5342 9320 -5302
rect 9290 -5362 9320 -5342
rect 9380 -5342 9430 -5302
rect 9380 -5362 9410 -5342
rect 9490 -5402 9550 -5142
rect 9150 -5412 9230 -5402
rect 9150 -5472 9160 -5412
rect 9220 -5422 9230 -5412
rect 9470 -5412 9550 -5402
rect 9470 -5422 9480 -5412
rect 9220 -5472 9480 -5422
rect 9540 -5472 9550 -5412
rect 9150 -5482 9550 -5472
rect 9606 -5062 10006 -5052
rect 9606 -5122 9616 -5062
rect 9676 -5112 9936 -5062
rect 9676 -5122 9686 -5112
rect 9606 -5132 9686 -5122
rect 9926 -5122 9936 -5112
rect 9996 -5122 10006 -5062
rect 9926 -5132 10006 -5122
rect 9606 -5402 9666 -5132
rect 9936 -5142 10006 -5132
rect 9746 -5192 9776 -5172
rect 9726 -5232 9776 -5192
rect 9836 -5192 9866 -5172
rect 9836 -5232 9886 -5192
rect 9726 -5302 9886 -5232
rect 9726 -5342 9776 -5302
rect 9746 -5362 9776 -5342
rect 9836 -5342 9886 -5302
rect 9836 -5362 9866 -5342
rect 9946 -5402 10006 -5142
rect 9606 -5412 9686 -5402
rect 9606 -5472 9616 -5412
rect 9676 -5422 9686 -5412
rect 9926 -5412 10006 -5402
rect 9926 -5422 9936 -5412
rect 9676 -5472 9936 -5422
rect 9996 -5472 10006 -5412
rect 9606 -5482 10006 -5472
rect 10062 -5062 10462 -5052
rect 10062 -5122 10072 -5062
rect 10132 -5112 10392 -5062
rect 10132 -5122 10142 -5112
rect 10062 -5132 10142 -5122
rect 10382 -5122 10392 -5112
rect 10452 -5122 10462 -5062
rect 10382 -5132 10462 -5122
rect 10062 -5402 10122 -5132
rect 10392 -5142 10462 -5132
rect 10202 -5192 10232 -5172
rect 10182 -5232 10232 -5192
rect 10292 -5192 10322 -5172
rect 10292 -5232 10342 -5192
rect 10182 -5302 10342 -5232
rect 10182 -5342 10232 -5302
rect 10202 -5362 10232 -5342
rect 10292 -5342 10342 -5302
rect 10292 -5362 10322 -5342
rect 10402 -5402 10462 -5142
rect 10062 -5412 10142 -5402
rect 10062 -5472 10072 -5412
rect 10132 -5422 10142 -5412
rect 10382 -5412 10462 -5402
rect 10382 -5422 10392 -5412
rect 10132 -5472 10392 -5422
rect 10452 -5472 10462 -5412
rect 10062 -5482 10462 -5472
rect 10520 -5062 10920 -5052
rect 10520 -5122 10530 -5062
rect 10590 -5112 10850 -5062
rect 10590 -5122 10600 -5112
rect 10520 -5132 10600 -5122
rect 10840 -5122 10850 -5112
rect 10910 -5122 10920 -5062
rect 10840 -5132 10920 -5122
rect 10520 -5402 10580 -5132
rect 10850 -5142 10920 -5132
rect 10660 -5192 10690 -5172
rect 10640 -5232 10690 -5192
rect 10750 -5192 10780 -5172
rect 10750 -5232 10800 -5192
rect 10640 -5302 10800 -5232
rect 10640 -5342 10690 -5302
rect 10660 -5362 10690 -5342
rect 10750 -5342 10800 -5302
rect 10750 -5362 10780 -5342
rect 10860 -5402 10920 -5142
rect 10520 -5412 10600 -5402
rect 10520 -5472 10530 -5412
rect 10590 -5422 10600 -5412
rect 10840 -5412 10920 -5402
rect 10840 -5422 10850 -5412
rect 10590 -5472 10850 -5422
rect 10910 -5472 10920 -5412
rect 10520 -5482 10920 -5472
rect 10976 -5062 11376 -5052
rect 10976 -5122 10986 -5062
rect 11046 -5112 11306 -5062
rect 11046 -5122 11056 -5112
rect 10976 -5132 11056 -5122
rect 11296 -5122 11306 -5112
rect 11366 -5122 11376 -5062
rect 11296 -5132 11376 -5122
rect 10976 -5402 11036 -5132
rect 11306 -5142 11376 -5132
rect 11116 -5192 11146 -5172
rect 11096 -5232 11146 -5192
rect 11206 -5192 11236 -5172
rect 11206 -5232 11256 -5192
rect 11096 -5302 11256 -5232
rect 11096 -5342 11146 -5302
rect 11116 -5362 11146 -5342
rect 11206 -5342 11256 -5302
rect 11206 -5362 11236 -5342
rect 11316 -5402 11376 -5142
rect 10976 -5412 11056 -5402
rect 10976 -5472 10986 -5412
rect 11046 -5422 11056 -5412
rect 11296 -5412 11376 -5402
rect 11296 -5422 11306 -5412
rect 11046 -5472 11306 -5422
rect 11366 -5472 11376 -5412
rect 10976 -5482 11376 -5472
rect 11432 -5062 11832 -5052
rect 11432 -5122 11442 -5062
rect 11502 -5112 11762 -5062
rect 11502 -5122 11512 -5112
rect 11432 -5132 11512 -5122
rect 11752 -5122 11762 -5112
rect 11822 -5122 11832 -5062
rect 11752 -5132 11832 -5122
rect 11432 -5402 11492 -5132
rect 11762 -5142 11832 -5132
rect 11572 -5192 11602 -5172
rect 11552 -5232 11602 -5192
rect 11662 -5192 11692 -5172
rect 11662 -5232 11712 -5192
rect 11552 -5302 11712 -5232
rect 11552 -5342 11602 -5302
rect 11572 -5362 11602 -5342
rect 11662 -5342 11712 -5302
rect 11662 -5362 11692 -5342
rect 11772 -5402 11832 -5142
rect 11432 -5412 11512 -5402
rect 11432 -5472 11442 -5412
rect 11502 -5422 11512 -5412
rect 11752 -5412 11832 -5402
rect 11752 -5422 11762 -5412
rect 11502 -5472 11762 -5422
rect 11822 -5472 11832 -5412
rect 11432 -5482 11832 -5472
rect 11890 -5062 12290 -5052
rect 11890 -5122 11900 -5062
rect 11960 -5112 12220 -5062
rect 11960 -5122 11970 -5112
rect 11890 -5132 11970 -5122
rect 12210 -5122 12220 -5112
rect 12280 -5122 12290 -5062
rect 12210 -5132 12290 -5122
rect 11890 -5402 11950 -5132
rect 12220 -5142 12290 -5132
rect 12030 -5192 12060 -5172
rect 12010 -5232 12060 -5192
rect 12120 -5192 12150 -5172
rect 12120 -5232 12170 -5192
rect 12010 -5302 12170 -5232
rect 12010 -5342 12060 -5302
rect 12030 -5362 12060 -5342
rect 12120 -5342 12170 -5302
rect 12120 -5362 12150 -5342
rect 12230 -5402 12290 -5142
rect 11890 -5412 11970 -5402
rect 11890 -5472 11900 -5412
rect 11960 -5422 11970 -5412
rect 12210 -5412 12290 -5402
rect 12210 -5422 12220 -5412
rect 11960 -5472 12220 -5422
rect 12280 -5472 12290 -5412
rect 11890 -5482 12290 -5472
rect 12346 -5062 12746 -5052
rect 12346 -5122 12356 -5062
rect 12416 -5112 12676 -5062
rect 12416 -5122 12426 -5112
rect 12346 -5132 12426 -5122
rect 12666 -5122 12676 -5112
rect 12736 -5122 12746 -5062
rect 12666 -5132 12746 -5122
rect 12346 -5402 12406 -5132
rect 12676 -5142 12746 -5132
rect 12486 -5192 12516 -5172
rect 12466 -5232 12516 -5192
rect 12576 -5192 12606 -5172
rect 12576 -5232 12626 -5192
rect 12466 -5302 12626 -5232
rect 12466 -5342 12516 -5302
rect 12486 -5362 12516 -5342
rect 12576 -5342 12626 -5302
rect 12576 -5362 12606 -5342
rect 12686 -5402 12746 -5142
rect 12346 -5412 12426 -5402
rect 12346 -5472 12356 -5412
rect 12416 -5422 12426 -5412
rect 12666 -5412 12746 -5402
rect 12666 -5422 12676 -5412
rect 12416 -5472 12676 -5422
rect 12736 -5472 12746 -5412
rect 12346 -5482 12746 -5472
rect 12802 -5062 13202 -5052
rect 12802 -5122 12812 -5062
rect 12872 -5112 13132 -5062
rect 12872 -5122 12882 -5112
rect 12802 -5132 12882 -5122
rect 13122 -5122 13132 -5112
rect 13192 -5122 13202 -5062
rect 13122 -5132 13202 -5122
rect 12802 -5402 12862 -5132
rect 13132 -5142 13202 -5132
rect 12942 -5192 12972 -5172
rect 12922 -5232 12972 -5192
rect 13032 -5192 13062 -5172
rect 13032 -5232 13082 -5192
rect 12922 -5302 13082 -5232
rect 12922 -5342 12972 -5302
rect 12942 -5362 12972 -5342
rect 13032 -5342 13082 -5302
rect 13032 -5362 13062 -5342
rect 13142 -5402 13202 -5142
rect 12802 -5412 12882 -5402
rect 12802 -5472 12812 -5412
rect 12872 -5422 12882 -5412
rect 13122 -5412 13202 -5402
rect 13122 -5422 13132 -5412
rect 12872 -5472 13132 -5422
rect 13192 -5472 13202 -5412
rect 12802 -5482 13202 -5472
rect 13260 -5062 13660 -5052
rect 13260 -5122 13270 -5062
rect 13330 -5112 13590 -5062
rect 13330 -5122 13340 -5112
rect 13260 -5132 13340 -5122
rect 13580 -5122 13590 -5112
rect 13650 -5122 13660 -5062
rect 13580 -5132 13660 -5122
rect 13260 -5402 13320 -5132
rect 13590 -5142 13660 -5132
rect 13400 -5192 13430 -5172
rect 13380 -5232 13430 -5192
rect 13490 -5192 13520 -5172
rect 13490 -5232 13540 -5192
rect 13380 -5302 13540 -5232
rect 13380 -5342 13430 -5302
rect 13400 -5362 13430 -5342
rect 13490 -5342 13540 -5302
rect 13490 -5362 13520 -5342
rect 13600 -5402 13660 -5142
rect 13260 -5412 13340 -5402
rect 13260 -5472 13270 -5412
rect 13330 -5422 13340 -5412
rect 13580 -5412 13660 -5402
rect 13580 -5422 13590 -5412
rect 13330 -5472 13590 -5422
rect 13650 -5472 13660 -5412
rect 13260 -5482 13660 -5472
rect 13716 -5062 14116 -5052
rect 13716 -5122 13726 -5062
rect 13786 -5112 14046 -5062
rect 13786 -5122 13796 -5112
rect 13716 -5132 13796 -5122
rect 14036 -5122 14046 -5112
rect 14106 -5122 14116 -5062
rect 14036 -5132 14116 -5122
rect 13716 -5402 13776 -5132
rect 14046 -5142 14116 -5132
rect 13856 -5192 13886 -5172
rect 13836 -5232 13886 -5192
rect 13946 -5192 13976 -5172
rect 13946 -5232 13996 -5192
rect 13836 -5302 13996 -5232
rect 13836 -5342 13886 -5302
rect 13856 -5362 13886 -5342
rect 13946 -5342 13996 -5302
rect 13946 -5362 13976 -5342
rect 14056 -5402 14116 -5142
rect 13716 -5412 13796 -5402
rect 13716 -5472 13726 -5412
rect 13786 -5422 13796 -5412
rect 14036 -5412 14116 -5402
rect 14036 -5422 14046 -5412
rect 13786 -5472 14046 -5422
rect 14106 -5472 14116 -5412
rect 13716 -5482 14116 -5472
rect 14172 -5062 14572 -5052
rect 14172 -5122 14182 -5062
rect 14242 -5112 14502 -5062
rect 14242 -5122 14252 -5112
rect 14172 -5132 14252 -5122
rect 14492 -5122 14502 -5112
rect 14562 -5122 14572 -5062
rect 14492 -5132 14572 -5122
rect 14172 -5402 14232 -5132
rect 14502 -5142 14572 -5132
rect 14312 -5192 14342 -5172
rect 14292 -5232 14342 -5192
rect 14402 -5192 14432 -5172
rect 14402 -5232 14452 -5192
rect 14292 -5302 14452 -5232
rect 14292 -5342 14342 -5302
rect 14312 -5362 14342 -5342
rect 14402 -5342 14452 -5302
rect 14402 -5362 14432 -5342
rect 14512 -5402 14572 -5142
rect 14172 -5412 14252 -5402
rect 14172 -5472 14182 -5412
rect 14242 -5422 14252 -5412
rect 14492 -5412 14572 -5402
rect 14492 -5422 14502 -5412
rect 14242 -5472 14502 -5422
rect 14562 -5472 14572 -5412
rect 14172 -5482 14572 -5472
rect 14630 -5062 15030 -5052
rect 14630 -5122 14640 -5062
rect 14700 -5112 14960 -5062
rect 14700 -5122 14710 -5112
rect 14630 -5132 14710 -5122
rect 14950 -5122 14960 -5112
rect 15020 -5122 15030 -5062
rect 14950 -5132 15030 -5122
rect 14630 -5402 14690 -5132
rect 14960 -5142 15030 -5132
rect 14770 -5192 14800 -5172
rect 14750 -5232 14800 -5192
rect 14860 -5192 14890 -5172
rect 14860 -5232 14910 -5192
rect 14750 -5302 14910 -5232
rect 14750 -5342 14800 -5302
rect 14770 -5362 14800 -5342
rect 14860 -5342 14910 -5302
rect 14860 -5362 14890 -5342
rect 14970 -5402 15030 -5142
rect 14630 -5412 14710 -5402
rect 14630 -5472 14640 -5412
rect 14700 -5422 14710 -5412
rect 14950 -5412 15030 -5402
rect 14950 -5422 14960 -5412
rect 14700 -5472 14960 -5422
rect 15020 -5472 15030 -5412
rect 14630 -5482 15030 -5472
rect 15086 -5062 15486 -5052
rect 15086 -5122 15096 -5062
rect 15156 -5112 15416 -5062
rect 15156 -5122 15166 -5112
rect 15086 -5132 15166 -5122
rect 15406 -5122 15416 -5112
rect 15476 -5122 15486 -5062
rect 15406 -5132 15486 -5122
rect 15086 -5402 15146 -5132
rect 15416 -5142 15486 -5132
rect 15226 -5192 15256 -5172
rect 15206 -5232 15256 -5192
rect 15316 -5192 15346 -5172
rect 15316 -5232 15366 -5192
rect 15206 -5302 15366 -5232
rect 15206 -5342 15256 -5302
rect 15226 -5362 15256 -5342
rect 15316 -5342 15366 -5302
rect 15316 -5362 15346 -5342
rect 15426 -5402 15486 -5142
rect 15086 -5412 15166 -5402
rect 15086 -5472 15096 -5412
rect 15156 -5422 15166 -5412
rect 15406 -5412 15486 -5402
rect 15406 -5422 15416 -5412
rect 15156 -5472 15416 -5422
rect 15476 -5472 15486 -5412
rect 15086 -5482 15486 -5472
rect 0 -5554 400 -5544
rect 0 -5614 10 -5554
rect 70 -5604 330 -5554
rect 70 -5614 80 -5604
rect 0 -5624 80 -5614
rect 320 -5614 330 -5604
rect 390 -5614 400 -5554
rect 320 -5624 400 -5614
rect 0 -5894 60 -5624
rect 330 -5634 400 -5624
rect 140 -5684 170 -5664
rect 120 -5724 170 -5684
rect 230 -5684 260 -5664
rect 230 -5724 280 -5684
rect 120 -5794 280 -5724
rect 120 -5834 170 -5794
rect 140 -5854 170 -5834
rect 230 -5834 280 -5794
rect 230 -5854 260 -5834
rect 340 -5894 400 -5634
rect 0 -5904 80 -5894
rect 0 -5964 10 -5904
rect 70 -5914 80 -5904
rect 320 -5904 400 -5894
rect 320 -5914 330 -5904
rect 70 -5964 330 -5914
rect 390 -5964 400 -5904
rect 0 -5974 400 -5964
rect 456 -5554 856 -5544
rect 456 -5614 466 -5554
rect 526 -5604 786 -5554
rect 526 -5614 536 -5604
rect 456 -5624 536 -5614
rect 776 -5614 786 -5604
rect 846 -5614 856 -5554
rect 776 -5624 856 -5614
rect 456 -5894 516 -5624
rect 786 -5634 856 -5624
rect 596 -5684 626 -5664
rect 576 -5724 626 -5684
rect 686 -5684 716 -5664
rect 686 -5724 736 -5684
rect 576 -5794 736 -5724
rect 576 -5834 626 -5794
rect 596 -5854 626 -5834
rect 686 -5834 736 -5794
rect 686 -5854 716 -5834
rect 796 -5894 856 -5634
rect 456 -5904 536 -5894
rect 456 -5964 466 -5904
rect 526 -5914 536 -5904
rect 776 -5904 856 -5894
rect 776 -5914 786 -5904
rect 526 -5964 786 -5914
rect 846 -5964 856 -5904
rect 456 -5974 856 -5964
rect 912 -5554 1312 -5544
rect 912 -5614 922 -5554
rect 982 -5604 1242 -5554
rect 982 -5614 992 -5604
rect 912 -5624 992 -5614
rect 1232 -5614 1242 -5604
rect 1302 -5614 1312 -5554
rect 1232 -5624 1312 -5614
rect 912 -5894 972 -5624
rect 1242 -5634 1312 -5624
rect 1052 -5684 1082 -5664
rect 1032 -5724 1082 -5684
rect 1142 -5684 1172 -5664
rect 1142 -5724 1192 -5684
rect 1032 -5794 1192 -5724
rect 1032 -5834 1082 -5794
rect 1052 -5854 1082 -5834
rect 1142 -5834 1192 -5794
rect 1142 -5854 1172 -5834
rect 1252 -5894 1312 -5634
rect 912 -5904 992 -5894
rect 912 -5964 922 -5904
rect 982 -5914 992 -5904
rect 1232 -5904 1312 -5894
rect 1232 -5914 1242 -5904
rect 982 -5964 1242 -5914
rect 1302 -5964 1312 -5904
rect 912 -5974 1312 -5964
rect 1370 -5554 1770 -5544
rect 1370 -5614 1380 -5554
rect 1440 -5604 1700 -5554
rect 1440 -5614 1450 -5604
rect 1370 -5624 1450 -5614
rect 1690 -5614 1700 -5604
rect 1760 -5614 1770 -5554
rect 1690 -5624 1770 -5614
rect 1370 -5894 1430 -5624
rect 1700 -5634 1770 -5624
rect 1510 -5684 1540 -5664
rect 1490 -5724 1540 -5684
rect 1600 -5684 1630 -5664
rect 1600 -5724 1650 -5684
rect 1490 -5794 1650 -5724
rect 1490 -5834 1540 -5794
rect 1510 -5854 1540 -5834
rect 1600 -5834 1650 -5794
rect 1600 -5854 1630 -5834
rect 1710 -5894 1770 -5634
rect 1370 -5904 1450 -5894
rect 1370 -5964 1380 -5904
rect 1440 -5914 1450 -5904
rect 1690 -5904 1770 -5894
rect 1690 -5914 1700 -5904
rect 1440 -5964 1700 -5914
rect 1760 -5964 1770 -5904
rect 1370 -5974 1770 -5964
rect 1826 -5554 2226 -5544
rect 1826 -5614 1836 -5554
rect 1896 -5604 2156 -5554
rect 1896 -5614 1906 -5604
rect 1826 -5624 1906 -5614
rect 2146 -5614 2156 -5604
rect 2216 -5614 2226 -5554
rect 2146 -5624 2226 -5614
rect 1826 -5894 1886 -5624
rect 2156 -5634 2226 -5624
rect 1966 -5684 1996 -5664
rect 1946 -5724 1996 -5684
rect 2056 -5684 2086 -5664
rect 2056 -5724 2106 -5684
rect 1946 -5794 2106 -5724
rect 1946 -5834 1996 -5794
rect 1966 -5854 1996 -5834
rect 2056 -5834 2106 -5794
rect 2056 -5854 2086 -5834
rect 2166 -5894 2226 -5634
rect 1826 -5904 1906 -5894
rect 1826 -5964 1836 -5904
rect 1896 -5914 1906 -5904
rect 2146 -5904 2226 -5894
rect 2146 -5914 2156 -5904
rect 1896 -5964 2156 -5914
rect 2216 -5964 2226 -5904
rect 1826 -5974 2226 -5964
rect 2282 -5554 2682 -5544
rect 2282 -5614 2292 -5554
rect 2352 -5604 2612 -5554
rect 2352 -5614 2362 -5604
rect 2282 -5624 2362 -5614
rect 2602 -5614 2612 -5604
rect 2672 -5614 2682 -5554
rect 2602 -5624 2682 -5614
rect 2282 -5894 2342 -5624
rect 2612 -5634 2682 -5624
rect 2422 -5684 2452 -5664
rect 2402 -5724 2452 -5684
rect 2512 -5684 2542 -5664
rect 2512 -5724 2562 -5684
rect 2402 -5794 2562 -5724
rect 2402 -5834 2452 -5794
rect 2422 -5854 2452 -5834
rect 2512 -5834 2562 -5794
rect 2512 -5854 2542 -5834
rect 2622 -5894 2682 -5634
rect 2282 -5904 2362 -5894
rect 2282 -5964 2292 -5904
rect 2352 -5914 2362 -5904
rect 2602 -5904 2682 -5894
rect 2602 -5914 2612 -5904
rect 2352 -5964 2612 -5914
rect 2672 -5964 2682 -5904
rect 2282 -5974 2682 -5964
rect 2740 -5554 3140 -5544
rect 2740 -5614 2750 -5554
rect 2810 -5604 3070 -5554
rect 2810 -5614 2820 -5604
rect 2740 -5624 2820 -5614
rect 3060 -5614 3070 -5604
rect 3130 -5614 3140 -5554
rect 3060 -5624 3140 -5614
rect 2740 -5894 2800 -5624
rect 3070 -5634 3140 -5624
rect 2880 -5684 2910 -5664
rect 2860 -5724 2910 -5684
rect 2970 -5684 3000 -5664
rect 2970 -5724 3020 -5684
rect 2860 -5794 3020 -5724
rect 2860 -5834 2910 -5794
rect 2880 -5854 2910 -5834
rect 2970 -5834 3020 -5794
rect 2970 -5854 3000 -5834
rect 3080 -5894 3140 -5634
rect 2740 -5904 2820 -5894
rect 2740 -5964 2750 -5904
rect 2810 -5914 2820 -5904
rect 3060 -5904 3140 -5894
rect 3060 -5914 3070 -5904
rect 2810 -5964 3070 -5914
rect 3130 -5964 3140 -5904
rect 2740 -5974 3140 -5964
rect 3196 -5554 3596 -5544
rect 3196 -5614 3206 -5554
rect 3266 -5604 3526 -5554
rect 3266 -5614 3276 -5604
rect 3196 -5624 3276 -5614
rect 3516 -5614 3526 -5604
rect 3586 -5614 3596 -5554
rect 3516 -5624 3596 -5614
rect 3196 -5894 3256 -5624
rect 3526 -5634 3596 -5624
rect 3336 -5684 3366 -5664
rect 3316 -5724 3366 -5684
rect 3426 -5684 3456 -5664
rect 3426 -5724 3476 -5684
rect 3316 -5794 3476 -5724
rect 3316 -5834 3366 -5794
rect 3336 -5854 3366 -5834
rect 3426 -5834 3476 -5794
rect 3426 -5854 3456 -5834
rect 3536 -5894 3596 -5634
rect 3196 -5904 3276 -5894
rect 3196 -5964 3206 -5904
rect 3266 -5914 3276 -5904
rect 3516 -5904 3596 -5894
rect 3516 -5914 3526 -5904
rect 3266 -5964 3526 -5914
rect 3586 -5964 3596 -5904
rect 3196 -5974 3596 -5964
rect 3652 -5554 4052 -5544
rect 3652 -5614 3662 -5554
rect 3722 -5604 3982 -5554
rect 3722 -5614 3732 -5604
rect 3652 -5624 3732 -5614
rect 3972 -5614 3982 -5604
rect 4042 -5614 4052 -5554
rect 3972 -5624 4052 -5614
rect 3652 -5894 3712 -5624
rect 3982 -5634 4052 -5624
rect 3792 -5684 3822 -5664
rect 3772 -5724 3822 -5684
rect 3882 -5684 3912 -5664
rect 3882 -5724 3932 -5684
rect 3772 -5794 3932 -5724
rect 3772 -5834 3822 -5794
rect 3792 -5854 3822 -5834
rect 3882 -5834 3932 -5794
rect 3882 -5854 3912 -5834
rect 3992 -5894 4052 -5634
rect 3652 -5904 3732 -5894
rect 3652 -5964 3662 -5904
rect 3722 -5914 3732 -5904
rect 3972 -5904 4052 -5894
rect 3972 -5914 3982 -5904
rect 3722 -5964 3982 -5914
rect 4042 -5964 4052 -5904
rect 3652 -5974 4052 -5964
rect 4110 -5554 4510 -5544
rect 4110 -5614 4120 -5554
rect 4180 -5604 4440 -5554
rect 4180 -5614 4190 -5604
rect 4110 -5624 4190 -5614
rect 4430 -5614 4440 -5604
rect 4500 -5614 4510 -5554
rect 4430 -5624 4510 -5614
rect 4110 -5894 4170 -5624
rect 4440 -5634 4510 -5624
rect 4250 -5684 4280 -5664
rect 4230 -5724 4280 -5684
rect 4340 -5684 4370 -5664
rect 4340 -5724 4390 -5684
rect 4230 -5794 4390 -5724
rect 4230 -5834 4280 -5794
rect 4250 -5854 4280 -5834
rect 4340 -5834 4390 -5794
rect 4340 -5854 4370 -5834
rect 4450 -5894 4510 -5634
rect 4110 -5904 4190 -5894
rect 4110 -5964 4120 -5904
rect 4180 -5914 4190 -5904
rect 4430 -5904 4510 -5894
rect 4430 -5914 4440 -5904
rect 4180 -5964 4440 -5914
rect 4500 -5964 4510 -5904
rect 4110 -5974 4510 -5964
rect 4566 -5554 4966 -5544
rect 4566 -5614 4576 -5554
rect 4636 -5604 4896 -5554
rect 4636 -5614 4646 -5604
rect 4566 -5624 4646 -5614
rect 4886 -5614 4896 -5604
rect 4956 -5614 4966 -5554
rect 4886 -5624 4966 -5614
rect 4566 -5894 4626 -5624
rect 4896 -5634 4966 -5624
rect 4706 -5684 4736 -5664
rect 4686 -5724 4736 -5684
rect 4796 -5684 4826 -5664
rect 4796 -5724 4846 -5684
rect 4686 -5794 4846 -5724
rect 4686 -5834 4736 -5794
rect 4706 -5854 4736 -5834
rect 4796 -5834 4846 -5794
rect 4796 -5854 4826 -5834
rect 4906 -5894 4966 -5634
rect 4566 -5904 4646 -5894
rect 4566 -5964 4576 -5904
rect 4636 -5914 4646 -5904
rect 4886 -5904 4966 -5894
rect 4886 -5914 4896 -5904
rect 4636 -5964 4896 -5914
rect 4956 -5964 4966 -5904
rect 4566 -5974 4966 -5964
rect 5022 -5554 5422 -5544
rect 5022 -5614 5032 -5554
rect 5092 -5604 5352 -5554
rect 5092 -5614 5102 -5604
rect 5022 -5624 5102 -5614
rect 5342 -5614 5352 -5604
rect 5412 -5614 5422 -5554
rect 5342 -5624 5422 -5614
rect 5022 -5894 5082 -5624
rect 5352 -5634 5422 -5624
rect 5162 -5684 5192 -5664
rect 5142 -5724 5192 -5684
rect 5252 -5684 5282 -5664
rect 5252 -5724 5302 -5684
rect 5142 -5794 5302 -5724
rect 5142 -5834 5192 -5794
rect 5162 -5854 5192 -5834
rect 5252 -5834 5302 -5794
rect 5252 -5854 5282 -5834
rect 5362 -5894 5422 -5634
rect 5022 -5904 5102 -5894
rect 5022 -5964 5032 -5904
rect 5092 -5914 5102 -5904
rect 5342 -5904 5422 -5894
rect 5342 -5914 5352 -5904
rect 5092 -5964 5352 -5914
rect 5412 -5964 5422 -5904
rect 5022 -5974 5422 -5964
rect 5480 -5554 5880 -5544
rect 5480 -5614 5490 -5554
rect 5550 -5604 5810 -5554
rect 5550 -5614 5560 -5604
rect 5480 -5624 5560 -5614
rect 5800 -5614 5810 -5604
rect 5870 -5614 5880 -5554
rect 5800 -5624 5880 -5614
rect 5480 -5894 5540 -5624
rect 5810 -5634 5880 -5624
rect 5620 -5684 5650 -5664
rect 5600 -5724 5650 -5684
rect 5710 -5684 5740 -5664
rect 5710 -5724 5760 -5684
rect 5600 -5794 5760 -5724
rect 5600 -5834 5650 -5794
rect 5620 -5854 5650 -5834
rect 5710 -5834 5760 -5794
rect 5710 -5854 5740 -5834
rect 5820 -5894 5880 -5634
rect 5480 -5904 5560 -5894
rect 5480 -5964 5490 -5904
rect 5550 -5914 5560 -5904
rect 5800 -5904 5880 -5894
rect 5800 -5914 5810 -5904
rect 5550 -5964 5810 -5914
rect 5870 -5964 5880 -5904
rect 5480 -5974 5880 -5964
rect 5936 -5554 6336 -5544
rect 5936 -5614 5946 -5554
rect 6006 -5604 6266 -5554
rect 6006 -5614 6016 -5604
rect 5936 -5624 6016 -5614
rect 6256 -5614 6266 -5604
rect 6326 -5614 6336 -5554
rect 6256 -5624 6336 -5614
rect 5936 -5894 5996 -5624
rect 6266 -5634 6336 -5624
rect 6076 -5684 6106 -5664
rect 6056 -5724 6106 -5684
rect 6166 -5684 6196 -5664
rect 6166 -5724 6216 -5684
rect 6056 -5794 6216 -5724
rect 6056 -5834 6106 -5794
rect 6076 -5854 6106 -5834
rect 6166 -5834 6216 -5794
rect 6166 -5854 6196 -5834
rect 6276 -5894 6336 -5634
rect 5936 -5904 6016 -5894
rect 5936 -5964 5946 -5904
rect 6006 -5914 6016 -5904
rect 6256 -5904 6336 -5894
rect 6256 -5914 6266 -5904
rect 6006 -5964 6266 -5914
rect 6326 -5964 6336 -5904
rect 5936 -5974 6336 -5964
rect 6392 -5554 6792 -5544
rect 6392 -5614 6402 -5554
rect 6462 -5604 6722 -5554
rect 6462 -5614 6472 -5604
rect 6392 -5624 6472 -5614
rect 6712 -5614 6722 -5604
rect 6782 -5614 6792 -5554
rect 6712 -5624 6792 -5614
rect 6392 -5894 6452 -5624
rect 6722 -5634 6792 -5624
rect 6532 -5684 6562 -5664
rect 6512 -5724 6562 -5684
rect 6622 -5684 6652 -5664
rect 6622 -5724 6672 -5684
rect 6512 -5794 6672 -5724
rect 6512 -5834 6562 -5794
rect 6532 -5854 6562 -5834
rect 6622 -5834 6672 -5794
rect 6622 -5854 6652 -5834
rect 6732 -5894 6792 -5634
rect 6392 -5904 6472 -5894
rect 6392 -5964 6402 -5904
rect 6462 -5914 6472 -5904
rect 6712 -5904 6792 -5894
rect 6712 -5914 6722 -5904
rect 6462 -5964 6722 -5914
rect 6782 -5964 6792 -5904
rect 6392 -5974 6792 -5964
rect 6850 -5554 7250 -5544
rect 6850 -5614 6860 -5554
rect 6920 -5604 7180 -5554
rect 6920 -5614 6930 -5604
rect 6850 -5624 6930 -5614
rect 7170 -5614 7180 -5604
rect 7240 -5614 7250 -5554
rect 7170 -5624 7250 -5614
rect 6850 -5894 6910 -5624
rect 7180 -5634 7250 -5624
rect 6990 -5684 7020 -5664
rect 6970 -5724 7020 -5684
rect 7080 -5684 7110 -5664
rect 7080 -5724 7130 -5684
rect 6970 -5794 7130 -5724
rect 6970 -5834 7020 -5794
rect 6990 -5854 7020 -5834
rect 7080 -5834 7130 -5794
rect 7080 -5854 7110 -5834
rect 7190 -5894 7250 -5634
rect 6850 -5904 6930 -5894
rect 6850 -5964 6860 -5904
rect 6920 -5914 6930 -5904
rect 7170 -5904 7250 -5894
rect 7170 -5914 7180 -5904
rect 6920 -5964 7180 -5914
rect 7240 -5964 7250 -5904
rect 6850 -5974 7250 -5964
rect 7306 -5554 7706 -5544
rect 7306 -5614 7316 -5554
rect 7376 -5604 7636 -5554
rect 7376 -5614 7386 -5604
rect 7306 -5624 7386 -5614
rect 7626 -5614 7636 -5604
rect 7696 -5614 7706 -5554
rect 7626 -5624 7706 -5614
rect 7306 -5894 7366 -5624
rect 7636 -5634 7706 -5624
rect 7446 -5684 7476 -5664
rect 7426 -5724 7476 -5684
rect 7536 -5684 7566 -5664
rect 7536 -5724 7586 -5684
rect 7426 -5794 7586 -5724
rect 7426 -5834 7476 -5794
rect 7446 -5854 7476 -5834
rect 7536 -5834 7586 -5794
rect 7536 -5854 7566 -5834
rect 7646 -5894 7706 -5634
rect 7306 -5904 7386 -5894
rect 7306 -5964 7316 -5904
rect 7376 -5914 7386 -5904
rect 7626 -5904 7706 -5894
rect 7626 -5914 7636 -5904
rect 7376 -5964 7636 -5914
rect 7696 -5964 7706 -5904
rect 7306 -5974 7706 -5964
rect 7762 -5554 8162 -5544
rect 7762 -5614 7772 -5554
rect 7832 -5604 8092 -5554
rect 7832 -5614 7842 -5604
rect 7762 -5624 7842 -5614
rect 8082 -5614 8092 -5604
rect 8152 -5614 8162 -5554
rect 8082 -5624 8162 -5614
rect 7762 -5894 7822 -5624
rect 8092 -5634 8162 -5624
rect 7902 -5684 7932 -5664
rect 7882 -5724 7932 -5684
rect 7992 -5684 8022 -5664
rect 7992 -5724 8042 -5684
rect 7882 -5794 8042 -5724
rect 7882 -5834 7932 -5794
rect 7902 -5854 7932 -5834
rect 7992 -5834 8042 -5794
rect 7992 -5854 8022 -5834
rect 8102 -5894 8162 -5634
rect 7762 -5904 7842 -5894
rect 7762 -5964 7772 -5904
rect 7832 -5914 7842 -5904
rect 8082 -5904 8162 -5894
rect 8082 -5914 8092 -5904
rect 7832 -5964 8092 -5914
rect 8152 -5964 8162 -5904
rect 7762 -5974 8162 -5964
rect 8236 -5554 8636 -5544
rect 8236 -5614 8246 -5554
rect 8306 -5604 8566 -5554
rect 8306 -5614 8316 -5604
rect 8236 -5624 8316 -5614
rect 8556 -5614 8566 -5604
rect 8626 -5614 8636 -5554
rect 8556 -5624 8636 -5614
rect 8236 -5894 8296 -5624
rect 8566 -5634 8636 -5624
rect 8376 -5684 8406 -5664
rect 8356 -5724 8406 -5684
rect 8466 -5684 8496 -5664
rect 8466 -5724 8516 -5684
rect 8356 -5794 8516 -5724
rect 8356 -5834 8406 -5794
rect 8376 -5854 8406 -5834
rect 8466 -5834 8516 -5794
rect 8466 -5854 8496 -5834
rect 8576 -5894 8636 -5634
rect 8236 -5904 8316 -5894
rect 8236 -5964 8246 -5904
rect 8306 -5914 8316 -5904
rect 8556 -5904 8636 -5894
rect 8556 -5914 8566 -5904
rect 8306 -5964 8566 -5914
rect 8626 -5964 8636 -5904
rect 8236 -5974 8636 -5964
rect 8692 -5554 9092 -5544
rect 8692 -5614 8702 -5554
rect 8762 -5604 9022 -5554
rect 8762 -5614 8772 -5604
rect 8692 -5624 8772 -5614
rect 9012 -5614 9022 -5604
rect 9082 -5614 9092 -5554
rect 9012 -5624 9092 -5614
rect 8692 -5894 8752 -5624
rect 9022 -5634 9092 -5624
rect 8832 -5684 8862 -5664
rect 8812 -5724 8862 -5684
rect 8922 -5684 8952 -5664
rect 8922 -5724 8972 -5684
rect 8812 -5794 8972 -5724
rect 8812 -5834 8862 -5794
rect 8832 -5854 8862 -5834
rect 8922 -5834 8972 -5794
rect 8922 -5854 8952 -5834
rect 9032 -5894 9092 -5634
rect 8692 -5904 8772 -5894
rect 8692 -5964 8702 -5904
rect 8762 -5914 8772 -5904
rect 9012 -5904 9092 -5894
rect 9012 -5914 9022 -5904
rect 8762 -5964 9022 -5914
rect 9082 -5964 9092 -5904
rect 8692 -5974 9092 -5964
rect 9150 -5554 9550 -5544
rect 9150 -5614 9160 -5554
rect 9220 -5604 9480 -5554
rect 9220 -5614 9230 -5604
rect 9150 -5624 9230 -5614
rect 9470 -5614 9480 -5604
rect 9540 -5614 9550 -5554
rect 9470 -5624 9550 -5614
rect 9150 -5894 9210 -5624
rect 9480 -5634 9550 -5624
rect 9290 -5684 9320 -5664
rect 9270 -5724 9320 -5684
rect 9380 -5684 9410 -5664
rect 9380 -5724 9430 -5684
rect 9270 -5794 9430 -5724
rect 9270 -5834 9320 -5794
rect 9290 -5854 9320 -5834
rect 9380 -5834 9430 -5794
rect 9380 -5854 9410 -5834
rect 9490 -5894 9550 -5634
rect 9150 -5904 9230 -5894
rect 9150 -5964 9160 -5904
rect 9220 -5914 9230 -5904
rect 9470 -5904 9550 -5894
rect 9470 -5914 9480 -5904
rect 9220 -5964 9480 -5914
rect 9540 -5964 9550 -5904
rect 9150 -5974 9550 -5964
rect 9606 -5554 10006 -5544
rect 9606 -5614 9616 -5554
rect 9676 -5604 9936 -5554
rect 9676 -5614 9686 -5604
rect 9606 -5624 9686 -5614
rect 9926 -5614 9936 -5604
rect 9996 -5614 10006 -5554
rect 9926 -5624 10006 -5614
rect 9606 -5894 9666 -5624
rect 9936 -5634 10006 -5624
rect 9746 -5684 9776 -5664
rect 9726 -5724 9776 -5684
rect 9836 -5684 9866 -5664
rect 9836 -5724 9886 -5684
rect 9726 -5794 9886 -5724
rect 9726 -5834 9776 -5794
rect 9746 -5854 9776 -5834
rect 9836 -5834 9886 -5794
rect 9836 -5854 9866 -5834
rect 9946 -5894 10006 -5634
rect 9606 -5904 9686 -5894
rect 9606 -5964 9616 -5904
rect 9676 -5914 9686 -5904
rect 9926 -5904 10006 -5894
rect 9926 -5914 9936 -5904
rect 9676 -5964 9936 -5914
rect 9996 -5964 10006 -5904
rect 9606 -5974 10006 -5964
rect 10062 -5554 10462 -5544
rect 10062 -5614 10072 -5554
rect 10132 -5604 10392 -5554
rect 10132 -5614 10142 -5604
rect 10062 -5624 10142 -5614
rect 10382 -5614 10392 -5604
rect 10452 -5614 10462 -5554
rect 10382 -5624 10462 -5614
rect 10062 -5894 10122 -5624
rect 10392 -5634 10462 -5624
rect 10202 -5684 10232 -5664
rect 10182 -5724 10232 -5684
rect 10292 -5684 10322 -5664
rect 10292 -5724 10342 -5684
rect 10182 -5794 10342 -5724
rect 10182 -5834 10232 -5794
rect 10202 -5854 10232 -5834
rect 10292 -5834 10342 -5794
rect 10292 -5854 10322 -5834
rect 10402 -5894 10462 -5634
rect 10062 -5904 10142 -5894
rect 10062 -5964 10072 -5904
rect 10132 -5914 10142 -5904
rect 10382 -5904 10462 -5894
rect 10382 -5914 10392 -5904
rect 10132 -5964 10392 -5914
rect 10452 -5964 10462 -5904
rect 10062 -5974 10462 -5964
rect 10520 -5554 10920 -5544
rect 10520 -5614 10530 -5554
rect 10590 -5604 10850 -5554
rect 10590 -5614 10600 -5604
rect 10520 -5624 10600 -5614
rect 10840 -5614 10850 -5604
rect 10910 -5614 10920 -5554
rect 10840 -5624 10920 -5614
rect 10520 -5894 10580 -5624
rect 10850 -5634 10920 -5624
rect 10660 -5684 10690 -5664
rect 10640 -5724 10690 -5684
rect 10750 -5684 10780 -5664
rect 10750 -5724 10800 -5684
rect 10640 -5794 10800 -5724
rect 10640 -5834 10690 -5794
rect 10660 -5854 10690 -5834
rect 10750 -5834 10800 -5794
rect 10750 -5854 10780 -5834
rect 10860 -5894 10920 -5634
rect 10520 -5904 10600 -5894
rect 10520 -5964 10530 -5904
rect 10590 -5914 10600 -5904
rect 10840 -5904 10920 -5894
rect 10840 -5914 10850 -5904
rect 10590 -5964 10850 -5914
rect 10910 -5964 10920 -5904
rect 10520 -5974 10920 -5964
rect 10976 -5554 11376 -5544
rect 10976 -5614 10986 -5554
rect 11046 -5604 11306 -5554
rect 11046 -5614 11056 -5604
rect 10976 -5624 11056 -5614
rect 11296 -5614 11306 -5604
rect 11366 -5614 11376 -5554
rect 11296 -5624 11376 -5614
rect 10976 -5894 11036 -5624
rect 11306 -5634 11376 -5624
rect 11116 -5684 11146 -5664
rect 11096 -5724 11146 -5684
rect 11206 -5684 11236 -5664
rect 11206 -5724 11256 -5684
rect 11096 -5794 11256 -5724
rect 11096 -5834 11146 -5794
rect 11116 -5854 11146 -5834
rect 11206 -5834 11256 -5794
rect 11206 -5854 11236 -5834
rect 11316 -5894 11376 -5634
rect 10976 -5904 11056 -5894
rect 10976 -5964 10986 -5904
rect 11046 -5914 11056 -5904
rect 11296 -5904 11376 -5894
rect 11296 -5914 11306 -5904
rect 11046 -5964 11306 -5914
rect 11366 -5964 11376 -5904
rect 10976 -5974 11376 -5964
rect 11432 -5554 11832 -5544
rect 11432 -5614 11442 -5554
rect 11502 -5604 11762 -5554
rect 11502 -5614 11512 -5604
rect 11432 -5624 11512 -5614
rect 11752 -5614 11762 -5604
rect 11822 -5614 11832 -5554
rect 11752 -5624 11832 -5614
rect 11432 -5894 11492 -5624
rect 11762 -5634 11832 -5624
rect 11572 -5684 11602 -5664
rect 11552 -5724 11602 -5684
rect 11662 -5684 11692 -5664
rect 11662 -5724 11712 -5684
rect 11552 -5794 11712 -5724
rect 11552 -5834 11602 -5794
rect 11572 -5854 11602 -5834
rect 11662 -5834 11712 -5794
rect 11662 -5854 11692 -5834
rect 11772 -5894 11832 -5634
rect 11432 -5904 11512 -5894
rect 11432 -5964 11442 -5904
rect 11502 -5914 11512 -5904
rect 11752 -5904 11832 -5894
rect 11752 -5914 11762 -5904
rect 11502 -5964 11762 -5914
rect 11822 -5964 11832 -5904
rect 11432 -5974 11832 -5964
rect 11890 -5554 12290 -5544
rect 11890 -5614 11900 -5554
rect 11960 -5604 12220 -5554
rect 11960 -5614 11970 -5604
rect 11890 -5624 11970 -5614
rect 12210 -5614 12220 -5604
rect 12280 -5614 12290 -5554
rect 12210 -5624 12290 -5614
rect 11890 -5894 11950 -5624
rect 12220 -5634 12290 -5624
rect 12030 -5684 12060 -5664
rect 12010 -5724 12060 -5684
rect 12120 -5684 12150 -5664
rect 12120 -5724 12170 -5684
rect 12010 -5794 12170 -5724
rect 12010 -5834 12060 -5794
rect 12030 -5854 12060 -5834
rect 12120 -5834 12170 -5794
rect 12120 -5854 12150 -5834
rect 12230 -5894 12290 -5634
rect 11890 -5904 11970 -5894
rect 11890 -5964 11900 -5904
rect 11960 -5914 11970 -5904
rect 12210 -5904 12290 -5894
rect 12210 -5914 12220 -5904
rect 11960 -5964 12220 -5914
rect 12280 -5964 12290 -5904
rect 11890 -5974 12290 -5964
rect 12346 -5554 12746 -5544
rect 12346 -5614 12356 -5554
rect 12416 -5604 12676 -5554
rect 12416 -5614 12426 -5604
rect 12346 -5624 12426 -5614
rect 12666 -5614 12676 -5604
rect 12736 -5614 12746 -5554
rect 12666 -5624 12746 -5614
rect 12346 -5894 12406 -5624
rect 12676 -5634 12746 -5624
rect 12486 -5684 12516 -5664
rect 12466 -5724 12516 -5684
rect 12576 -5684 12606 -5664
rect 12576 -5724 12626 -5684
rect 12466 -5794 12626 -5724
rect 12466 -5834 12516 -5794
rect 12486 -5854 12516 -5834
rect 12576 -5834 12626 -5794
rect 12576 -5854 12606 -5834
rect 12686 -5894 12746 -5634
rect 12346 -5904 12426 -5894
rect 12346 -5964 12356 -5904
rect 12416 -5914 12426 -5904
rect 12666 -5904 12746 -5894
rect 12666 -5914 12676 -5904
rect 12416 -5964 12676 -5914
rect 12736 -5964 12746 -5904
rect 12346 -5974 12746 -5964
rect 12802 -5554 13202 -5544
rect 12802 -5614 12812 -5554
rect 12872 -5604 13132 -5554
rect 12872 -5614 12882 -5604
rect 12802 -5624 12882 -5614
rect 13122 -5614 13132 -5604
rect 13192 -5614 13202 -5554
rect 13122 -5624 13202 -5614
rect 12802 -5894 12862 -5624
rect 13132 -5634 13202 -5624
rect 12942 -5684 12972 -5664
rect 12922 -5724 12972 -5684
rect 13032 -5684 13062 -5664
rect 13032 -5724 13082 -5684
rect 12922 -5794 13082 -5724
rect 12922 -5834 12972 -5794
rect 12942 -5854 12972 -5834
rect 13032 -5834 13082 -5794
rect 13032 -5854 13062 -5834
rect 13142 -5894 13202 -5634
rect 12802 -5904 12882 -5894
rect 12802 -5964 12812 -5904
rect 12872 -5914 12882 -5904
rect 13122 -5904 13202 -5894
rect 13122 -5914 13132 -5904
rect 12872 -5964 13132 -5914
rect 13192 -5964 13202 -5904
rect 12802 -5974 13202 -5964
rect 13260 -5554 13660 -5544
rect 13260 -5614 13270 -5554
rect 13330 -5604 13590 -5554
rect 13330 -5614 13340 -5604
rect 13260 -5624 13340 -5614
rect 13580 -5614 13590 -5604
rect 13650 -5614 13660 -5554
rect 13580 -5624 13660 -5614
rect 13260 -5894 13320 -5624
rect 13590 -5634 13660 -5624
rect 13400 -5684 13430 -5664
rect 13380 -5724 13430 -5684
rect 13490 -5684 13520 -5664
rect 13490 -5724 13540 -5684
rect 13380 -5794 13540 -5724
rect 13380 -5834 13430 -5794
rect 13400 -5854 13430 -5834
rect 13490 -5834 13540 -5794
rect 13490 -5854 13520 -5834
rect 13600 -5894 13660 -5634
rect 13260 -5904 13340 -5894
rect 13260 -5964 13270 -5904
rect 13330 -5914 13340 -5904
rect 13580 -5904 13660 -5894
rect 13580 -5914 13590 -5904
rect 13330 -5964 13590 -5914
rect 13650 -5964 13660 -5904
rect 13260 -5974 13660 -5964
rect 13716 -5554 14116 -5544
rect 13716 -5614 13726 -5554
rect 13786 -5604 14046 -5554
rect 13786 -5614 13796 -5604
rect 13716 -5624 13796 -5614
rect 14036 -5614 14046 -5604
rect 14106 -5614 14116 -5554
rect 14036 -5624 14116 -5614
rect 13716 -5894 13776 -5624
rect 14046 -5634 14116 -5624
rect 13856 -5684 13886 -5664
rect 13836 -5724 13886 -5684
rect 13946 -5684 13976 -5664
rect 13946 -5724 13996 -5684
rect 13836 -5794 13996 -5724
rect 13836 -5834 13886 -5794
rect 13856 -5854 13886 -5834
rect 13946 -5834 13996 -5794
rect 13946 -5854 13976 -5834
rect 14056 -5894 14116 -5634
rect 13716 -5904 13796 -5894
rect 13716 -5964 13726 -5904
rect 13786 -5914 13796 -5904
rect 14036 -5904 14116 -5894
rect 14036 -5914 14046 -5904
rect 13786 -5964 14046 -5914
rect 14106 -5964 14116 -5904
rect 13716 -5974 14116 -5964
rect 14172 -5554 14572 -5544
rect 14172 -5614 14182 -5554
rect 14242 -5604 14502 -5554
rect 14242 -5614 14252 -5604
rect 14172 -5624 14252 -5614
rect 14492 -5614 14502 -5604
rect 14562 -5614 14572 -5554
rect 14492 -5624 14572 -5614
rect 14172 -5894 14232 -5624
rect 14502 -5634 14572 -5624
rect 14312 -5684 14342 -5664
rect 14292 -5724 14342 -5684
rect 14402 -5684 14432 -5664
rect 14402 -5724 14452 -5684
rect 14292 -5794 14452 -5724
rect 14292 -5834 14342 -5794
rect 14312 -5854 14342 -5834
rect 14402 -5834 14452 -5794
rect 14402 -5854 14432 -5834
rect 14512 -5894 14572 -5634
rect 14172 -5904 14252 -5894
rect 14172 -5964 14182 -5904
rect 14242 -5914 14252 -5904
rect 14492 -5904 14572 -5894
rect 14492 -5914 14502 -5904
rect 14242 -5964 14502 -5914
rect 14562 -5964 14572 -5904
rect 14172 -5974 14572 -5964
rect 14630 -5554 15030 -5544
rect 14630 -5614 14640 -5554
rect 14700 -5604 14960 -5554
rect 14700 -5614 14710 -5604
rect 14630 -5624 14710 -5614
rect 14950 -5614 14960 -5604
rect 15020 -5614 15030 -5554
rect 14950 -5624 15030 -5614
rect 14630 -5894 14690 -5624
rect 14960 -5634 15030 -5624
rect 14770 -5684 14800 -5664
rect 14750 -5724 14800 -5684
rect 14860 -5684 14890 -5664
rect 14860 -5724 14910 -5684
rect 14750 -5794 14910 -5724
rect 14750 -5834 14800 -5794
rect 14770 -5854 14800 -5834
rect 14860 -5834 14910 -5794
rect 14860 -5854 14890 -5834
rect 14970 -5894 15030 -5634
rect 14630 -5904 14710 -5894
rect 14630 -5964 14640 -5904
rect 14700 -5914 14710 -5904
rect 14950 -5904 15030 -5894
rect 14950 -5914 14960 -5904
rect 14700 -5964 14960 -5914
rect 15020 -5964 15030 -5904
rect 14630 -5974 15030 -5964
rect 15086 -5554 15486 -5544
rect 15086 -5614 15096 -5554
rect 15156 -5604 15416 -5554
rect 15156 -5614 15166 -5604
rect 15086 -5624 15166 -5614
rect 15406 -5614 15416 -5604
rect 15476 -5614 15486 -5554
rect 15406 -5624 15486 -5614
rect 15086 -5894 15146 -5624
rect 15416 -5634 15486 -5624
rect 15226 -5684 15256 -5664
rect 15206 -5724 15256 -5684
rect 15316 -5684 15346 -5664
rect 15316 -5724 15366 -5684
rect 15206 -5794 15366 -5724
rect 15206 -5834 15256 -5794
rect 15226 -5854 15256 -5834
rect 15316 -5834 15366 -5794
rect 15316 -5854 15346 -5834
rect 15426 -5894 15486 -5634
rect 15086 -5904 15166 -5894
rect 15086 -5964 15096 -5904
rect 15156 -5914 15166 -5904
rect 15406 -5904 15486 -5894
rect 15406 -5914 15416 -5904
rect 15156 -5964 15416 -5914
rect 15476 -5964 15486 -5904
rect 15086 -5974 15486 -5964
rect 1 -6051 401 -6041
rect 1 -6111 11 -6051
rect 71 -6101 331 -6051
rect 71 -6111 81 -6101
rect 1 -6121 81 -6111
rect 321 -6111 331 -6101
rect 391 -6111 401 -6051
rect 321 -6121 401 -6111
rect 1 -6391 61 -6121
rect 331 -6131 401 -6121
rect 141 -6181 171 -6161
rect 121 -6221 171 -6181
rect 231 -6181 261 -6161
rect 231 -6221 281 -6181
rect 121 -6291 281 -6221
rect 121 -6331 171 -6291
rect 141 -6351 171 -6331
rect 231 -6331 281 -6291
rect 231 -6351 261 -6331
rect 341 -6391 401 -6131
rect 1 -6401 81 -6391
rect 1 -6461 11 -6401
rect 71 -6411 81 -6401
rect 321 -6401 401 -6391
rect 321 -6411 331 -6401
rect 71 -6461 331 -6411
rect 391 -6461 401 -6401
rect 1 -6471 401 -6461
rect 457 -6051 857 -6041
rect 457 -6111 467 -6051
rect 527 -6101 787 -6051
rect 527 -6111 537 -6101
rect 457 -6121 537 -6111
rect 777 -6111 787 -6101
rect 847 -6111 857 -6051
rect 777 -6121 857 -6111
rect 457 -6391 517 -6121
rect 787 -6131 857 -6121
rect 597 -6181 627 -6161
rect 577 -6221 627 -6181
rect 687 -6181 717 -6161
rect 687 -6221 737 -6181
rect 577 -6291 737 -6221
rect 577 -6331 627 -6291
rect 597 -6351 627 -6331
rect 687 -6331 737 -6291
rect 687 -6351 717 -6331
rect 797 -6391 857 -6131
rect 457 -6401 537 -6391
rect 457 -6461 467 -6401
rect 527 -6411 537 -6401
rect 777 -6401 857 -6391
rect 777 -6411 787 -6401
rect 527 -6461 787 -6411
rect 847 -6461 857 -6401
rect 457 -6471 857 -6461
rect 913 -6051 1313 -6041
rect 913 -6111 923 -6051
rect 983 -6101 1243 -6051
rect 983 -6111 993 -6101
rect 913 -6121 993 -6111
rect 1233 -6111 1243 -6101
rect 1303 -6111 1313 -6051
rect 1233 -6121 1313 -6111
rect 913 -6391 973 -6121
rect 1243 -6131 1313 -6121
rect 1053 -6181 1083 -6161
rect 1033 -6221 1083 -6181
rect 1143 -6181 1173 -6161
rect 1143 -6221 1193 -6181
rect 1033 -6291 1193 -6221
rect 1033 -6331 1083 -6291
rect 1053 -6351 1083 -6331
rect 1143 -6331 1193 -6291
rect 1143 -6351 1173 -6331
rect 1253 -6391 1313 -6131
rect 913 -6401 993 -6391
rect 913 -6461 923 -6401
rect 983 -6411 993 -6401
rect 1233 -6401 1313 -6391
rect 1233 -6411 1243 -6401
rect 983 -6461 1243 -6411
rect 1303 -6461 1313 -6401
rect 913 -6471 1313 -6461
rect 1371 -6051 1771 -6041
rect 1371 -6111 1381 -6051
rect 1441 -6101 1701 -6051
rect 1441 -6111 1451 -6101
rect 1371 -6121 1451 -6111
rect 1691 -6111 1701 -6101
rect 1761 -6111 1771 -6051
rect 1691 -6121 1771 -6111
rect 1371 -6391 1431 -6121
rect 1701 -6131 1771 -6121
rect 1511 -6181 1541 -6161
rect 1491 -6221 1541 -6181
rect 1601 -6181 1631 -6161
rect 1601 -6221 1651 -6181
rect 1491 -6291 1651 -6221
rect 1491 -6331 1541 -6291
rect 1511 -6351 1541 -6331
rect 1601 -6331 1651 -6291
rect 1601 -6351 1631 -6331
rect 1711 -6391 1771 -6131
rect 1371 -6401 1451 -6391
rect 1371 -6461 1381 -6401
rect 1441 -6411 1451 -6401
rect 1691 -6401 1771 -6391
rect 1691 -6411 1701 -6401
rect 1441 -6461 1701 -6411
rect 1761 -6461 1771 -6401
rect 1371 -6471 1771 -6461
rect 1827 -6051 2227 -6041
rect 1827 -6111 1837 -6051
rect 1897 -6101 2157 -6051
rect 1897 -6111 1907 -6101
rect 1827 -6121 1907 -6111
rect 2147 -6111 2157 -6101
rect 2217 -6111 2227 -6051
rect 2147 -6121 2227 -6111
rect 1827 -6391 1887 -6121
rect 2157 -6131 2227 -6121
rect 1967 -6181 1997 -6161
rect 1947 -6221 1997 -6181
rect 2057 -6181 2087 -6161
rect 2057 -6221 2107 -6181
rect 1947 -6291 2107 -6221
rect 1947 -6331 1997 -6291
rect 1967 -6351 1997 -6331
rect 2057 -6331 2107 -6291
rect 2057 -6351 2087 -6331
rect 2167 -6391 2227 -6131
rect 1827 -6401 1907 -6391
rect 1827 -6461 1837 -6401
rect 1897 -6411 1907 -6401
rect 2147 -6401 2227 -6391
rect 2147 -6411 2157 -6401
rect 1897 -6461 2157 -6411
rect 2217 -6461 2227 -6401
rect 1827 -6471 2227 -6461
rect 2283 -6051 2683 -6041
rect 2283 -6111 2293 -6051
rect 2353 -6101 2613 -6051
rect 2353 -6111 2363 -6101
rect 2283 -6121 2363 -6111
rect 2603 -6111 2613 -6101
rect 2673 -6111 2683 -6051
rect 2603 -6121 2683 -6111
rect 2283 -6391 2343 -6121
rect 2613 -6131 2683 -6121
rect 2423 -6181 2453 -6161
rect 2403 -6221 2453 -6181
rect 2513 -6181 2543 -6161
rect 2513 -6221 2563 -6181
rect 2403 -6291 2563 -6221
rect 2403 -6331 2453 -6291
rect 2423 -6351 2453 -6331
rect 2513 -6331 2563 -6291
rect 2513 -6351 2543 -6331
rect 2623 -6391 2683 -6131
rect 2283 -6401 2363 -6391
rect 2283 -6461 2293 -6401
rect 2353 -6411 2363 -6401
rect 2603 -6401 2683 -6391
rect 2603 -6411 2613 -6401
rect 2353 -6461 2613 -6411
rect 2673 -6461 2683 -6401
rect 2283 -6471 2683 -6461
rect 2741 -6051 3141 -6041
rect 2741 -6111 2751 -6051
rect 2811 -6101 3071 -6051
rect 2811 -6111 2821 -6101
rect 2741 -6121 2821 -6111
rect 3061 -6111 3071 -6101
rect 3131 -6111 3141 -6051
rect 3061 -6121 3141 -6111
rect 2741 -6391 2801 -6121
rect 3071 -6131 3141 -6121
rect 2881 -6181 2911 -6161
rect 2861 -6221 2911 -6181
rect 2971 -6181 3001 -6161
rect 2971 -6221 3021 -6181
rect 2861 -6291 3021 -6221
rect 2861 -6331 2911 -6291
rect 2881 -6351 2911 -6331
rect 2971 -6331 3021 -6291
rect 2971 -6351 3001 -6331
rect 3081 -6391 3141 -6131
rect 2741 -6401 2821 -6391
rect 2741 -6461 2751 -6401
rect 2811 -6411 2821 -6401
rect 3061 -6401 3141 -6391
rect 3061 -6411 3071 -6401
rect 2811 -6461 3071 -6411
rect 3131 -6461 3141 -6401
rect 2741 -6471 3141 -6461
rect 3197 -6051 3597 -6041
rect 3197 -6111 3207 -6051
rect 3267 -6101 3527 -6051
rect 3267 -6111 3277 -6101
rect 3197 -6121 3277 -6111
rect 3517 -6111 3527 -6101
rect 3587 -6111 3597 -6051
rect 3517 -6121 3597 -6111
rect 3197 -6391 3257 -6121
rect 3527 -6131 3597 -6121
rect 3337 -6181 3367 -6161
rect 3317 -6221 3367 -6181
rect 3427 -6181 3457 -6161
rect 3427 -6221 3477 -6181
rect 3317 -6291 3477 -6221
rect 3317 -6331 3367 -6291
rect 3337 -6351 3367 -6331
rect 3427 -6331 3477 -6291
rect 3427 -6351 3457 -6331
rect 3537 -6391 3597 -6131
rect 3197 -6401 3277 -6391
rect 3197 -6461 3207 -6401
rect 3267 -6411 3277 -6401
rect 3517 -6401 3597 -6391
rect 3517 -6411 3527 -6401
rect 3267 -6461 3527 -6411
rect 3587 -6461 3597 -6401
rect 3197 -6471 3597 -6461
rect 3653 -6051 4053 -6041
rect 3653 -6111 3663 -6051
rect 3723 -6101 3983 -6051
rect 3723 -6111 3733 -6101
rect 3653 -6121 3733 -6111
rect 3973 -6111 3983 -6101
rect 4043 -6111 4053 -6051
rect 3973 -6121 4053 -6111
rect 3653 -6391 3713 -6121
rect 3983 -6131 4053 -6121
rect 3793 -6181 3823 -6161
rect 3773 -6221 3823 -6181
rect 3883 -6181 3913 -6161
rect 3883 -6221 3933 -6181
rect 3773 -6291 3933 -6221
rect 3773 -6331 3823 -6291
rect 3793 -6351 3823 -6331
rect 3883 -6331 3933 -6291
rect 3883 -6351 3913 -6331
rect 3993 -6391 4053 -6131
rect 3653 -6401 3733 -6391
rect 3653 -6461 3663 -6401
rect 3723 -6411 3733 -6401
rect 3973 -6401 4053 -6391
rect 3973 -6411 3983 -6401
rect 3723 -6461 3983 -6411
rect 4043 -6461 4053 -6401
rect 3653 -6471 4053 -6461
rect 4111 -6051 4511 -6041
rect 4111 -6111 4121 -6051
rect 4181 -6101 4441 -6051
rect 4181 -6111 4191 -6101
rect 4111 -6121 4191 -6111
rect 4431 -6111 4441 -6101
rect 4501 -6111 4511 -6051
rect 4431 -6121 4511 -6111
rect 4111 -6391 4171 -6121
rect 4441 -6131 4511 -6121
rect 4251 -6181 4281 -6161
rect 4231 -6221 4281 -6181
rect 4341 -6181 4371 -6161
rect 4341 -6221 4391 -6181
rect 4231 -6291 4391 -6221
rect 4231 -6331 4281 -6291
rect 4251 -6351 4281 -6331
rect 4341 -6331 4391 -6291
rect 4341 -6351 4371 -6331
rect 4451 -6391 4511 -6131
rect 4111 -6401 4191 -6391
rect 4111 -6461 4121 -6401
rect 4181 -6411 4191 -6401
rect 4431 -6401 4511 -6391
rect 4431 -6411 4441 -6401
rect 4181 -6461 4441 -6411
rect 4501 -6461 4511 -6401
rect 4111 -6471 4511 -6461
rect 4567 -6051 4967 -6041
rect 4567 -6111 4577 -6051
rect 4637 -6101 4897 -6051
rect 4637 -6111 4647 -6101
rect 4567 -6121 4647 -6111
rect 4887 -6111 4897 -6101
rect 4957 -6111 4967 -6051
rect 4887 -6121 4967 -6111
rect 4567 -6391 4627 -6121
rect 4897 -6131 4967 -6121
rect 4707 -6181 4737 -6161
rect 4687 -6221 4737 -6181
rect 4797 -6181 4827 -6161
rect 4797 -6221 4847 -6181
rect 4687 -6291 4847 -6221
rect 4687 -6331 4737 -6291
rect 4707 -6351 4737 -6331
rect 4797 -6331 4847 -6291
rect 4797 -6351 4827 -6331
rect 4907 -6391 4967 -6131
rect 4567 -6401 4647 -6391
rect 4567 -6461 4577 -6401
rect 4637 -6411 4647 -6401
rect 4887 -6401 4967 -6391
rect 4887 -6411 4897 -6401
rect 4637 -6461 4897 -6411
rect 4957 -6461 4967 -6401
rect 4567 -6471 4967 -6461
rect 5023 -6051 5423 -6041
rect 5023 -6111 5033 -6051
rect 5093 -6101 5353 -6051
rect 5093 -6111 5103 -6101
rect 5023 -6121 5103 -6111
rect 5343 -6111 5353 -6101
rect 5413 -6111 5423 -6051
rect 5343 -6121 5423 -6111
rect 5023 -6391 5083 -6121
rect 5353 -6131 5423 -6121
rect 5163 -6181 5193 -6161
rect 5143 -6221 5193 -6181
rect 5253 -6181 5283 -6161
rect 5253 -6221 5303 -6181
rect 5143 -6291 5303 -6221
rect 5143 -6331 5193 -6291
rect 5163 -6351 5193 -6331
rect 5253 -6331 5303 -6291
rect 5253 -6351 5283 -6331
rect 5363 -6391 5423 -6131
rect 5023 -6401 5103 -6391
rect 5023 -6461 5033 -6401
rect 5093 -6411 5103 -6401
rect 5343 -6401 5423 -6391
rect 5343 -6411 5353 -6401
rect 5093 -6461 5353 -6411
rect 5413 -6461 5423 -6401
rect 5023 -6471 5423 -6461
rect 5481 -6051 5881 -6041
rect 5481 -6111 5491 -6051
rect 5551 -6101 5811 -6051
rect 5551 -6111 5561 -6101
rect 5481 -6121 5561 -6111
rect 5801 -6111 5811 -6101
rect 5871 -6111 5881 -6051
rect 5801 -6121 5881 -6111
rect 5481 -6391 5541 -6121
rect 5811 -6131 5881 -6121
rect 5621 -6181 5651 -6161
rect 5601 -6221 5651 -6181
rect 5711 -6181 5741 -6161
rect 5711 -6221 5761 -6181
rect 5601 -6291 5761 -6221
rect 5601 -6331 5651 -6291
rect 5621 -6351 5651 -6331
rect 5711 -6331 5761 -6291
rect 5711 -6351 5741 -6331
rect 5821 -6391 5881 -6131
rect 5481 -6401 5561 -6391
rect 5481 -6461 5491 -6401
rect 5551 -6411 5561 -6401
rect 5801 -6401 5881 -6391
rect 5801 -6411 5811 -6401
rect 5551 -6461 5811 -6411
rect 5871 -6461 5881 -6401
rect 5481 -6471 5881 -6461
rect 5937 -6051 6337 -6041
rect 5937 -6111 5947 -6051
rect 6007 -6101 6267 -6051
rect 6007 -6111 6017 -6101
rect 5937 -6121 6017 -6111
rect 6257 -6111 6267 -6101
rect 6327 -6111 6337 -6051
rect 6257 -6121 6337 -6111
rect 5937 -6391 5997 -6121
rect 6267 -6131 6337 -6121
rect 6077 -6181 6107 -6161
rect 6057 -6221 6107 -6181
rect 6167 -6181 6197 -6161
rect 6167 -6221 6217 -6181
rect 6057 -6291 6217 -6221
rect 6057 -6331 6107 -6291
rect 6077 -6351 6107 -6331
rect 6167 -6331 6217 -6291
rect 6167 -6351 6197 -6331
rect 6277 -6391 6337 -6131
rect 5937 -6401 6017 -6391
rect 5937 -6461 5947 -6401
rect 6007 -6411 6017 -6401
rect 6257 -6401 6337 -6391
rect 6257 -6411 6267 -6401
rect 6007 -6461 6267 -6411
rect 6327 -6461 6337 -6401
rect 5937 -6471 6337 -6461
rect 6393 -6051 6793 -6041
rect 6393 -6111 6403 -6051
rect 6463 -6101 6723 -6051
rect 6463 -6111 6473 -6101
rect 6393 -6121 6473 -6111
rect 6713 -6111 6723 -6101
rect 6783 -6111 6793 -6051
rect 6713 -6121 6793 -6111
rect 6393 -6391 6453 -6121
rect 6723 -6131 6793 -6121
rect 6533 -6181 6563 -6161
rect 6513 -6221 6563 -6181
rect 6623 -6181 6653 -6161
rect 6623 -6221 6673 -6181
rect 6513 -6291 6673 -6221
rect 6513 -6331 6563 -6291
rect 6533 -6351 6563 -6331
rect 6623 -6331 6673 -6291
rect 6623 -6351 6653 -6331
rect 6733 -6391 6793 -6131
rect 6393 -6401 6473 -6391
rect 6393 -6461 6403 -6401
rect 6463 -6411 6473 -6401
rect 6713 -6401 6793 -6391
rect 6713 -6411 6723 -6401
rect 6463 -6461 6723 -6411
rect 6783 -6461 6793 -6401
rect 6393 -6471 6793 -6461
rect 6851 -6051 7251 -6041
rect 6851 -6111 6861 -6051
rect 6921 -6101 7181 -6051
rect 6921 -6111 6931 -6101
rect 6851 -6121 6931 -6111
rect 7171 -6111 7181 -6101
rect 7241 -6111 7251 -6051
rect 7171 -6121 7251 -6111
rect 6851 -6391 6911 -6121
rect 7181 -6131 7251 -6121
rect 6991 -6181 7021 -6161
rect 6971 -6221 7021 -6181
rect 7081 -6181 7111 -6161
rect 7081 -6221 7131 -6181
rect 6971 -6291 7131 -6221
rect 6971 -6331 7021 -6291
rect 6991 -6351 7021 -6331
rect 7081 -6331 7131 -6291
rect 7081 -6351 7111 -6331
rect 7191 -6391 7251 -6131
rect 6851 -6401 6931 -6391
rect 6851 -6461 6861 -6401
rect 6921 -6411 6931 -6401
rect 7171 -6401 7251 -6391
rect 7171 -6411 7181 -6401
rect 6921 -6461 7181 -6411
rect 7241 -6461 7251 -6401
rect 6851 -6471 7251 -6461
rect 7307 -6051 7707 -6041
rect 7307 -6111 7317 -6051
rect 7377 -6101 7637 -6051
rect 7377 -6111 7387 -6101
rect 7307 -6121 7387 -6111
rect 7627 -6111 7637 -6101
rect 7697 -6111 7707 -6051
rect 7627 -6121 7707 -6111
rect 7307 -6391 7367 -6121
rect 7637 -6131 7707 -6121
rect 7447 -6181 7477 -6161
rect 7427 -6221 7477 -6181
rect 7537 -6181 7567 -6161
rect 7537 -6221 7587 -6181
rect 7427 -6291 7587 -6221
rect 7427 -6331 7477 -6291
rect 7447 -6351 7477 -6331
rect 7537 -6331 7587 -6291
rect 7537 -6351 7567 -6331
rect 7647 -6391 7707 -6131
rect 7307 -6401 7387 -6391
rect 7307 -6461 7317 -6401
rect 7377 -6411 7387 -6401
rect 7627 -6401 7707 -6391
rect 7627 -6411 7637 -6401
rect 7377 -6461 7637 -6411
rect 7697 -6461 7707 -6401
rect 7307 -6471 7707 -6461
rect 7763 -6051 8163 -6041
rect 7763 -6111 7773 -6051
rect 7833 -6101 8093 -6051
rect 7833 -6111 7843 -6101
rect 7763 -6121 7843 -6111
rect 8083 -6111 8093 -6101
rect 8153 -6111 8163 -6051
rect 8083 -6121 8163 -6111
rect 7763 -6391 7823 -6121
rect 8093 -6131 8163 -6121
rect 7903 -6181 7933 -6161
rect 7883 -6221 7933 -6181
rect 7993 -6181 8023 -6161
rect 7993 -6221 8043 -6181
rect 7883 -6291 8043 -6221
rect 7883 -6331 7933 -6291
rect 7903 -6351 7933 -6331
rect 7993 -6331 8043 -6291
rect 7993 -6351 8023 -6331
rect 8103 -6391 8163 -6131
rect 7763 -6401 7843 -6391
rect 7763 -6461 7773 -6401
rect 7833 -6411 7843 -6401
rect 8083 -6401 8163 -6391
rect 8083 -6411 8093 -6401
rect 7833 -6461 8093 -6411
rect 8153 -6461 8163 -6401
rect 7763 -6471 8163 -6461
rect 8237 -6051 8637 -6041
rect 8237 -6111 8247 -6051
rect 8307 -6101 8567 -6051
rect 8307 -6111 8317 -6101
rect 8237 -6121 8317 -6111
rect 8557 -6111 8567 -6101
rect 8627 -6111 8637 -6051
rect 8557 -6121 8637 -6111
rect 8237 -6391 8297 -6121
rect 8567 -6131 8637 -6121
rect 8377 -6181 8407 -6161
rect 8357 -6221 8407 -6181
rect 8467 -6181 8497 -6161
rect 8467 -6221 8517 -6181
rect 8357 -6291 8517 -6221
rect 8357 -6331 8407 -6291
rect 8377 -6351 8407 -6331
rect 8467 -6331 8517 -6291
rect 8467 -6351 8497 -6331
rect 8577 -6391 8637 -6131
rect 8237 -6401 8317 -6391
rect 8237 -6461 8247 -6401
rect 8307 -6411 8317 -6401
rect 8557 -6401 8637 -6391
rect 8557 -6411 8567 -6401
rect 8307 -6461 8567 -6411
rect 8627 -6461 8637 -6401
rect 8237 -6471 8637 -6461
rect 8693 -6051 9093 -6041
rect 8693 -6111 8703 -6051
rect 8763 -6101 9023 -6051
rect 8763 -6111 8773 -6101
rect 8693 -6121 8773 -6111
rect 9013 -6111 9023 -6101
rect 9083 -6111 9093 -6051
rect 9013 -6121 9093 -6111
rect 8693 -6391 8753 -6121
rect 9023 -6131 9093 -6121
rect 8833 -6181 8863 -6161
rect 8813 -6221 8863 -6181
rect 8923 -6181 8953 -6161
rect 8923 -6221 8973 -6181
rect 8813 -6291 8973 -6221
rect 8813 -6331 8863 -6291
rect 8833 -6351 8863 -6331
rect 8923 -6331 8973 -6291
rect 8923 -6351 8953 -6331
rect 9033 -6391 9093 -6131
rect 8693 -6401 8773 -6391
rect 8693 -6461 8703 -6401
rect 8763 -6411 8773 -6401
rect 9013 -6401 9093 -6391
rect 9013 -6411 9023 -6401
rect 8763 -6461 9023 -6411
rect 9083 -6461 9093 -6401
rect 8693 -6471 9093 -6461
rect 9151 -6051 9551 -6041
rect 9151 -6111 9161 -6051
rect 9221 -6101 9481 -6051
rect 9221 -6111 9231 -6101
rect 9151 -6121 9231 -6111
rect 9471 -6111 9481 -6101
rect 9541 -6111 9551 -6051
rect 9471 -6121 9551 -6111
rect 9151 -6391 9211 -6121
rect 9481 -6131 9551 -6121
rect 9291 -6181 9321 -6161
rect 9271 -6221 9321 -6181
rect 9381 -6181 9411 -6161
rect 9381 -6221 9431 -6181
rect 9271 -6291 9431 -6221
rect 9271 -6331 9321 -6291
rect 9291 -6351 9321 -6331
rect 9381 -6331 9431 -6291
rect 9381 -6351 9411 -6331
rect 9491 -6391 9551 -6131
rect 9151 -6401 9231 -6391
rect 9151 -6461 9161 -6401
rect 9221 -6411 9231 -6401
rect 9471 -6401 9551 -6391
rect 9471 -6411 9481 -6401
rect 9221 -6461 9481 -6411
rect 9541 -6461 9551 -6401
rect 9151 -6471 9551 -6461
rect 9607 -6051 10007 -6041
rect 9607 -6111 9617 -6051
rect 9677 -6101 9937 -6051
rect 9677 -6111 9687 -6101
rect 9607 -6121 9687 -6111
rect 9927 -6111 9937 -6101
rect 9997 -6111 10007 -6051
rect 9927 -6121 10007 -6111
rect 9607 -6391 9667 -6121
rect 9937 -6131 10007 -6121
rect 9747 -6181 9777 -6161
rect 9727 -6221 9777 -6181
rect 9837 -6181 9867 -6161
rect 9837 -6221 9887 -6181
rect 9727 -6291 9887 -6221
rect 9727 -6331 9777 -6291
rect 9747 -6351 9777 -6331
rect 9837 -6331 9887 -6291
rect 9837 -6351 9867 -6331
rect 9947 -6391 10007 -6131
rect 9607 -6401 9687 -6391
rect 9607 -6461 9617 -6401
rect 9677 -6411 9687 -6401
rect 9927 -6401 10007 -6391
rect 9927 -6411 9937 -6401
rect 9677 -6461 9937 -6411
rect 9997 -6461 10007 -6401
rect 9607 -6471 10007 -6461
rect 10063 -6051 10463 -6041
rect 10063 -6111 10073 -6051
rect 10133 -6101 10393 -6051
rect 10133 -6111 10143 -6101
rect 10063 -6121 10143 -6111
rect 10383 -6111 10393 -6101
rect 10453 -6111 10463 -6051
rect 10383 -6121 10463 -6111
rect 10063 -6391 10123 -6121
rect 10393 -6131 10463 -6121
rect 10203 -6181 10233 -6161
rect 10183 -6221 10233 -6181
rect 10293 -6181 10323 -6161
rect 10293 -6221 10343 -6181
rect 10183 -6291 10343 -6221
rect 10183 -6331 10233 -6291
rect 10203 -6351 10233 -6331
rect 10293 -6331 10343 -6291
rect 10293 -6351 10323 -6331
rect 10403 -6391 10463 -6131
rect 10063 -6401 10143 -6391
rect 10063 -6461 10073 -6401
rect 10133 -6411 10143 -6401
rect 10383 -6401 10463 -6391
rect 10383 -6411 10393 -6401
rect 10133 -6461 10393 -6411
rect 10453 -6461 10463 -6401
rect 10063 -6471 10463 -6461
rect 10521 -6051 10921 -6041
rect 10521 -6111 10531 -6051
rect 10591 -6101 10851 -6051
rect 10591 -6111 10601 -6101
rect 10521 -6121 10601 -6111
rect 10841 -6111 10851 -6101
rect 10911 -6111 10921 -6051
rect 10841 -6121 10921 -6111
rect 10521 -6391 10581 -6121
rect 10851 -6131 10921 -6121
rect 10661 -6181 10691 -6161
rect 10641 -6221 10691 -6181
rect 10751 -6181 10781 -6161
rect 10751 -6221 10801 -6181
rect 10641 -6291 10801 -6221
rect 10641 -6331 10691 -6291
rect 10661 -6351 10691 -6331
rect 10751 -6331 10801 -6291
rect 10751 -6351 10781 -6331
rect 10861 -6391 10921 -6131
rect 10521 -6401 10601 -6391
rect 10521 -6461 10531 -6401
rect 10591 -6411 10601 -6401
rect 10841 -6401 10921 -6391
rect 10841 -6411 10851 -6401
rect 10591 -6461 10851 -6411
rect 10911 -6461 10921 -6401
rect 10521 -6471 10921 -6461
rect 10977 -6051 11377 -6041
rect 10977 -6111 10987 -6051
rect 11047 -6101 11307 -6051
rect 11047 -6111 11057 -6101
rect 10977 -6121 11057 -6111
rect 11297 -6111 11307 -6101
rect 11367 -6111 11377 -6051
rect 11297 -6121 11377 -6111
rect 10977 -6391 11037 -6121
rect 11307 -6131 11377 -6121
rect 11117 -6181 11147 -6161
rect 11097 -6221 11147 -6181
rect 11207 -6181 11237 -6161
rect 11207 -6221 11257 -6181
rect 11097 -6291 11257 -6221
rect 11097 -6331 11147 -6291
rect 11117 -6351 11147 -6331
rect 11207 -6331 11257 -6291
rect 11207 -6351 11237 -6331
rect 11317 -6391 11377 -6131
rect 10977 -6401 11057 -6391
rect 10977 -6461 10987 -6401
rect 11047 -6411 11057 -6401
rect 11297 -6401 11377 -6391
rect 11297 -6411 11307 -6401
rect 11047 -6461 11307 -6411
rect 11367 -6461 11377 -6401
rect 10977 -6471 11377 -6461
rect 11433 -6051 11833 -6041
rect 11433 -6111 11443 -6051
rect 11503 -6101 11763 -6051
rect 11503 -6111 11513 -6101
rect 11433 -6121 11513 -6111
rect 11753 -6111 11763 -6101
rect 11823 -6111 11833 -6051
rect 11753 -6121 11833 -6111
rect 11433 -6391 11493 -6121
rect 11763 -6131 11833 -6121
rect 11573 -6181 11603 -6161
rect 11553 -6221 11603 -6181
rect 11663 -6181 11693 -6161
rect 11663 -6221 11713 -6181
rect 11553 -6291 11713 -6221
rect 11553 -6331 11603 -6291
rect 11573 -6351 11603 -6331
rect 11663 -6331 11713 -6291
rect 11663 -6351 11693 -6331
rect 11773 -6391 11833 -6131
rect 11433 -6401 11513 -6391
rect 11433 -6461 11443 -6401
rect 11503 -6411 11513 -6401
rect 11753 -6401 11833 -6391
rect 11753 -6411 11763 -6401
rect 11503 -6461 11763 -6411
rect 11823 -6461 11833 -6401
rect 11433 -6471 11833 -6461
rect 11891 -6051 12291 -6041
rect 11891 -6111 11901 -6051
rect 11961 -6101 12221 -6051
rect 11961 -6111 11971 -6101
rect 11891 -6121 11971 -6111
rect 12211 -6111 12221 -6101
rect 12281 -6111 12291 -6051
rect 12211 -6121 12291 -6111
rect 11891 -6391 11951 -6121
rect 12221 -6131 12291 -6121
rect 12031 -6181 12061 -6161
rect 12011 -6221 12061 -6181
rect 12121 -6181 12151 -6161
rect 12121 -6221 12171 -6181
rect 12011 -6291 12171 -6221
rect 12011 -6331 12061 -6291
rect 12031 -6351 12061 -6331
rect 12121 -6331 12171 -6291
rect 12121 -6351 12151 -6331
rect 12231 -6391 12291 -6131
rect 11891 -6401 11971 -6391
rect 11891 -6461 11901 -6401
rect 11961 -6411 11971 -6401
rect 12211 -6401 12291 -6391
rect 12211 -6411 12221 -6401
rect 11961 -6461 12221 -6411
rect 12281 -6461 12291 -6401
rect 11891 -6471 12291 -6461
rect 12347 -6051 12747 -6041
rect 12347 -6111 12357 -6051
rect 12417 -6101 12677 -6051
rect 12417 -6111 12427 -6101
rect 12347 -6121 12427 -6111
rect 12667 -6111 12677 -6101
rect 12737 -6111 12747 -6051
rect 12667 -6121 12747 -6111
rect 12347 -6391 12407 -6121
rect 12677 -6131 12747 -6121
rect 12487 -6181 12517 -6161
rect 12467 -6221 12517 -6181
rect 12577 -6181 12607 -6161
rect 12577 -6221 12627 -6181
rect 12467 -6291 12627 -6221
rect 12467 -6331 12517 -6291
rect 12487 -6351 12517 -6331
rect 12577 -6331 12627 -6291
rect 12577 -6351 12607 -6331
rect 12687 -6391 12747 -6131
rect 12347 -6401 12427 -6391
rect 12347 -6461 12357 -6401
rect 12417 -6411 12427 -6401
rect 12667 -6401 12747 -6391
rect 12667 -6411 12677 -6401
rect 12417 -6461 12677 -6411
rect 12737 -6461 12747 -6401
rect 12347 -6471 12747 -6461
rect 12803 -6051 13203 -6041
rect 12803 -6111 12813 -6051
rect 12873 -6101 13133 -6051
rect 12873 -6111 12883 -6101
rect 12803 -6121 12883 -6111
rect 13123 -6111 13133 -6101
rect 13193 -6111 13203 -6051
rect 13123 -6121 13203 -6111
rect 12803 -6391 12863 -6121
rect 13133 -6131 13203 -6121
rect 12943 -6181 12973 -6161
rect 12923 -6221 12973 -6181
rect 13033 -6181 13063 -6161
rect 13033 -6221 13083 -6181
rect 12923 -6291 13083 -6221
rect 12923 -6331 12973 -6291
rect 12943 -6351 12973 -6331
rect 13033 -6331 13083 -6291
rect 13033 -6351 13063 -6331
rect 13143 -6391 13203 -6131
rect 12803 -6401 12883 -6391
rect 12803 -6461 12813 -6401
rect 12873 -6411 12883 -6401
rect 13123 -6401 13203 -6391
rect 13123 -6411 13133 -6401
rect 12873 -6461 13133 -6411
rect 13193 -6461 13203 -6401
rect 12803 -6471 13203 -6461
rect 13261 -6051 13661 -6041
rect 13261 -6111 13271 -6051
rect 13331 -6101 13591 -6051
rect 13331 -6111 13341 -6101
rect 13261 -6121 13341 -6111
rect 13581 -6111 13591 -6101
rect 13651 -6111 13661 -6051
rect 13581 -6121 13661 -6111
rect 13261 -6391 13321 -6121
rect 13591 -6131 13661 -6121
rect 13401 -6181 13431 -6161
rect 13381 -6221 13431 -6181
rect 13491 -6181 13521 -6161
rect 13491 -6221 13541 -6181
rect 13381 -6291 13541 -6221
rect 13381 -6331 13431 -6291
rect 13401 -6351 13431 -6331
rect 13491 -6331 13541 -6291
rect 13491 -6351 13521 -6331
rect 13601 -6391 13661 -6131
rect 13261 -6401 13341 -6391
rect 13261 -6461 13271 -6401
rect 13331 -6411 13341 -6401
rect 13581 -6401 13661 -6391
rect 13581 -6411 13591 -6401
rect 13331 -6461 13591 -6411
rect 13651 -6461 13661 -6401
rect 13261 -6471 13661 -6461
rect 13717 -6051 14117 -6041
rect 13717 -6111 13727 -6051
rect 13787 -6101 14047 -6051
rect 13787 -6111 13797 -6101
rect 13717 -6121 13797 -6111
rect 14037 -6111 14047 -6101
rect 14107 -6111 14117 -6051
rect 14037 -6121 14117 -6111
rect 13717 -6391 13777 -6121
rect 14047 -6131 14117 -6121
rect 13857 -6181 13887 -6161
rect 13837 -6221 13887 -6181
rect 13947 -6181 13977 -6161
rect 13947 -6221 13997 -6181
rect 13837 -6291 13997 -6221
rect 13837 -6331 13887 -6291
rect 13857 -6351 13887 -6331
rect 13947 -6331 13997 -6291
rect 13947 -6351 13977 -6331
rect 14057 -6391 14117 -6131
rect 13717 -6401 13797 -6391
rect 13717 -6461 13727 -6401
rect 13787 -6411 13797 -6401
rect 14037 -6401 14117 -6391
rect 14037 -6411 14047 -6401
rect 13787 -6461 14047 -6411
rect 14107 -6461 14117 -6401
rect 13717 -6471 14117 -6461
rect 14173 -6051 14573 -6041
rect 14173 -6111 14183 -6051
rect 14243 -6101 14503 -6051
rect 14243 -6111 14253 -6101
rect 14173 -6121 14253 -6111
rect 14493 -6111 14503 -6101
rect 14563 -6111 14573 -6051
rect 14493 -6121 14573 -6111
rect 14173 -6391 14233 -6121
rect 14503 -6131 14573 -6121
rect 14313 -6181 14343 -6161
rect 14293 -6221 14343 -6181
rect 14403 -6181 14433 -6161
rect 14403 -6221 14453 -6181
rect 14293 -6291 14453 -6221
rect 14293 -6331 14343 -6291
rect 14313 -6351 14343 -6331
rect 14403 -6331 14453 -6291
rect 14403 -6351 14433 -6331
rect 14513 -6391 14573 -6131
rect 14173 -6401 14253 -6391
rect 14173 -6461 14183 -6401
rect 14243 -6411 14253 -6401
rect 14493 -6401 14573 -6391
rect 14493 -6411 14503 -6401
rect 14243 -6461 14503 -6411
rect 14563 -6461 14573 -6401
rect 14173 -6471 14573 -6461
rect 14631 -6051 15031 -6041
rect 14631 -6111 14641 -6051
rect 14701 -6101 14961 -6051
rect 14701 -6111 14711 -6101
rect 14631 -6121 14711 -6111
rect 14951 -6111 14961 -6101
rect 15021 -6111 15031 -6051
rect 14951 -6121 15031 -6111
rect 14631 -6391 14691 -6121
rect 14961 -6131 15031 -6121
rect 14771 -6181 14801 -6161
rect 14751 -6221 14801 -6181
rect 14861 -6181 14891 -6161
rect 14861 -6221 14911 -6181
rect 14751 -6291 14911 -6221
rect 14751 -6331 14801 -6291
rect 14771 -6351 14801 -6331
rect 14861 -6331 14911 -6291
rect 14861 -6351 14891 -6331
rect 14971 -6391 15031 -6131
rect 14631 -6401 14711 -6391
rect 14631 -6461 14641 -6401
rect 14701 -6411 14711 -6401
rect 14951 -6401 15031 -6391
rect 14951 -6411 14961 -6401
rect 14701 -6461 14961 -6411
rect 15021 -6461 15031 -6401
rect 14631 -6471 15031 -6461
rect 15087 -6051 15487 -6041
rect 15087 -6111 15097 -6051
rect 15157 -6101 15417 -6051
rect 15157 -6111 15167 -6101
rect 15087 -6121 15167 -6111
rect 15407 -6111 15417 -6101
rect 15477 -6111 15487 -6051
rect 15407 -6121 15487 -6111
rect 15087 -6391 15147 -6121
rect 15417 -6131 15487 -6121
rect 15227 -6181 15257 -6161
rect 15207 -6221 15257 -6181
rect 15317 -6181 15347 -6161
rect 15317 -6221 15367 -6181
rect 15207 -6291 15367 -6221
rect 15207 -6331 15257 -6291
rect 15227 -6351 15257 -6331
rect 15317 -6331 15367 -6291
rect 15317 -6351 15347 -6331
rect 15427 -6391 15487 -6131
rect 15087 -6401 15167 -6391
rect 15087 -6461 15097 -6401
rect 15157 -6411 15167 -6401
rect 15407 -6401 15487 -6391
rect 15407 -6411 15417 -6401
rect 15157 -6461 15417 -6411
rect 15477 -6461 15487 -6401
rect 15087 -6471 15487 -6461
rect 1 -6543 401 -6533
rect 1 -6603 11 -6543
rect 71 -6593 331 -6543
rect 71 -6603 81 -6593
rect 1 -6613 81 -6603
rect 321 -6603 331 -6593
rect 391 -6603 401 -6543
rect 321 -6613 401 -6603
rect 1 -6883 61 -6613
rect 331 -6623 401 -6613
rect 141 -6673 171 -6653
rect 121 -6713 171 -6673
rect 231 -6673 261 -6653
rect 231 -6713 281 -6673
rect 121 -6783 281 -6713
rect 121 -6823 171 -6783
rect 141 -6843 171 -6823
rect 231 -6823 281 -6783
rect 231 -6843 261 -6823
rect 341 -6883 401 -6623
rect 1 -6893 81 -6883
rect 1 -6953 11 -6893
rect 71 -6903 81 -6893
rect 321 -6893 401 -6883
rect 321 -6903 331 -6893
rect 71 -6953 331 -6903
rect 391 -6953 401 -6893
rect 1 -6963 401 -6953
rect 457 -6543 857 -6533
rect 457 -6603 467 -6543
rect 527 -6593 787 -6543
rect 527 -6603 537 -6593
rect 457 -6613 537 -6603
rect 777 -6603 787 -6593
rect 847 -6603 857 -6543
rect 777 -6613 857 -6603
rect 457 -6883 517 -6613
rect 787 -6623 857 -6613
rect 597 -6673 627 -6653
rect 577 -6713 627 -6673
rect 687 -6673 717 -6653
rect 687 -6713 737 -6673
rect 577 -6783 737 -6713
rect 577 -6823 627 -6783
rect 597 -6843 627 -6823
rect 687 -6823 737 -6783
rect 687 -6843 717 -6823
rect 797 -6883 857 -6623
rect 457 -6893 537 -6883
rect 457 -6953 467 -6893
rect 527 -6903 537 -6893
rect 777 -6893 857 -6883
rect 777 -6903 787 -6893
rect 527 -6953 787 -6903
rect 847 -6953 857 -6893
rect 457 -6963 857 -6953
rect 913 -6543 1313 -6533
rect 913 -6603 923 -6543
rect 983 -6593 1243 -6543
rect 983 -6603 993 -6593
rect 913 -6613 993 -6603
rect 1233 -6603 1243 -6593
rect 1303 -6603 1313 -6543
rect 1233 -6613 1313 -6603
rect 913 -6883 973 -6613
rect 1243 -6623 1313 -6613
rect 1053 -6673 1083 -6653
rect 1033 -6713 1083 -6673
rect 1143 -6673 1173 -6653
rect 1143 -6713 1193 -6673
rect 1033 -6783 1193 -6713
rect 1033 -6823 1083 -6783
rect 1053 -6843 1083 -6823
rect 1143 -6823 1193 -6783
rect 1143 -6843 1173 -6823
rect 1253 -6883 1313 -6623
rect 913 -6893 993 -6883
rect 913 -6953 923 -6893
rect 983 -6903 993 -6893
rect 1233 -6893 1313 -6883
rect 1233 -6903 1243 -6893
rect 983 -6953 1243 -6903
rect 1303 -6953 1313 -6893
rect 913 -6963 1313 -6953
rect 1371 -6543 1771 -6533
rect 1371 -6603 1381 -6543
rect 1441 -6593 1701 -6543
rect 1441 -6603 1451 -6593
rect 1371 -6613 1451 -6603
rect 1691 -6603 1701 -6593
rect 1761 -6603 1771 -6543
rect 1691 -6613 1771 -6603
rect 1371 -6883 1431 -6613
rect 1701 -6623 1771 -6613
rect 1511 -6673 1541 -6653
rect 1491 -6713 1541 -6673
rect 1601 -6673 1631 -6653
rect 1601 -6713 1651 -6673
rect 1491 -6783 1651 -6713
rect 1491 -6823 1541 -6783
rect 1511 -6843 1541 -6823
rect 1601 -6823 1651 -6783
rect 1601 -6843 1631 -6823
rect 1711 -6883 1771 -6623
rect 1371 -6893 1451 -6883
rect 1371 -6953 1381 -6893
rect 1441 -6903 1451 -6893
rect 1691 -6893 1771 -6883
rect 1691 -6903 1701 -6893
rect 1441 -6953 1701 -6903
rect 1761 -6953 1771 -6893
rect 1371 -6963 1771 -6953
rect 1827 -6543 2227 -6533
rect 1827 -6603 1837 -6543
rect 1897 -6593 2157 -6543
rect 1897 -6603 1907 -6593
rect 1827 -6613 1907 -6603
rect 2147 -6603 2157 -6593
rect 2217 -6603 2227 -6543
rect 2147 -6613 2227 -6603
rect 1827 -6883 1887 -6613
rect 2157 -6623 2227 -6613
rect 1967 -6673 1997 -6653
rect 1947 -6713 1997 -6673
rect 2057 -6673 2087 -6653
rect 2057 -6713 2107 -6673
rect 1947 -6783 2107 -6713
rect 1947 -6823 1997 -6783
rect 1967 -6843 1997 -6823
rect 2057 -6823 2107 -6783
rect 2057 -6843 2087 -6823
rect 2167 -6883 2227 -6623
rect 1827 -6893 1907 -6883
rect 1827 -6953 1837 -6893
rect 1897 -6903 1907 -6893
rect 2147 -6893 2227 -6883
rect 2147 -6903 2157 -6893
rect 1897 -6953 2157 -6903
rect 2217 -6953 2227 -6893
rect 1827 -6963 2227 -6953
rect 2283 -6543 2683 -6533
rect 2283 -6603 2293 -6543
rect 2353 -6593 2613 -6543
rect 2353 -6603 2363 -6593
rect 2283 -6613 2363 -6603
rect 2603 -6603 2613 -6593
rect 2673 -6603 2683 -6543
rect 2603 -6613 2683 -6603
rect 2283 -6883 2343 -6613
rect 2613 -6623 2683 -6613
rect 2423 -6673 2453 -6653
rect 2403 -6713 2453 -6673
rect 2513 -6673 2543 -6653
rect 2513 -6713 2563 -6673
rect 2403 -6783 2563 -6713
rect 2403 -6823 2453 -6783
rect 2423 -6843 2453 -6823
rect 2513 -6823 2563 -6783
rect 2513 -6843 2543 -6823
rect 2623 -6883 2683 -6623
rect 2283 -6893 2363 -6883
rect 2283 -6953 2293 -6893
rect 2353 -6903 2363 -6893
rect 2603 -6893 2683 -6883
rect 2603 -6903 2613 -6893
rect 2353 -6953 2613 -6903
rect 2673 -6953 2683 -6893
rect 2283 -6963 2683 -6953
rect 2741 -6543 3141 -6533
rect 2741 -6603 2751 -6543
rect 2811 -6593 3071 -6543
rect 2811 -6603 2821 -6593
rect 2741 -6613 2821 -6603
rect 3061 -6603 3071 -6593
rect 3131 -6603 3141 -6543
rect 3061 -6613 3141 -6603
rect 2741 -6883 2801 -6613
rect 3071 -6623 3141 -6613
rect 2881 -6673 2911 -6653
rect 2861 -6713 2911 -6673
rect 2971 -6673 3001 -6653
rect 2971 -6713 3021 -6673
rect 2861 -6783 3021 -6713
rect 2861 -6823 2911 -6783
rect 2881 -6843 2911 -6823
rect 2971 -6823 3021 -6783
rect 2971 -6843 3001 -6823
rect 3081 -6883 3141 -6623
rect 2741 -6893 2821 -6883
rect 2741 -6953 2751 -6893
rect 2811 -6903 2821 -6893
rect 3061 -6893 3141 -6883
rect 3061 -6903 3071 -6893
rect 2811 -6953 3071 -6903
rect 3131 -6953 3141 -6893
rect 2741 -6963 3141 -6953
rect 3197 -6543 3597 -6533
rect 3197 -6603 3207 -6543
rect 3267 -6593 3527 -6543
rect 3267 -6603 3277 -6593
rect 3197 -6613 3277 -6603
rect 3517 -6603 3527 -6593
rect 3587 -6603 3597 -6543
rect 3517 -6613 3597 -6603
rect 3197 -6883 3257 -6613
rect 3527 -6623 3597 -6613
rect 3337 -6673 3367 -6653
rect 3317 -6713 3367 -6673
rect 3427 -6673 3457 -6653
rect 3427 -6713 3477 -6673
rect 3317 -6783 3477 -6713
rect 3317 -6823 3367 -6783
rect 3337 -6843 3367 -6823
rect 3427 -6823 3477 -6783
rect 3427 -6843 3457 -6823
rect 3537 -6883 3597 -6623
rect 3197 -6893 3277 -6883
rect 3197 -6953 3207 -6893
rect 3267 -6903 3277 -6893
rect 3517 -6893 3597 -6883
rect 3517 -6903 3527 -6893
rect 3267 -6953 3527 -6903
rect 3587 -6953 3597 -6893
rect 3197 -6963 3597 -6953
rect 3653 -6543 4053 -6533
rect 3653 -6603 3663 -6543
rect 3723 -6593 3983 -6543
rect 3723 -6603 3733 -6593
rect 3653 -6613 3733 -6603
rect 3973 -6603 3983 -6593
rect 4043 -6603 4053 -6543
rect 3973 -6613 4053 -6603
rect 3653 -6883 3713 -6613
rect 3983 -6623 4053 -6613
rect 3793 -6673 3823 -6653
rect 3773 -6713 3823 -6673
rect 3883 -6673 3913 -6653
rect 3883 -6713 3933 -6673
rect 3773 -6783 3933 -6713
rect 3773 -6823 3823 -6783
rect 3793 -6843 3823 -6823
rect 3883 -6823 3933 -6783
rect 3883 -6843 3913 -6823
rect 3993 -6883 4053 -6623
rect 3653 -6893 3733 -6883
rect 3653 -6953 3663 -6893
rect 3723 -6903 3733 -6893
rect 3973 -6893 4053 -6883
rect 3973 -6903 3983 -6893
rect 3723 -6953 3983 -6903
rect 4043 -6953 4053 -6893
rect 3653 -6963 4053 -6953
rect 4111 -6543 4511 -6533
rect 4111 -6603 4121 -6543
rect 4181 -6593 4441 -6543
rect 4181 -6603 4191 -6593
rect 4111 -6613 4191 -6603
rect 4431 -6603 4441 -6593
rect 4501 -6603 4511 -6543
rect 4431 -6613 4511 -6603
rect 4111 -6883 4171 -6613
rect 4441 -6623 4511 -6613
rect 4251 -6673 4281 -6653
rect 4231 -6713 4281 -6673
rect 4341 -6673 4371 -6653
rect 4341 -6713 4391 -6673
rect 4231 -6783 4391 -6713
rect 4231 -6823 4281 -6783
rect 4251 -6843 4281 -6823
rect 4341 -6823 4391 -6783
rect 4341 -6843 4371 -6823
rect 4451 -6883 4511 -6623
rect 4111 -6893 4191 -6883
rect 4111 -6953 4121 -6893
rect 4181 -6903 4191 -6893
rect 4431 -6893 4511 -6883
rect 4431 -6903 4441 -6893
rect 4181 -6953 4441 -6903
rect 4501 -6953 4511 -6893
rect 4111 -6963 4511 -6953
rect 4567 -6543 4967 -6533
rect 4567 -6603 4577 -6543
rect 4637 -6593 4897 -6543
rect 4637 -6603 4647 -6593
rect 4567 -6613 4647 -6603
rect 4887 -6603 4897 -6593
rect 4957 -6603 4967 -6543
rect 4887 -6613 4967 -6603
rect 4567 -6883 4627 -6613
rect 4897 -6623 4967 -6613
rect 4707 -6673 4737 -6653
rect 4687 -6713 4737 -6673
rect 4797 -6673 4827 -6653
rect 4797 -6713 4847 -6673
rect 4687 -6783 4847 -6713
rect 4687 -6823 4737 -6783
rect 4707 -6843 4737 -6823
rect 4797 -6823 4847 -6783
rect 4797 -6843 4827 -6823
rect 4907 -6883 4967 -6623
rect 4567 -6893 4647 -6883
rect 4567 -6953 4577 -6893
rect 4637 -6903 4647 -6893
rect 4887 -6893 4967 -6883
rect 4887 -6903 4897 -6893
rect 4637 -6953 4897 -6903
rect 4957 -6953 4967 -6893
rect 4567 -6963 4967 -6953
rect 5023 -6543 5423 -6533
rect 5023 -6603 5033 -6543
rect 5093 -6593 5353 -6543
rect 5093 -6603 5103 -6593
rect 5023 -6613 5103 -6603
rect 5343 -6603 5353 -6593
rect 5413 -6603 5423 -6543
rect 5343 -6613 5423 -6603
rect 5023 -6883 5083 -6613
rect 5353 -6623 5423 -6613
rect 5163 -6673 5193 -6653
rect 5143 -6713 5193 -6673
rect 5253 -6673 5283 -6653
rect 5253 -6713 5303 -6673
rect 5143 -6783 5303 -6713
rect 5143 -6823 5193 -6783
rect 5163 -6843 5193 -6823
rect 5253 -6823 5303 -6783
rect 5253 -6843 5283 -6823
rect 5363 -6883 5423 -6623
rect 5023 -6893 5103 -6883
rect 5023 -6953 5033 -6893
rect 5093 -6903 5103 -6893
rect 5343 -6893 5423 -6883
rect 5343 -6903 5353 -6893
rect 5093 -6953 5353 -6903
rect 5413 -6953 5423 -6893
rect 5023 -6963 5423 -6953
rect 5481 -6543 5881 -6533
rect 5481 -6603 5491 -6543
rect 5551 -6593 5811 -6543
rect 5551 -6603 5561 -6593
rect 5481 -6613 5561 -6603
rect 5801 -6603 5811 -6593
rect 5871 -6603 5881 -6543
rect 5801 -6613 5881 -6603
rect 5481 -6883 5541 -6613
rect 5811 -6623 5881 -6613
rect 5621 -6673 5651 -6653
rect 5601 -6713 5651 -6673
rect 5711 -6673 5741 -6653
rect 5711 -6713 5761 -6673
rect 5601 -6783 5761 -6713
rect 5601 -6823 5651 -6783
rect 5621 -6843 5651 -6823
rect 5711 -6823 5761 -6783
rect 5711 -6843 5741 -6823
rect 5821 -6883 5881 -6623
rect 5481 -6893 5561 -6883
rect 5481 -6953 5491 -6893
rect 5551 -6903 5561 -6893
rect 5801 -6893 5881 -6883
rect 5801 -6903 5811 -6893
rect 5551 -6953 5811 -6903
rect 5871 -6953 5881 -6893
rect 5481 -6963 5881 -6953
rect 5937 -6543 6337 -6533
rect 5937 -6603 5947 -6543
rect 6007 -6593 6267 -6543
rect 6007 -6603 6017 -6593
rect 5937 -6613 6017 -6603
rect 6257 -6603 6267 -6593
rect 6327 -6603 6337 -6543
rect 6257 -6613 6337 -6603
rect 5937 -6883 5997 -6613
rect 6267 -6623 6337 -6613
rect 6077 -6673 6107 -6653
rect 6057 -6713 6107 -6673
rect 6167 -6673 6197 -6653
rect 6167 -6713 6217 -6673
rect 6057 -6783 6217 -6713
rect 6057 -6823 6107 -6783
rect 6077 -6843 6107 -6823
rect 6167 -6823 6217 -6783
rect 6167 -6843 6197 -6823
rect 6277 -6883 6337 -6623
rect 5937 -6893 6017 -6883
rect 5937 -6953 5947 -6893
rect 6007 -6903 6017 -6893
rect 6257 -6893 6337 -6883
rect 6257 -6903 6267 -6893
rect 6007 -6953 6267 -6903
rect 6327 -6953 6337 -6893
rect 5937 -6963 6337 -6953
rect 6393 -6543 6793 -6533
rect 6393 -6603 6403 -6543
rect 6463 -6593 6723 -6543
rect 6463 -6603 6473 -6593
rect 6393 -6613 6473 -6603
rect 6713 -6603 6723 -6593
rect 6783 -6603 6793 -6543
rect 6713 -6613 6793 -6603
rect 6393 -6883 6453 -6613
rect 6723 -6623 6793 -6613
rect 6533 -6673 6563 -6653
rect 6513 -6713 6563 -6673
rect 6623 -6673 6653 -6653
rect 6623 -6713 6673 -6673
rect 6513 -6783 6673 -6713
rect 6513 -6823 6563 -6783
rect 6533 -6843 6563 -6823
rect 6623 -6823 6673 -6783
rect 6623 -6843 6653 -6823
rect 6733 -6883 6793 -6623
rect 6393 -6893 6473 -6883
rect 6393 -6953 6403 -6893
rect 6463 -6903 6473 -6893
rect 6713 -6893 6793 -6883
rect 6713 -6903 6723 -6893
rect 6463 -6953 6723 -6903
rect 6783 -6953 6793 -6893
rect 6393 -6963 6793 -6953
rect 6851 -6543 7251 -6533
rect 6851 -6603 6861 -6543
rect 6921 -6593 7181 -6543
rect 6921 -6603 6931 -6593
rect 6851 -6613 6931 -6603
rect 7171 -6603 7181 -6593
rect 7241 -6603 7251 -6543
rect 7171 -6613 7251 -6603
rect 6851 -6883 6911 -6613
rect 7181 -6623 7251 -6613
rect 6991 -6673 7021 -6653
rect 6971 -6713 7021 -6673
rect 7081 -6673 7111 -6653
rect 7081 -6713 7131 -6673
rect 6971 -6783 7131 -6713
rect 6971 -6823 7021 -6783
rect 6991 -6843 7021 -6823
rect 7081 -6823 7131 -6783
rect 7081 -6843 7111 -6823
rect 7191 -6883 7251 -6623
rect 6851 -6893 6931 -6883
rect 6851 -6953 6861 -6893
rect 6921 -6903 6931 -6893
rect 7171 -6893 7251 -6883
rect 7171 -6903 7181 -6893
rect 6921 -6953 7181 -6903
rect 7241 -6953 7251 -6893
rect 6851 -6963 7251 -6953
rect 7307 -6543 7707 -6533
rect 7307 -6603 7317 -6543
rect 7377 -6593 7637 -6543
rect 7377 -6603 7387 -6593
rect 7307 -6613 7387 -6603
rect 7627 -6603 7637 -6593
rect 7697 -6603 7707 -6543
rect 7627 -6613 7707 -6603
rect 7307 -6883 7367 -6613
rect 7637 -6623 7707 -6613
rect 7447 -6673 7477 -6653
rect 7427 -6713 7477 -6673
rect 7537 -6673 7567 -6653
rect 7537 -6713 7587 -6673
rect 7427 -6783 7587 -6713
rect 7427 -6823 7477 -6783
rect 7447 -6843 7477 -6823
rect 7537 -6823 7587 -6783
rect 7537 -6843 7567 -6823
rect 7647 -6883 7707 -6623
rect 7307 -6893 7387 -6883
rect 7307 -6953 7317 -6893
rect 7377 -6903 7387 -6893
rect 7627 -6893 7707 -6883
rect 7627 -6903 7637 -6893
rect 7377 -6953 7637 -6903
rect 7697 -6953 7707 -6893
rect 7307 -6963 7707 -6953
rect 7763 -6543 8163 -6533
rect 7763 -6603 7773 -6543
rect 7833 -6593 8093 -6543
rect 7833 -6603 7843 -6593
rect 7763 -6613 7843 -6603
rect 8083 -6603 8093 -6593
rect 8153 -6603 8163 -6543
rect 8083 -6613 8163 -6603
rect 7763 -6883 7823 -6613
rect 8093 -6623 8163 -6613
rect 7903 -6673 7933 -6653
rect 7883 -6713 7933 -6673
rect 7993 -6673 8023 -6653
rect 7993 -6713 8043 -6673
rect 7883 -6783 8043 -6713
rect 7883 -6823 7933 -6783
rect 7903 -6843 7933 -6823
rect 7993 -6823 8043 -6783
rect 7993 -6843 8023 -6823
rect 8103 -6883 8163 -6623
rect 7763 -6893 7843 -6883
rect 7763 -6953 7773 -6893
rect 7833 -6903 7843 -6893
rect 8083 -6893 8163 -6883
rect 8083 -6903 8093 -6893
rect 7833 -6953 8093 -6903
rect 8153 -6953 8163 -6893
rect 7763 -6963 8163 -6953
rect 8237 -6543 8637 -6533
rect 8237 -6603 8247 -6543
rect 8307 -6593 8567 -6543
rect 8307 -6603 8317 -6593
rect 8237 -6613 8317 -6603
rect 8557 -6603 8567 -6593
rect 8627 -6603 8637 -6543
rect 8557 -6613 8637 -6603
rect 8237 -6883 8297 -6613
rect 8567 -6623 8637 -6613
rect 8377 -6673 8407 -6653
rect 8357 -6713 8407 -6673
rect 8467 -6673 8497 -6653
rect 8467 -6713 8517 -6673
rect 8357 -6783 8517 -6713
rect 8357 -6823 8407 -6783
rect 8377 -6843 8407 -6823
rect 8467 -6823 8517 -6783
rect 8467 -6843 8497 -6823
rect 8577 -6883 8637 -6623
rect 8237 -6893 8317 -6883
rect 8237 -6953 8247 -6893
rect 8307 -6903 8317 -6893
rect 8557 -6893 8637 -6883
rect 8557 -6903 8567 -6893
rect 8307 -6953 8567 -6903
rect 8627 -6953 8637 -6893
rect 8237 -6963 8637 -6953
rect 8693 -6543 9093 -6533
rect 8693 -6603 8703 -6543
rect 8763 -6593 9023 -6543
rect 8763 -6603 8773 -6593
rect 8693 -6613 8773 -6603
rect 9013 -6603 9023 -6593
rect 9083 -6603 9093 -6543
rect 9013 -6613 9093 -6603
rect 8693 -6883 8753 -6613
rect 9023 -6623 9093 -6613
rect 8833 -6673 8863 -6653
rect 8813 -6713 8863 -6673
rect 8923 -6673 8953 -6653
rect 8923 -6713 8973 -6673
rect 8813 -6783 8973 -6713
rect 8813 -6823 8863 -6783
rect 8833 -6843 8863 -6823
rect 8923 -6823 8973 -6783
rect 8923 -6843 8953 -6823
rect 9033 -6883 9093 -6623
rect 8693 -6893 8773 -6883
rect 8693 -6953 8703 -6893
rect 8763 -6903 8773 -6893
rect 9013 -6893 9093 -6883
rect 9013 -6903 9023 -6893
rect 8763 -6953 9023 -6903
rect 9083 -6953 9093 -6893
rect 8693 -6963 9093 -6953
rect 9151 -6543 9551 -6533
rect 9151 -6603 9161 -6543
rect 9221 -6593 9481 -6543
rect 9221 -6603 9231 -6593
rect 9151 -6613 9231 -6603
rect 9471 -6603 9481 -6593
rect 9541 -6603 9551 -6543
rect 9471 -6613 9551 -6603
rect 9151 -6883 9211 -6613
rect 9481 -6623 9551 -6613
rect 9291 -6673 9321 -6653
rect 9271 -6713 9321 -6673
rect 9381 -6673 9411 -6653
rect 9381 -6713 9431 -6673
rect 9271 -6783 9431 -6713
rect 9271 -6823 9321 -6783
rect 9291 -6843 9321 -6823
rect 9381 -6823 9431 -6783
rect 9381 -6843 9411 -6823
rect 9491 -6883 9551 -6623
rect 9151 -6893 9231 -6883
rect 9151 -6953 9161 -6893
rect 9221 -6903 9231 -6893
rect 9471 -6893 9551 -6883
rect 9471 -6903 9481 -6893
rect 9221 -6953 9481 -6903
rect 9541 -6953 9551 -6893
rect 9151 -6963 9551 -6953
rect 9607 -6543 10007 -6533
rect 9607 -6603 9617 -6543
rect 9677 -6593 9937 -6543
rect 9677 -6603 9687 -6593
rect 9607 -6613 9687 -6603
rect 9927 -6603 9937 -6593
rect 9997 -6603 10007 -6543
rect 9927 -6613 10007 -6603
rect 9607 -6883 9667 -6613
rect 9937 -6623 10007 -6613
rect 9747 -6673 9777 -6653
rect 9727 -6713 9777 -6673
rect 9837 -6673 9867 -6653
rect 9837 -6713 9887 -6673
rect 9727 -6783 9887 -6713
rect 9727 -6823 9777 -6783
rect 9747 -6843 9777 -6823
rect 9837 -6823 9887 -6783
rect 9837 -6843 9867 -6823
rect 9947 -6883 10007 -6623
rect 9607 -6893 9687 -6883
rect 9607 -6953 9617 -6893
rect 9677 -6903 9687 -6893
rect 9927 -6893 10007 -6883
rect 9927 -6903 9937 -6893
rect 9677 -6953 9937 -6903
rect 9997 -6953 10007 -6893
rect 9607 -6963 10007 -6953
rect 10063 -6543 10463 -6533
rect 10063 -6603 10073 -6543
rect 10133 -6593 10393 -6543
rect 10133 -6603 10143 -6593
rect 10063 -6613 10143 -6603
rect 10383 -6603 10393 -6593
rect 10453 -6603 10463 -6543
rect 10383 -6613 10463 -6603
rect 10063 -6883 10123 -6613
rect 10393 -6623 10463 -6613
rect 10203 -6673 10233 -6653
rect 10183 -6713 10233 -6673
rect 10293 -6673 10323 -6653
rect 10293 -6713 10343 -6673
rect 10183 -6783 10343 -6713
rect 10183 -6823 10233 -6783
rect 10203 -6843 10233 -6823
rect 10293 -6823 10343 -6783
rect 10293 -6843 10323 -6823
rect 10403 -6883 10463 -6623
rect 10063 -6893 10143 -6883
rect 10063 -6953 10073 -6893
rect 10133 -6903 10143 -6893
rect 10383 -6893 10463 -6883
rect 10383 -6903 10393 -6893
rect 10133 -6953 10393 -6903
rect 10453 -6953 10463 -6893
rect 10063 -6963 10463 -6953
rect 10521 -6543 10921 -6533
rect 10521 -6603 10531 -6543
rect 10591 -6593 10851 -6543
rect 10591 -6603 10601 -6593
rect 10521 -6613 10601 -6603
rect 10841 -6603 10851 -6593
rect 10911 -6603 10921 -6543
rect 10841 -6613 10921 -6603
rect 10521 -6883 10581 -6613
rect 10851 -6623 10921 -6613
rect 10661 -6673 10691 -6653
rect 10641 -6713 10691 -6673
rect 10751 -6673 10781 -6653
rect 10751 -6713 10801 -6673
rect 10641 -6783 10801 -6713
rect 10641 -6823 10691 -6783
rect 10661 -6843 10691 -6823
rect 10751 -6823 10801 -6783
rect 10751 -6843 10781 -6823
rect 10861 -6883 10921 -6623
rect 10521 -6893 10601 -6883
rect 10521 -6953 10531 -6893
rect 10591 -6903 10601 -6893
rect 10841 -6893 10921 -6883
rect 10841 -6903 10851 -6893
rect 10591 -6953 10851 -6903
rect 10911 -6953 10921 -6893
rect 10521 -6963 10921 -6953
rect 10977 -6543 11377 -6533
rect 10977 -6603 10987 -6543
rect 11047 -6593 11307 -6543
rect 11047 -6603 11057 -6593
rect 10977 -6613 11057 -6603
rect 11297 -6603 11307 -6593
rect 11367 -6603 11377 -6543
rect 11297 -6613 11377 -6603
rect 10977 -6883 11037 -6613
rect 11307 -6623 11377 -6613
rect 11117 -6673 11147 -6653
rect 11097 -6713 11147 -6673
rect 11207 -6673 11237 -6653
rect 11207 -6713 11257 -6673
rect 11097 -6783 11257 -6713
rect 11097 -6823 11147 -6783
rect 11117 -6843 11147 -6823
rect 11207 -6823 11257 -6783
rect 11207 -6843 11237 -6823
rect 11317 -6883 11377 -6623
rect 10977 -6893 11057 -6883
rect 10977 -6953 10987 -6893
rect 11047 -6903 11057 -6893
rect 11297 -6893 11377 -6883
rect 11297 -6903 11307 -6893
rect 11047 -6953 11307 -6903
rect 11367 -6953 11377 -6893
rect 10977 -6963 11377 -6953
rect 11433 -6543 11833 -6533
rect 11433 -6603 11443 -6543
rect 11503 -6593 11763 -6543
rect 11503 -6603 11513 -6593
rect 11433 -6613 11513 -6603
rect 11753 -6603 11763 -6593
rect 11823 -6603 11833 -6543
rect 11753 -6613 11833 -6603
rect 11433 -6883 11493 -6613
rect 11763 -6623 11833 -6613
rect 11573 -6673 11603 -6653
rect 11553 -6713 11603 -6673
rect 11663 -6673 11693 -6653
rect 11663 -6713 11713 -6673
rect 11553 -6783 11713 -6713
rect 11553 -6823 11603 -6783
rect 11573 -6843 11603 -6823
rect 11663 -6823 11713 -6783
rect 11663 -6843 11693 -6823
rect 11773 -6883 11833 -6623
rect 11433 -6893 11513 -6883
rect 11433 -6953 11443 -6893
rect 11503 -6903 11513 -6893
rect 11753 -6893 11833 -6883
rect 11753 -6903 11763 -6893
rect 11503 -6953 11763 -6903
rect 11823 -6953 11833 -6893
rect 11433 -6963 11833 -6953
rect 11891 -6543 12291 -6533
rect 11891 -6603 11901 -6543
rect 11961 -6593 12221 -6543
rect 11961 -6603 11971 -6593
rect 11891 -6613 11971 -6603
rect 12211 -6603 12221 -6593
rect 12281 -6603 12291 -6543
rect 12211 -6613 12291 -6603
rect 11891 -6883 11951 -6613
rect 12221 -6623 12291 -6613
rect 12031 -6673 12061 -6653
rect 12011 -6713 12061 -6673
rect 12121 -6673 12151 -6653
rect 12121 -6713 12171 -6673
rect 12011 -6783 12171 -6713
rect 12011 -6823 12061 -6783
rect 12031 -6843 12061 -6823
rect 12121 -6823 12171 -6783
rect 12121 -6843 12151 -6823
rect 12231 -6883 12291 -6623
rect 11891 -6893 11971 -6883
rect 11891 -6953 11901 -6893
rect 11961 -6903 11971 -6893
rect 12211 -6893 12291 -6883
rect 12211 -6903 12221 -6893
rect 11961 -6953 12221 -6903
rect 12281 -6953 12291 -6893
rect 11891 -6963 12291 -6953
rect 12347 -6543 12747 -6533
rect 12347 -6603 12357 -6543
rect 12417 -6593 12677 -6543
rect 12417 -6603 12427 -6593
rect 12347 -6613 12427 -6603
rect 12667 -6603 12677 -6593
rect 12737 -6603 12747 -6543
rect 12667 -6613 12747 -6603
rect 12347 -6883 12407 -6613
rect 12677 -6623 12747 -6613
rect 12487 -6673 12517 -6653
rect 12467 -6713 12517 -6673
rect 12577 -6673 12607 -6653
rect 12577 -6713 12627 -6673
rect 12467 -6783 12627 -6713
rect 12467 -6823 12517 -6783
rect 12487 -6843 12517 -6823
rect 12577 -6823 12627 -6783
rect 12577 -6843 12607 -6823
rect 12687 -6883 12747 -6623
rect 12347 -6893 12427 -6883
rect 12347 -6953 12357 -6893
rect 12417 -6903 12427 -6893
rect 12667 -6893 12747 -6883
rect 12667 -6903 12677 -6893
rect 12417 -6953 12677 -6903
rect 12737 -6953 12747 -6893
rect 12347 -6963 12747 -6953
rect 12803 -6543 13203 -6533
rect 12803 -6603 12813 -6543
rect 12873 -6593 13133 -6543
rect 12873 -6603 12883 -6593
rect 12803 -6613 12883 -6603
rect 13123 -6603 13133 -6593
rect 13193 -6603 13203 -6543
rect 13123 -6613 13203 -6603
rect 12803 -6883 12863 -6613
rect 13133 -6623 13203 -6613
rect 12943 -6673 12973 -6653
rect 12923 -6713 12973 -6673
rect 13033 -6673 13063 -6653
rect 13033 -6713 13083 -6673
rect 12923 -6783 13083 -6713
rect 12923 -6823 12973 -6783
rect 12943 -6843 12973 -6823
rect 13033 -6823 13083 -6783
rect 13033 -6843 13063 -6823
rect 13143 -6883 13203 -6623
rect 12803 -6893 12883 -6883
rect 12803 -6953 12813 -6893
rect 12873 -6903 12883 -6893
rect 13123 -6893 13203 -6883
rect 13123 -6903 13133 -6893
rect 12873 -6953 13133 -6903
rect 13193 -6953 13203 -6893
rect 12803 -6963 13203 -6953
rect 13261 -6543 13661 -6533
rect 13261 -6603 13271 -6543
rect 13331 -6593 13591 -6543
rect 13331 -6603 13341 -6593
rect 13261 -6613 13341 -6603
rect 13581 -6603 13591 -6593
rect 13651 -6603 13661 -6543
rect 13581 -6613 13661 -6603
rect 13261 -6883 13321 -6613
rect 13591 -6623 13661 -6613
rect 13401 -6673 13431 -6653
rect 13381 -6713 13431 -6673
rect 13491 -6673 13521 -6653
rect 13491 -6713 13541 -6673
rect 13381 -6783 13541 -6713
rect 13381 -6823 13431 -6783
rect 13401 -6843 13431 -6823
rect 13491 -6823 13541 -6783
rect 13491 -6843 13521 -6823
rect 13601 -6883 13661 -6623
rect 13261 -6893 13341 -6883
rect 13261 -6953 13271 -6893
rect 13331 -6903 13341 -6893
rect 13581 -6893 13661 -6883
rect 13581 -6903 13591 -6893
rect 13331 -6953 13591 -6903
rect 13651 -6953 13661 -6893
rect 13261 -6963 13661 -6953
rect 13717 -6543 14117 -6533
rect 13717 -6603 13727 -6543
rect 13787 -6593 14047 -6543
rect 13787 -6603 13797 -6593
rect 13717 -6613 13797 -6603
rect 14037 -6603 14047 -6593
rect 14107 -6603 14117 -6543
rect 14037 -6613 14117 -6603
rect 13717 -6883 13777 -6613
rect 14047 -6623 14117 -6613
rect 13857 -6673 13887 -6653
rect 13837 -6713 13887 -6673
rect 13947 -6673 13977 -6653
rect 13947 -6713 13997 -6673
rect 13837 -6783 13997 -6713
rect 13837 -6823 13887 -6783
rect 13857 -6843 13887 -6823
rect 13947 -6823 13997 -6783
rect 13947 -6843 13977 -6823
rect 14057 -6883 14117 -6623
rect 13717 -6893 13797 -6883
rect 13717 -6953 13727 -6893
rect 13787 -6903 13797 -6893
rect 14037 -6893 14117 -6883
rect 14037 -6903 14047 -6893
rect 13787 -6953 14047 -6903
rect 14107 -6953 14117 -6893
rect 13717 -6963 14117 -6953
rect 14173 -6543 14573 -6533
rect 14173 -6603 14183 -6543
rect 14243 -6593 14503 -6543
rect 14243 -6603 14253 -6593
rect 14173 -6613 14253 -6603
rect 14493 -6603 14503 -6593
rect 14563 -6603 14573 -6543
rect 14493 -6613 14573 -6603
rect 14173 -6883 14233 -6613
rect 14503 -6623 14573 -6613
rect 14313 -6673 14343 -6653
rect 14293 -6713 14343 -6673
rect 14403 -6673 14433 -6653
rect 14403 -6713 14453 -6673
rect 14293 -6783 14453 -6713
rect 14293 -6823 14343 -6783
rect 14313 -6843 14343 -6823
rect 14403 -6823 14453 -6783
rect 14403 -6843 14433 -6823
rect 14513 -6883 14573 -6623
rect 14173 -6893 14253 -6883
rect 14173 -6953 14183 -6893
rect 14243 -6903 14253 -6893
rect 14493 -6893 14573 -6883
rect 14493 -6903 14503 -6893
rect 14243 -6953 14503 -6903
rect 14563 -6953 14573 -6893
rect 14173 -6963 14573 -6953
rect 14631 -6543 15031 -6533
rect 14631 -6603 14641 -6543
rect 14701 -6593 14961 -6543
rect 14701 -6603 14711 -6593
rect 14631 -6613 14711 -6603
rect 14951 -6603 14961 -6593
rect 15021 -6603 15031 -6543
rect 14951 -6613 15031 -6603
rect 14631 -6883 14691 -6613
rect 14961 -6623 15031 -6613
rect 14771 -6673 14801 -6653
rect 14751 -6713 14801 -6673
rect 14861 -6673 14891 -6653
rect 14861 -6713 14911 -6673
rect 14751 -6783 14911 -6713
rect 14751 -6823 14801 -6783
rect 14771 -6843 14801 -6823
rect 14861 -6823 14911 -6783
rect 14861 -6843 14891 -6823
rect 14971 -6883 15031 -6623
rect 14631 -6893 14711 -6883
rect 14631 -6953 14641 -6893
rect 14701 -6903 14711 -6893
rect 14951 -6893 15031 -6883
rect 14951 -6903 14961 -6893
rect 14701 -6953 14961 -6903
rect 15021 -6953 15031 -6893
rect 14631 -6963 15031 -6953
rect 15087 -6543 15487 -6533
rect 15087 -6603 15097 -6543
rect 15157 -6593 15417 -6543
rect 15157 -6603 15167 -6593
rect 15087 -6613 15167 -6603
rect 15407 -6603 15417 -6593
rect 15477 -6603 15487 -6543
rect 15407 -6613 15487 -6603
rect 15087 -6883 15147 -6613
rect 15417 -6623 15487 -6613
rect 15227 -6673 15257 -6653
rect 15207 -6713 15257 -6673
rect 15317 -6673 15347 -6653
rect 15317 -6713 15367 -6673
rect 15207 -6783 15367 -6713
rect 15207 -6823 15257 -6783
rect 15227 -6843 15257 -6823
rect 15317 -6823 15367 -6783
rect 15317 -6843 15347 -6823
rect 15427 -6883 15487 -6623
rect 15087 -6893 15167 -6883
rect 15087 -6953 15097 -6893
rect 15157 -6903 15167 -6893
rect 15407 -6893 15487 -6883
rect 15407 -6903 15417 -6893
rect 15157 -6953 15417 -6903
rect 15477 -6953 15487 -6893
rect 15087 -6963 15487 -6953
rect 1 -7059 401 -7049
rect 1 -7119 11 -7059
rect 71 -7109 331 -7059
rect 71 -7119 81 -7109
rect 1 -7129 81 -7119
rect 321 -7119 331 -7109
rect 391 -7119 401 -7059
rect 321 -7129 401 -7119
rect 1 -7399 61 -7129
rect 331 -7139 401 -7129
rect 141 -7189 171 -7169
rect 121 -7229 171 -7189
rect 231 -7189 261 -7169
rect 231 -7229 281 -7189
rect 121 -7299 281 -7229
rect 121 -7339 171 -7299
rect 141 -7359 171 -7339
rect 231 -7339 281 -7299
rect 231 -7359 261 -7339
rect 341 -7399 401 -7139
rect 1 -7409 81 -7399
rect 1 -7469 11 -7409
rect 71 -7419 81 -7409
rect 321 -7409 401 -7399
rect 321 -7419 331 -7409
rect 71 -7469 331 -7419
rect 391 -7469 401 -7409
rect 1 -7479 401 -7469
rect 457 -7059 857 -7049
rect 457 -7119 467 -7059
rect 527 -7109 787 -7059
rect 527 -7119 537 -7109
rect 457 -7129 537 -7119
rect 777 -7119 787 -7109
rect 847 -7119 857 -7059
rect 777 -7129 857 -7119
rect 457 -7399 517 -7129
rect 787 -7139 857 -7129
rect 597 -7189 627 -7169
rect 577 -7229 627 -7189
rect 687 -7189 717 -7169
rect 687 -7229 737 -7189
rect 577 -7299 737 -7229
rect 577 -7339 627 -7299
rect 597 -7359 627 -7339
rect 687 -7339 737 -7299
rect 687 -7359 717 -7339
rect 797 -7399 857 -7139
rect 457 -7409 537 -7399
rect 457 -7469 467 -7409
rect 527 -7419 537 -7409
rect 777 -7409 857 -7399
rect 777 -7419 787 -7409
rect 527 -7469 787 -7419
rect 847 -7469 857 -7409
rect 457 -7479 857 -7469
rect 913 -7059 1313 -7049
rect 913 -7119 923 -7059
rect 983 -7109 1243 -7059
rect 983 -7119 993 -7109
rect 913 -7129 993 -7119
rect 1233 -7119 1243 -7109
rect 1303 -7119 1313 -7059
rect 1233 -7129 1313 -7119
rect 913 -7399 973 -7129
rect 1243 -7139 1313 -7129
rect 1053 -7189 1083 -7169
rect 1033 -7229 1083 -7189
rect 1143 -7189 1173 -7169
rect 1143 -7229 1193 -7189
rect 1033 -7299 1193 -7229
rect 1033 -7339 1083 -7299
rect 1053 -7359 1083 -7339
rect 1143 -7339 1193 -7299
rect 1143 -7359 1173 -7339
rect 1253 -7399 1313 -7139
rect 913 -7409 993 -7399
rect 913 -7469 923 -7409
rect 983 -7419 993 -7409
rect 1233 -7409 1313 -7399
rect 1233 -7419 1243 -7409
rect 983 -7469 1243 -7419
rect 1303 -7469 1313 -7409
rect 913 -7479 1313 -7469
rect 1371 -7059 1771 -7049
rect 1371 -7119 1381 -7059
rect 1441 -7109 1701 -7059
rect 1441 -7119 1451 -7109
rect 1371 -7129 1451 -7119
rect 1691 -7119 1701 -7109
rect 1761 -7119 1771 -7059
rect 1691 -7129 1771 -7119
rect 1371 -7399 1431 -7129
rect 1701 -7139 1771 -7129
rect 1511 -7189 1541 -7169
rect 1491 -7229 1541 -7189
rect 1601 -7189 1631 -7169
rect 1601 -7229 1651 -7189
rect 1491 -7299 1651 -7229
rect 1491 -7339 1541 -7299
rect 1511 -7359 1541 -7339
rect 1601 -7339 1651 -7299
rect 1601 -7359 1631 -7339
rect 1711 -7399 1771 -7139
rect 1371 -7409 1451 -7399
rect 1371 -7469 1381 -7409
rect 1441 -7419 1451 -7409
rect 1691 -7409 1771 -7399
rect 1691 -7419 1701 -7409
rect 1441 -7469 1701 -7419
rect 1761 -7469 1771 -7409
rect 1371 -7479 1771 -7469
rect 1827 -7059 2227 -7049
rect 1827 -7119 1837 -7059
rect 1897 -7109 2157 -7059
rect 1897 -7119 1907 -7109
rect 1827 -7129 1907 -7119
rect 2147 -7119 2157 -7109
rect 2217 -7119 2227 -7059
rect 2147 -7129 2227 -7119
rect 1827 -7399 1887 -7129
rect 2157 -7139 2227 -7129
rect 1967 -7189 1997 -7169
rect 1947 -7229 1997 -7189
rect 2057 -7189 2087 -7169
rect 2057 -7229 2107 -7189
rect 1947 -7299 2107 -7229
rect 1947 -7339 1997 -7299
rect 1967 -7359 1997 -7339
rect 2057 -7339 2107 -7299
rect 2057 -7359 2087 -7339
rect 2167 -7399 2227 -7139
rect 1827 -7409 1907 -7399
rect 1827 -7469 1837 -7409
rect 1897 -7419 1907 -7409
rect 2147 -7409 2227 -7399
rect 2147 -7419 2157 -7409
rect 1897 -7469 2157 -7419
rect 2217 -7469 2227 -7409
rect 1827 -7479 2227 -7469
rect 2283 -7059 2683 -7049
rect 2283 -7119 2293 -7059
rect 2353 -7109 2613 -7059
rect 2353 -7119 2363 -7109
rect 2283 -7129 2363 -7119
rect 2603 -7119 2613 -7109
rect 2673 -7119 2683 -7059
rect 2603 -7129 2683 -7119
rect 2283 -7399 2343 -7129
rect 2613 -7139 2683 -7129
rect 2423 -7189 2453 -7169
rect 2403 -7229 2453 -7189
rect 2513 -7189 2543 -7169
rect 2513 -7229 2563 -7189
rect 2403 -7299 2563 -7229
rect 2403 -7339 2453 -7299
rect 2423 -7359 2453 -7339
rect 2513 -7339 2563 -7299
rect 2513 -7359 2543 -7339
rect 2623 -7399 2683 -7139
rect 2283 -7409 2363 -7399
rect 2283 -7469 2293 -7409
rect 2353 -7419 2363 -7409
rect 2603 -7409 2683 -7399
rect 2603 -7419 2613 -7409
rect 2353 -7469 2613 -7419
rect 2673 -7469 2683 -7409
rect 2283 -7479 2683 -7469
rect 2741 -7059 3141 -7049
rect 2741 -7119 2751 -7059
rect 2811 -7109 3071 -7059
rect 2811 -7119 2821 -7109
rect 2741 -7129 2821 -7119
rect 3061 -7119 3071 -7109
rect 3131 -7119 3141 -7059
rect 3061 -7129 3141 -7119
rect 2741 -7399 2801 -7129
rect 3071 -7139 3141 -7129
rect 2881 -7189 2911 -7169
rect 2861 -7229 2911 -7189
rect 2971 -7189 3001 -7169
rect 2971 -7229 3021 -7189
rect 2861 -7299 3021 -7229
rect 2861 -7339 2911 -7299
rect 2881 -7359 2911 -7339
rect 2971 -7339 3021 -7299
rect 2971 -7359 3001 -7339
rect 3081 -7399 3141 -7139
rect 2741 -7409 2821 -7399
rect 2741 -7469 2751 -7409
rect 2811 -7419 2821 -7409
rect 3061 -7409 3141 -7399
rect 3061 -7419 3071 -7409
rect 2811 -7469 3071 -7419
rect 3131 -7469 3141 -7409
rect 2741 -7479 3141 -7469
rect 3197 -7059 3597 -7049
rect 3197 -7119 3207 -7059
rect 3267 -7109 3527 -7059
rect 3267 -7119 3277 -7109
rect 3197 -7129 3277 -7119
rect 3517 -7119 3527 -7109
rect 3587 -7119 3597 -7059
rect 3517 -7129 3597 -7119
rect 3197 -7399 3257 -7129
rect 3527 -7139 3597 -7129
rect 3337 -7189 3367 -7169
rect 3317 -7229 3367 -7189
rect 3427 -7189 3457 -7169
rect 3427 -7229 3477 -7189
rect 3317 -7299 3477 -7229
rect 3317 -7339 3367 -7299
rect 3337 -7359 3367 -7339
rect 3427 -7339 3477 -7299
rect 3427 -7359 3457 -7339
rect 3537 -7399 3597 -7139
rect 3197 -7409 3277 -7399
rect 3197 -7469 3207 -7409
rect 3267 -7419 3277 -7409
rect 3517 -7409 3597 -7399
rect 3517 -7419 3527 -7409
rect 3267 -7469 3527 -7419
rect 3587 -7469 3597 -7409
rect 3197 -7479 3597 -7469
rect 3653 -7059 4053 -7049
rect 3653 -7119 3663 -7059
rect 3723 -7109 3983 -7059
rect 3723 -7119 3733 -7109
rect 3653 -7129 3733 -7119
rect 3973 -7119 3983 -7109
rect 4043 -7119 4053 -7059
rect 3973 -7129 4053 -7119
rect 3653 -7399 3713 -7129
rect 3983 -7139 4053 -7129
rect 3793 -7189 3823 -7169
rect 3773 -7229 3823 -7189
rect 3883 -7189 3913 -7169
rect 3883 -7229 3933 -7189
rect 3773 -7299 3933 -7229
rect 3773 -7339 3823 -7299
rect 3793 -7359 3823 -7339
rect 3883 -7339 3933 -7299
rect 3883 -7359 3913 -7339
rect 3993 -7399 4053 -7139
rect 3653 -7409 3733 -7399
rect 3653 -7469 3663 -7409
rect 3723 -7419 3733 -7409
rect 3973 -7409 4053 -7399
rect 3973 -7419 3983 -7409
rect 3723 -7469 3983 -7419
rect 4043 -7469 4053 -7409
rect 3653 -7479 4053 -7469
rect 4111 -7059 4511 -7049
rect 4111 -7119 4121 -7059
rect 4181 -7109 4441 -7059
rect 4181 -7119 4191 -7109
rect 4111 -7129 4191 -7119
rect 4431 -7119 4441 -7109
rect 4501 -7119 4511 -7059
rect 4431 -7129 4511 -7119
rect 4111 -7399 4171 -7129
rect 4441 -7139 4511 -7129
rect 4251 -7189 4281 -7169
rect 4231 -7229 4281 -7189
rect 4341 -7189 4371 -7169
rect 4341 -7229 4391 -7189
rect 4231 -7299 4391 -7229
rect 4231 -7339 4281 -7299
rect 4251 -7359 4281 -7339
rect 4341 -7339 4391 -7299
rect 4341 -7359 4371 -7339
rect 4451 -7399 4511 -7139
rect 4111 -7409 4191 -7399
rect 4111 -7469 4121 -7409
rect 4181 -7419 4191 -7409
rect 4431 -7409 4511 -7399
rect 4431 -7419 4441 -7409
rect 4181 -7469 4441 -7419
rect 4501 -7469 4511 -7409
rect 4111 -7479 4511 -7469
rect 4567 -7059 4967 -7049
rect 4567 -7119 4577 -7059
rect 4637 -7109 4897 -7059
rect 4637 -7119 4647 -7109
rect 4567 -7129 4647 -7119
rect 4887 -7119 4897 -7109
rect 4957 -7119 4967 -7059
rect 4887 -7129 4967 -7119
rect 4567 -7399 4627 -7129
rect 4897 -7139 4967 -7129
rect 4707 -7189 4737 -7169
rect 4687 -7229 4737 -7189
rect 4797 -7189 4827 -7169
rect 4797 -7229 4847 -7189
rect 4687 -7299 4847 -7229
rect 4687 -7339 4737 -7299
rect 4707 -7359 4737 -7339
rect 4797 -7339 4847 -7299
rect 4797 -7359 4827 -7339
rect 4907 -7399 4967 -7139
rect 4567 -7409 4647 -7399
rect 4567 -7469 4577 -7409
rect 4637 -7419 4647 -7409
rect 4887 -7409 4967 -7399
rect 4887 -7419 4897 -7409
rect 4637 -7469 4897 -7419
rect 4957 -7469 4967 -7409
rect 4567 -7479 4967 -7469
rect 5023 -7059 5423 -7049
rect 5023 -7119 5033 -7059
rect 5093 -7109 5353 -7059
rect 5093 -7119 5103 -7109
rect 5023 -7129 5103 -7119
rect 5343 -7119 5353 -7109
rect 5413 -7119 5423 -7059
rect 5343 -7129 5423 -7119
rect 5023 -7399 5083 -7129
rect 5353 -7139 5423 -7129
rect 5163 -7189 5193 -7169
rect 5143 -7229 5193 -7189
rect 5253 -7189 5283 -7169
rect 5253 -7229 5303 -7189
rect 5143 -7299 5303 -7229
rect 5143 -7339 5193 -7299
rect 5163 -7359 5193 -7339
rect 5253 -7339 5303 -7299
rect 5253 -7359 5283 -7339
rect 5363 -7399 5423 -7139
rect 5023 -7409 5103 -7399
rect 5023 -7469 5033 -7409
rect 5093 -7419 5103 -7409
rect 5343 -7409 5423 -7399
rect 5343 -7419 5353 -7409
rect 5093 -7469 5353 -7419
rect 5413 -7469 5423 -7409
rect 5023 -7479 5423 -7469
rect 5481 -7059 5881 -7049
rect 5481 -7119 5491 -7059
rect 5551 -7109 5811 -7059
rect 5551 -7119 5561 -7109
rect 5481 -7129 5561 -7119
rect 5801 -7119 5811 -7109
rect 5871 -7119 5881 -7059
rect 5801 -7129 5881 -7119
rect 5481 -7399 5541 -7129
rect 5811 -7139 5881 -7129
rect 5621 -7189 5651 -7169
rect 5601 -7229 5651 -7189
rect 5711 -7189 5741 -7169
rect 5711 -7229 5761 -7189
rect 5601 -7299 5761 -7229
rect 5601 -7339 5651 -7299
rect 5621 -7359 5651 -7339
rect 5711 -7339 5761 -7299
rect 5711 -7359 5741 -7339
rect 5821 -7399 5881 -7139
rect 5481 -7409 5561 -7399
rect 5481 -7469 5491 -7409
rect 5551 -7419 5561 -7409
rect 5801 -7409 5881 -7399
rect 5801 -7419 5811 -7409
rect 5551 -7469 5811 -7419
rect 5871 -7469 5881 -7409
rect 5481 -7479 5881 -7469
rect 5937 -7059 6337 -7049
rect 5937 -7119 5947 -7059
rect 6007 -7109 6267 -7059
rect 6007 -7119 6017 -7109
rect 5937 -7129 6017 -7119
rect 6257 -7119 6267 -7109
rect 6327 -7119 6337 -7059
rect 6257 -7129 6337 -7119
rect 5937 -7399 5997 -7129
rect 6267 -7139 6337 -7129
rect 6077 -7189 6107 -7169
rect 6057 -7229 6107 -7189
rect 6167 -7189 6197 -7169
rect 6167 -7229 6217 -7189
rect 6057 -7299 6217 -7229
rect 6057 -7339 6107 -7299
rect 6077 -7359 6107 -7339
rect 6167 -7339 6217 -7299
rect 6167 -7359 6197 -7339
rect 6277 -7399 6337 -7139
rect 5937 -7409 6017 -7399
rect 5937 -7469 5947 -7409
rect 6007 -7419 6017 -7409
rect 6257 -7409 6337 -7399
rect 6257 -7419 6267 -7409
rect 6007 -7469 6267 -7419
rect 6327 -7469 6337 -7409
rect 5937 -7479 6337 -7469
rect 6393 -7059 6793 -7049
rect 6393 -7119 6403 -7059
rect 6463 -7109 6723 -7059
rect 6463 -7119 6473 -7109
rect 6393 -7129 6473 -7119
rect 6713 -7119 6723 -7109
rect 6783 -7119 6793 -7059
rect 6713 -7129 6793 -7119
rect 6393 -7399 6453 -7129
rect 6723 -7139 6793 -7129
rect 6533 -7189 6563 -7169
rect 6513 -7229 6563 -7189
rect 6623 -7189 6653 -7169
rect 6623 -7229 6673 -7189
rect 6513 -7299 6673 -7229
rect 6513 -7339 6563 -7299
rect 6533 -7359 6563 -7339
rect 6623 -7339 6673 -7299
rect 6623 -7359 6653 -7339
rect 6733 -7399 6793 -7139
rect 6393 -7409 6473 -7399
rect 6393 -7469 6403 -7409
rect 6463 -7419 6473 -7409
rect 6713 -7409 6793 -7399
rect 6713 -7419 6723 -7409
rect 6463 -7469 6723 -7419
rect 6783 -7469 6793 -7409
rect 6393 -7479 6793 -7469
rect 6851 -7059 7251 -7049
rect 6851 -7119 6861 -7059
rect 6921 -7109 7181 -7059
rect 6921 -7119 6931 -7109
rect 6851 -7129 6931 -7119
rect 7171 -7119 7181 -7109
rect 7241 -7119 7251 -7059
rect 7171 -7129 7251 -7119
rect 6851 -7399 6911 -7129
rect 7181 -7139 7251 -7129
rect 6991 -7189 7021 -7169
rect 6971 -7229 7021 -7189
rect 7081 -7189 7111 -7169
rect 7081 -7229 7131 -7189
rect 6971 -7299 7131 -7229
rect 6971 -7339 7021 -7299
rect 6991 -7359 7021 -7339
rect 7081 -7339 7131 -7299
rect 7081 -7359 7111 -7339
rect 7191 -7399 7251 -7139
rect 6851 -7409 6931 -7399
rect 6851 -7469 6861 -7409
rect 6921 -7419 6931 -7409
rect 7171 -7409 7251 -7399
rect 7171 -7419 7181 -7409
rect 6921 -7469 7181 -7419
rect 7241 -7469 7251 -7409
rect 6851 -7479 7251 -7469
rect 7307 -7059 7707 -7049
rect 7307 -7119 7317 -7059
rect 7377 -7109 7637 -7059
rect 7377 -7119 7387 -7109
rect 7307 -7129 7387 -7119
rect 7627 -7119 7637 -7109
rect 7697 -7119 7707 -7059
rect 7627 -7129 7707 -7119
rect 7307 -7399 7367 -7129
rect 7637 -7139 7707 -7129
rect 7447 -7189 7477 -7169
rect 7427 -7229 7477 -7189
rect 7537 -7189 7567 -7169
rect 7537 -7229 7587 -7189
rect 7427 -7299 7587 -7229
rect 7427 -7339 7477 -7299
rect 7447 -7359 7477 -7339
rect 7537 -7339 7587 -7299
rect 7537 -7359 7567 -7339
rect 7647 -7399 7707 -7139
rect 7307 -7409 7387 -7399
rect 7307 -7469 7317 -7409
rect 7377 -7419 7387 -7409
rect 7627 -7409 7707 -7399
rect 7627 -7419 7637 -7409
rect 7377 -7469 7637 -7419
rect 7697 -7469 7707 -7409
rect 7307 -7479 7707 -7469
rect 7763 -7059 8163 -7049
rect 7763 -7119 7773 -7059
rect 7833 -7109 8093 -7059
rect 7833 -7119 7843 -7109
rect 7763 -7129 7843 -7119
rect 8083 -7119 8093 -7109
rect 8153 -7119 8163 -7059
rect 8083 -7129 8163 -7119
rect 7763 -7399 7823 -7129
rect 8093 -7139 8163 -7129
rect 7903 -7189 7933 -7169
rect 7883 -7229 7933 -7189
rect 7993 -7189 8023 -7169
rect 7993 -7229 8043 -7189
rect 7883 -7299 8043 -7229
rect 7883 -7339 7933 -7299
rect 7903 -7359 7933 -7339
rect 7993 -7339 8043 -7299
rect 7993 -7359 8023 -7339
rect 8103 -7399 8163 -7139
rect 7763 -7409 7843 -7399
rect 7763 -7469 7773 -7409
rect 7833 -7419 7843 -7409
rect 8083 -7409 8163 -7399
rect 8083 -7419 8093 -7409
rect 7833 -7469 8093 -7419
rect 8153 -7469 8163 -7409
rect 7763 -7479 8163 -7469
rect 8237 -7059 8637 -7049
rect 8237 -7119 8247 -7059
rect 8307 -7109 8567 -7059
rect 8307 -7119 8317 -7109
rect 8237 -7129 8317 -7119
rect 8557 -7119 8567 -7109
rect 8627 -7119 8637 -7059
rect 8557 -7129 8637 -7119
rect 8237 -7399 8297 -7129
rect 8567 -7139 8637 -7129
rect 8377 -7189 8407 -7169
rect 8357 -7229 8407 -7189
rect 8467 -7189 8497 -7169
rect 8467 -7229 8517 -7189
rect 8357 -7299 8517 -7229
rect 8357 -7339 8407 -7299
rect 8377 -7359 8407 -7339
rect 8467 -7339 8517 -7299
rect 8467 -7359 8497 -7339
rect 8577 -7399 8637 -7139
rect 8237 -7409 8317 -7399
rect 8237 -7469 8247 -7409
rect 8307 -7419 8317 -7409
rect 8557 -7409 8637 -7399
rect 8557 -7419 8567 -7409
rect 8307 -7469 8567 -7419
rect 8627 -7469 8637 -7409
rect 8237 -7479 8637 -7469
rect 8693 -7059 9093 -7049
rect 8693 -7119 8703 -7059
rect 8763 -7109 9023 -7059
rect 8763 -7119 8773 -7109
rect 8693 -7129 8773 -7119
rect 9013 -7119 9023 -7109
rect 9083 -7119 9093 -7059
rect 9013 -7129 9093 -7119
rect 8693 -7399 8753 -7129
rect 9023 -7139 9093 -7129
rect 8833 -7189 8863 -7169
rect 8813 -7229 8863 -7189
rect 8923 -7189 8953 -7169
rect 8923 -7229 8973 -7189
rect 8813 -7299 8973 -7229
rect 8813 -7339 8863 -7299
rect 8833 -7359 8863 -7339
rect 8923 -7339 8973 -7299
rect 8923 -7359 8953 -7339
rect 9033 -7399 9093 -7139
rect 8693 -7409 8773 -7399
rect 8693 -7469 8703 -7409
rect 8763 -7419 8773 -7409
rect 9013 -7409 9093 -7399
rect 9013 -7419 9023 -7409
rect 8763 -7469 9023 -7419
rect 9083 -7469 9093 -7409
rect 8693 -7479 9093 -7469
rect 9151 -7059 9551 -7049
rect 9151 -7119 9161 -7059
rect 9221 -7109 9481 -7059
rect 9221 -7119 9231 -7109
rect 9151 -7129 9231 -7119
rect 9471 -7119 9481 -7109
rect 9541 -7119 9551 -7059
rect 9471 -7129 9551 -7119
rect 9151 -7399 9211 -7129
rect 9481 -7139 9551 -7129
rect 9291 -7189 9321 -7169
rect 9271 -7229 9321 -7189
rect 9381 -7189 9411 -7169
rect 9381 -7229 9431 -7189
rect 9271 -7299 9431 -7229
rect 9271 -7339 9321 -7299
rect 9291 -7359 9321 -7339
rect 9381 -7339 9431 -7299
rect 9381 -7359 9411 -7339
rect 9491 -7399 9551 -7139
rect 9151 -7409 9231 -7399
rect 9151 -7469 9161 -7409
rect 9221 -7419 9231 -7409
rect 9471 -7409 9551 -7399
rect 9471 -7419 9481 -7409
rect 9221 -7469 9481 -7419
rect 9541 -7469 9551 -7409
rect 9151 -7479 9551 -7469
rect 9607 -7059 10007 -7049
rect 9607 -7119 9617 -7059
rect 9677 -7109 9937 -7059
rect 9677 -7119 9687 -7109
rect 9607 -7129 9687 -7119
rect 9927 -7119 9937 -7109
rect 9997 -7119 10007 -7059
rect 9927 -7129 10007 -7119
rect 9607 -7399 9667 -7129
rect 9937 -7139 10007 -7129
rect 9747 -7189 9777 -7169
rect 9727 -7229 9777 -7189
rect 9837 -7189 9867 -7169
rect 9837 -7229 9887 -7189
rect 9727 -7299 9887 -7229
rect 9727 -7339 9777 -7299
rect 9747 -7359 9777 -7339
rect 9837 -7339 9887 -7299
rect 9837 -7359 9867 -7339
rect 9947 -7399 10007 -7139
rect 9607 -7409 9687 -7399
rect 9607 -7469 9617 -7409
rect 9677 -7419 9687 -7409
rect 9927 -7409 10007 -7399
rect 9927 -7419 9937 -7409
rect 9677 -7469 9937 -7419
rect 9997 -7469 10007 -7409
rect 9607 -7479 10007 -7469
rect 10063 -7059 10463 -7049
rect 10063 -7119 10073 -7059
rect 10133 -7109 10393 -7059
rect 10133 -7119 10143 -7109
rect 10063 -7129 10143 -7119
rect 10383 -7119 10393 -7109
rect 10453 -7119 10463 -7059
rect 10383 -7129 10463 -7119
rect 10063 -7399 10123 -7129
rect 10393 -7139 10463 -7129
rect 10203 -7189 10233 -7169
rect 10183 -7229 10233 -7189
rect 10293 -7189 10323 -7169
rect 10293 -7229 10343 -7189
rect 10183 -7299 10343 -7229
rect 10183 -7339 10233 -7299
rect 10203 -7359 10233 -7339
rect 10293 -7339 10343 -7299
rect 10293 -7359 10323 -7339
rect 10403 -7399 10463 -7139
rect 10063 -7409 10143 -7399
rect 10063 -7469 10073 -7409
rect 10133 -7419 10143 -7409
rect 10383 -7409 10463 -7399
rect 10383 -7419 10393 -7409
rect 10133 -7469 10393 -7419
rect 10453 -7469 10463 -7409
rect 10063 -7479 10463 -7469
rect 10521 -7059 10921 -7049
rect 10521 -7119 10531 -7059
rect 10591 -7109 10851 -7059
rect 10591 -7119 10601 -7109
rect 10521 -7129 10601 -7119
rect 10841 -7119 10851 -7109
rect 10911 -7119 10921 -7059
rect 10841 -7129 10921 -7119
rect 10521 -7399 10581 -7129
rect 10851 -7139 10921 -7129
rect 10661 -7189 10691 -7169
rect 10641 -7229 10691 -7189
rect 10751 -7189 10781 -7169
rect 10751 -7229 10801 -7189
rect 10641 -7299 10801 -7229
rect 10641 -7339 10691 -7299
rect 10661 -7359 10691 -7339
rect 10751 -7339 10801 -7299
rect 10751 -7359 10781 -7339
rect 10861 -7399 10921 -7139
rect 10521 -7409 10601 -7399
rect 10521 -7469 10531 -7409
rect 10591 -7419 10601 -7409
rect 10841 -7409 10921 -7399
rect 10841 -7419 10851 -7409
rect 10591 -7469 10851 -7419
rect 10911 -7469 10921 -7409
rect 10521 -7479 10921 -7469
rect 10977 -7059 11377 -7049
rect 10977 -7119 10987 -7059
rect 11047 -7109 11307 -7059
rect 11047 -7119 11057 -7109
rect 10977 -7129 11057 -7119
rect 11297 -7119 11307 -7109
rect 11367 -7119 11377 -7059
rect 11297 -7129 11377 -7119
rect 10977 -7399 11037 -7129
rect 11307 -7139 11377 -7129
rect 11117 -7189 11147 -7169
rect 11097 -7229 11147 -7189
rect 11207 -7189 11237 -7169
rect 11207 -7229 11257 -7189
rect 11097 -7299 11257 -7229
rect 11097 -7339 11147 -7299
rect 11117 -7359 11147 -7339
rect 11207 -7339 11257 -7299
rect 11207 -7359 11237 -7339
rect 11317 -7399 11377 -7139
rect 10977 -7409 11057 -7399
rect 10977 -7469 10987 -7409
rect 11047 -7419 11057 -7409
rect 11297 -7409 11377 -7399
rect 11297 -7419 11307 -7409
rect 11047 -7469 11307 -7419
rect 11367 -7469 11377 -7409
rect 10977 -7479 11377 -7469
rect 11433 -7059 11833 -7049
rect 11433 -7119 11443 -7059
rect 11503 -7109 11763 -7059
rect 11503 -7119 11513 -7109
rect 11433 -7129 11513 -7119
rect 11753 -7119 11763 -7109
rect 11823 -7119 11833 -7059
rect 11753 -7129 11833 -7119
rect 11433 -7399 11493 -7129
rect 11763 -7139 11833 -7129
rect 11573 -7189 11603 -7169
rect 11553 -7229 11603 -7189
rect 11663 -7189 11693 -7169
rect 11663 -7229 11713 -7189
rect 11553 -7299 11713 -7229
rect 11553 -7339 11603 -7299
rect 11573 -7359 11603 -7339
rect 11663 -7339 11713 -7299
rect 11663 -7359 11693 -7339
rect 11773 -7399 11833 -7139
rect 11433 -7409 11513 -7399
rect 11433 -7469 11443 -7409
rect 11503 -7419 11513 -7409
rect 11753 -7409 11833 -7399
rect 11753 -7419 11763 -7409
rect 11503 -7469 11763 -7419
rect 11823 -7469 11833 -7409
rect 11433 -7479 11833 -7469
rect 11891 -7059 12291 -7049
rect 11891 -7119 11901 -7059
rect 11961 -7109 12221 -7059
rect 11961 -7119 11971 -7109
rect 11891 -7129 11971 -7119
rect 12211 -7119 12221 -7109
rect 12281 -7119 12291 -7059
rect 12211 -7129 12291 -7119
rect 11891 -7399 11951 -7129
rect 12221 -7139 12291 -7129
rect 12031 -7189 12061 -7169
rect 12011 -7229 12061 -7189
rect 12121 -7189 12151 -7169
rect 12121 -7229 12171 -7189
rect 12011 -7299 12171 -7229
rect 12011 -7339 12061 -7299
rect 12031 -7359 12061 -7339
rect 12121 -7339 12171 -7299
rect 12121 -7359 12151 -7339
rect 12231 -7399 12291 -7139
rect 11891 -7409 11971 -7399
rect 11891 -7469 11901 -7409
rect 11961 -7419 11971 -7409
rect 12211 -7409 12291 -7399
rect 12211 -7419 12221 -7409
rect 11961 -7469 12221 -7419
rect 12281 -7469 12291 -7409
rect 11891 -7479 12291 -7469
rect 12347 -7059 12747 -7049
rect 12347 -7119 12357 -7059
rect 12417 -7109 12677 -7059
rect 12417 -7119 12427 -7109
rect 12347 -7129 12427 -7119
rect 12667 -7119 12677 -7109
rect 12737 -7119 12747 -7059
rect 12667 -7129 12747 -7119
rect 12347 -7399 12407 -7129
rect 12677 -7139 12747 -7129
rect 12487 -7189 12517 -7169
rect 12467 -7229 12517 -7189
rect 12577 -7189 12607 -7169
rect 12577 -7229 12627 -7189
rect 12467 -7299 12627 -7229
rect 12467 -7339 12517 -7299
rect 12487 -7359 12517 -7339
rect 12577 -7339 12627 -7299
rect 12577 -7359 12607 -7339
rect 12687 -7399 12747 -7139
rect 12347 -7409 12427 -7399
rect 12347 -7469 12357 -7409
rect 12417 -7419 12427 -7409
rect 12667 -7409 12747 -7399
rect 12667 -7419 12677 -7409
rect 12417 -7469 12677 -7419
rect 12737 -7469 12747 -7409
rect 12347 -7479 12747 -7469
rect 12803 -7059 13203 -7049
rect 12803 -7119 12813 -7059
rect 12873 -7109 13133 -7059
rect 12873 -7119 12883 -7109
rect 12803 -7129 12883 -7119
rect 13123 -7119 13133 -7109
rect 13193 -7119 13203 -7059
rect 13123 -7129 13203 -7119
rect 12803 -7399 12863 -7129
rect 13133 -7139 13203 -7129
rect 12943 -7189 12973 -7169
rect 12923 -7229 12973 -7189
rect 13033 -7189 13063 -7169
rect 13033 -7229 13083 -7189
rect 12923 -7299 13083 -7229
rect 12923 -7339 12973 -7299
rect 12943 -7359 12973 -7339
rect 13033 -7339 13083 -7299
rect 13033 -7359 13063 -7339
rect 13143 -7399 13203 -7139
rect 12803 -7409 12883 -7399
rect 12803 -7469 12813 -7409
rect 12873 -7419 12883 -7409
rect 13123 -7409 13203 -7399
rect 13123 -7419 13133 -7409
rect 12873 -7469 13133 -7419
rect 13193 -7469 13203 -7409
rect 12803 -7479 13203 -7469
rect 13261 -7059 13661 -7049
rect 13261 -7119 13271 -7059
rect 13331 -7109 13591 -7059
rect 13331 -7119 13341 -7109
rect 13261 -7129 13341 -7119
rect 13581 -7119 13591 -7109
rect 13651 -7119 13661 -7059
rect 13581 -7129 13661 -7119
rect 13261 -7399 13321 -7129
rect 13591 -7139 13661 -7129
rect 13401 -7189 13431 -7169
rect 13381 -7229 13431 -7189
rect 13491 -7189 13521 -7169
rect 13491 -7229 13541 -7189
rect 13381 -7299 13541 -7229
rect 13381 -7339 13431 -7299
rect 13401 -7359 13431 -7339
rect 13491 -7339 13541 -7299
rect 13491 -7359 13521 -7339
rect 13601 -7399 13661 -7139
rect 13261 -7409 13341 -7399
rect 13261 -7469 13271 -7409
rect 13331 -7419 13341 -7409
rect 13581 -7409 13661 -7399
rect 13581 -7419 13591 -7409
rect 13331 -7469 13591 -7419
rect 13651 -7469 13661 -7409
rect 13261 -7479 13661 -7469
rect 13717 -7059 14117 -7049
rect 13717 -7119 13727 -7059
rect 13787 -7109 14047 -7059
rect 13787 -7119 13797 -7109
rect 13717 -7129 13797 -7119
rect 14037 -7119 14047 -7109
rect 14107 -7119 14117 -7059
rect 14037 -7129 14117 -7119
rect 13717 -7399 13777 -7129
rect 14047 -7139 14117 -7129
rect 13857 -7189 13887 -7169
rect 13837 -7229 13887 -7189
rect 13947 -7189 13977 -7169
rect 13947 -7229 13997 -7189
rect 13837 -7299 13997 -7229
rect 13837 -7339 13887 -7299
rect 13857 -7359 13887 -7339
rect 13947 -7339 13997 -7299
rect 13947 -7359 13977 -7339
rect 14057 -7399 14117 -7139
rect 13717 -7409 13797 -7399
rect 13717 -7469 13727 -7409
rect 13787 -7419 13797 -7409
rect 14037 -7409 14117 -7399
rect 14037 -7419 14047 -7409
rect 13787 -7469 14047 -7419
rect 14107 -7469 14117 -7409
rect 13717 -7479 14117 -7469
rect 14173 -7059 14573 -7049
rect 14173 -7119 14183 -7059
rect 14243 -7109 14503 -7059
rect 14243 -7119 14253 -7109
rect 14173 -7129 14253 -7119
rect 14493 -7119 14503 -7109
rect 14563 -7119 14573 -7059
rect 14493 -7129 14573 -7119
rect 14173 -7399 14233 -7129
rect 14503 -7139 14573 -7129
rect 14313 -7189 14343 -7169
rect 14293 -7229 14343 -7189
rect 14403 -7189 14433 -7169
rect 14403 -7229 14453 -7189
rect 14293 -7299 14453 -7229
rect 14293 -7339 14343 -7299
rect 14313 -7359 14343 -7339
rect 14403 -7339 14453 -7299
rect 14403 -7359 14433 -7339
rect 14513 -7399 14573 -7139
rect 14173 -7409 14253 -7399
rect 14173 -7469 14183 -7409
rect 14243 -7419 14253 -7409
rect 14493 -7409 14573 -7399
rect 14493 -7419 14503 -7409
rect 14243 -7469 14503 -7419
rect 14563 -7469 14573 -7409
rect 14173 -7479 14573 -7469
rect 14631 -7059 15031 -7049
rect 14631 -7119 14641 -7059
rect 14701 -7109 14961 -7059
rect 14701 -7119 14711 -7109
rect 14631 -7129 14711 -7119
rect 14951 -7119 14961 -7109
rect 15021 -7119 15031 -7059
rect 14951 -7129 15031 -7119
rect 14631 -7399 14691 -7129
rect 14961 -7139 15031 -7129
rect 14771 -7189 14801 -7169
rect 14751 -7229 14801 -7189
rect 14861 -7189 14891 -7169
rect 14861 -7229 14911 -7189
rect 14751 -7299 14911 -7229
rect 14751 -7339 14801 -7299
rect 14771 -7359 14801 -7339
rect 14861 -7339 14911 -7299
rect 14861 -7359 14891 -7339
rect 14971 -7399 15031 -7139
rect 14631 -7409 14711 -7399
rect 14631 -7469 14641 -7409
rect 14701 -7419 14711 -7409
rect 14951 -7409 15031 -7399
rect 14951 -7419 14961 -7409
rect 14701 -7469 14961 -7419
rect 15021 -7469 15031 -7409
rect 14631 -7479 15031 -7469
rect 15087 -7059 15487 -7049
rect 15087 -7119 15097 -7059
rect 15157 -7109 15417 -7059
rect 15157 -7119 15167 -7109
rect 15087 -7129 15167 -7119
rect 15407 -7119 15417 -7109
rect 15477 -7119 15487 -7059
rect 15407 -7129 15487 -7119
rect 15087 -7399 15147 -7129
rect 15417 -7139 15487 -7129
rect 15227 -7189 15257 -7169
rect 15207 -7229 15257 -7189
rect 15317 -7189 15347 -7169
rect 15317 -7229 15367 -7189
rect 15207 -7299 15367 -7229
rect 15207 -7339 15257 -7299
rect 15227 -7359 15257 -7339
rect 15317 -7339 15367 -7299
rect 15317 -7359 15347 -7339
rect 15427 -7399 15487 -7139
rect 15087 -7409 15167 -7399
rect 15087 -7469 15097 -7409
rect 15157 -7419 15167 -7409
rect 15407 -7409 15487 -7399
rect 15407 -7419 15417 -7409
rect 15157 -7469 15417 -7419
rect 15477 -7469 15487 -7409
rect 15087 -7479 15487 -7469
rect 1 -7561 401 -7551
rect 1 -7621 11 -7561
rect 71 -7611 331 -7561
rect 71 -7621 81 -7611
rect 1 -7631 81 -7621
rect 321 -7621 331 -7611
rect 391 -7621 401 -7561
rect 321 -7631 401 -7621
rect 1 -7901 61 -7631
rect 331 -7641 401 -7631
rect 141 -7691 171 -7671
rect 121 -7731 171 -7691
rect 231 -7691 261 -7671
rect 231 -7731 281 -7691
rect 121 -7801 281 -7731
rect 121 -7841 171 -7801
rect 141 -7861 171 -7841
rect 231 -7841 281 -7801
rect 231 -7861 261 -7841
rect 341 -7901 401 -7641
rect 1 -7911 81 -7901
rect 1 -7971 11 -7911
rect 71 -7921 81 -7911
rect 321 -7911 401 -7901
rect 321 -7921 331 -7911
rect 71 -7971 331 -7921
rect 391 -7971 401 -7911
rect 1 -7981 401 -7971
rect 457 -7561 857 -7551
rect 457 -7621 467 -7561
rect 527 -7611 787 -7561
rect 527 -7621 537 -7611
rect 457 -7631 537 -7621
rect 777 -7621 787 -7611
rect 847 -7621 857 -7561
rect 777 -7631 857 -7621
rect 457 -7901 517 -7631
rect 787 -7641 857 -7631
rect 597 -7691 627 -7671
rect 577 -7731 627 -7691
rect 687 -7691 717 -7671
rect 687 -7731 737 -7691
rect 577 -7801 737 -7731
rect 577 -7841 627 -7801
rect 597 -7861 627 -7841
rect 687 -7841 737 -7801
rect 687 -7861 717 -7841
rect 797 -7901 857 -7641
rect 457 -7911 537 -7901
rect 457 -7971 467 -7911
rect 527 -7921 537 -7911
rect 777 -7911 857 -7901
rect 777 -7921 787 -7911
rect 527 -7971 787 -7921
rect 847 -7971 857 -7911
rect 457 -7981 857 -7971
rect 913 -7561 1313 -7551
rect 913 -7621 923 -7561
rect 983 -7611 1243 -7561
rect 983 -7621 993 -7611
rect 913 -7631 993 -7621
rect 1233 -7621 1243 -7611
rect 1303 -7621 1313 -7561
rect 1233 -7631 1313 -7621
rect 913 -7901 973 -7631
rect 1243 -7641 1313 -7631
rect 1053 -7691 1083 -7671
rect 1033 -7731 1083 -7691
rect 1143 -7691 1173 -7671
rect 1143 -7731 1193 -7691
rect 1033 -7801 1193 -7731
rect 1033 -7841 1083 -7801
rect 1053 -7861 1083 -7841
rect 1143 -7841 1193 -7801
rect 1143 -7861 1173 -7841
rect 1253 -7901 1313 -7641
rect 913 -7911 993 -7901
rect 913 -7971 923 -7911
rect 983 -7921 993 -7911
rect 1233 -7911 1313 -7901
rect 1233 -7921 1243 -7911
rect 983 -7971 1243 -7921
rect 1303 -7971 1313 -7911
rect 913 -7981 1313 -7971
rect 1371 -7561 1771 -7551
rect 1371 -7621 1381 -7561
rect 1441 -7611 1701 -7561
rect 1441 -7621 1451 -7611
rect 1371 -7631 1451 -7621
rect 1691 -7621 1701 -7611
rect 1761 -7621 1771 -7561
rect 1691 -7631 1771 -7621
rect 1371 -7901 1431 -7631
rect 1701 -7641 1771 -7631
rect 1511 -7691 1541 -7671
rect 1491 -7731 1541 -7691
rect 1601 -7691 1631 -7671
rect 1601 -7731 1651 -7691
rect 1491 -7801 1651 -7731
rect 1491 -7841 1541 -7801
rect 1511 -7861 1541 -7841
rect 1601 -7841 1651 -7801
rect 1601 -7861 1631 -7841
rect 1711 -7901 1771 -7641
rect 1371 -7911 1451 -7901
rect 1371 -7971 1381 -7911
rect 1441 -7921 1451 -7911
rect 1691 -7911 1771 -7901
rect 1691 -7921 1701 -7911
rect 1441 -7971 1701 -7921
rect 1761 -7971 1771 -7911
rect 1371 -7981 1771 -7971
rect 1827 -7561 2227 -7551
rect 1827 -7621 1837 -7561
rect 1897 -7611 2157 -7561
rect 1897 -7621 1907 -7611
rect 1827 -7631 1907 -7621
rect 2147 -7621 2157 -7611
rect 2217 -7621 2227 -7561
rect 2147 -7631 2227 -7621
rect 1827 -7901 1887 -7631
rect 2157 -7641 2227 -7631
rect 1967 -7691 1997 -7671
rect 1947 -7731 1997 -7691
rect 2057 -7691 2087 -7671
rect 2057 -7731 2107 -7691
rect 1947 -7801 2107 -7731
rect 1947 -7841 1997 -7801
rect 1967 -7861 1997 -7841
rect 2057 -7841 2107 -7801
rect 2057 -7861 2087 -7841
rect 2167 -7901 2227 -7641
rect 1827 -7911 1907 -7901
rect 1827 -7971 1837 -7911
rect 1897 -7921 1907 -7911
rect 2147 -7911 2227 -7901
rect 2147 -7921 2157 -7911
rect 1897 -7971 2157 -7921
rect 2217 -7971 2227 -7911
rect 1827 -7981 2227 -7971
rect 2283 -7561 2683 -7551
rect 2283 -7621 2293 -7561
rect 2353 -7611 2613 -7561
rect 2353 -7621 2363 -7611
rect 2283 -7631 2363 -7621
rect 2603 -7621 2613 -7611
rect 2673 -7621 2683 -7561
rect 2603 -7631 2683 -7621
rect 2283 -7901 2343 -7631
rect 2613 -7641 2683 -7631
rect 2423 -7691 2453 -7671
rect 2403 -7731 2453 -7691
rect 2513 -7691 2543 -7671
rect 2513 -7731 2563 -7691
rect 2403 -7801 2563 -7731
rect 2403 -7841 2453 -7801
rect 2423 -7861 2453 -7841
rect 2513 -7841 2563 -7801
rect 2513 -7861 2543 -7841
rect 2623 -7901 2683 -7641
rect 2283 -7911 2363 -7901
rect 2283 -7971 2293 -7911
rect 2353 -7921 2363 -7911
rect 2603 -7911 2683 -7901
rect 2603 -7921 2613 -7911
rect 2353 -7971 2613 -7921
rect 2673 -7971 2683 -7911
rect 2283 -7981 2683 -7971
rect 2741 -7561 3141 -7551
rect 2741 -7621 2751 -7561
rect 2811 -7611 3071 -7561
rect 2811 -7621 2821 -7611
rect 2741 -7631 2821 -7621
rect 3061 -7621 3071 -7611
rect 3131 -7621 3141 -7561
rect 3061 -7631 3141 -7621
rect 2741 -7901 2801 -7631
rect 3071 -7641 3141 -7631
rect 2881 -7691 2911 -7671
rect 2861 -7731 2911 -7691
rect 2971 -7691 3001 -7671
rect 2971 -7731 3021 -7691
rect 2861 -7801 3021 -7731
rect 2861 -7841 2911 -7801
rect 2881 -7861 2911 -7841
rect 2971 -7841 3021 -7801
rect 2971 -7861 3001 -7841
rect 3081 -7901 3141 -7641
rect 2741 -7911 2821 -7901
rect 2741 -7971 2751 -7911
rect 2811 -7921 2821 -7911
rect 3061 -7911 3141 -7901
rect 3061 -7921 3071 -7911
rect 2811 -7971 3071 -7921
rect 3131 -7971 3141 -7911
rect 2741 -7981 3141 -7971
rect 3197 -7561 3597 -7551
rect 3197 -7621 3207 -7561
rect 3267 -7611 3527 -7561
rect 3267 -7621 3277 -7611
rect 3197 -7631 3277 -7621
rect 3517 -7621 3527 -7611
rect 3587 -7621 3597 -7561
rect 3517 -7631 3597 -7621
rect 3197 -7901 3257 -7631
rect 3527 -7641 3597 -7631
rect 3337 -7691 3367 -7671
rect 3317 -7731 3367 -7691
rect 3427 -7691 3457 -7671
rect 3427 -7731 3477 -7691
rect 3317 -7801 3477 -7731
rect 3317 -7841 3367 -7801
rect 3337 -7861 3367 -7841
rect 3427 -7841 3477 -7801
rect 3427 -7861 3457 -7841
rect 3537 -7901 3597 -7641
rect 3197 -7911 3277 -7901
rect 3197 -7971 3207 -7911
rect 3267 -7921 3277 -7911
rect 3517 -7911 3597 -7901
rect 3517 -7921 3527 -7911
rect 3267 -7971 3527 -7921
rect 3587 -7971 3597 -7911
rect 3197 -7981 3597 -7971
rect 3653 -7561 4053 -7551
rect 3653 -7621 3663 -7561
rect 3723 -7611 3983 -7561
rect 3723 -7621 3733 -7611
rect 3653 -7631 3733 -7621
rect 3973 -7621 3983 -7611
rect 4043 -7621 4053 -7561
rect 3973 -7631 4053 -7621
rect 3653 -7901 3713 -7631
rect 3983 -7641 4053 -7631
rect 3793 -7691 3823 -7671
rect 3773 -7731 3823 -7691
rect 3883 -7691 3913 -7671
rect 3883 -7731 3933 -7691
rect 3773 -7801 3933 -7731
rect 3773 -7841 3823 -7801
rect 3793 -7861 3823 -7841
rect 3883 -7841 3933 -7801
rect 3883 -7861 3913 -7841
rect 3993 -7901 4053 -7641
rect 3653 -7911 3733 -7901
rect 3653 -7971 3663 -7911
rect 3723 -7921 3733 -7911
rect 3973 -7911 4053 -7901
rect 3973 -7921 3983 -7911
rect 3723 -7971 3983 -7921
rect 4043 -7971 4053 -7911
rect 3653 -7981 4053 -7971
rect 4111 -7561 4511 -7551
rect 4111 -7621 4121 -7561
rect 4181 -7611 4441 -7561
rect 4181 -7621 4191 -7611
rect 4111 -7631 4191 -7621
rect 4431 -7621 4441 -7611
rect 4501 -7621 4511 -7561
rect 4431 -7631 4511 -7621
rect 4111 -7901 4171 -7631
rect 4441 -7641 4511 -7631
rect 4251 -7691 4281 -7671
rect 4231 -7731 4281 -7691
rect 4341 -7691 4371 -7671
rect 4341 -7731 4391 -7691
rect 4231 -7801 4391 -7731
rect 4231 -7841 4281 -7801
rect 4251 -7861 4281 -7841
rect 4341 -7841 4391 -7801
rect 4341 -7861 4371 -7841
rect 4451 -7901 4511 -7641
rect 4111 -7911 4191 -7901
rect 4111 -7971 4121 -7911
rect 4181 -7921 4191 -7911
rect 4431 -7911 4511 -7901
rect 4431 -7921 4441 -7911
rect 4181 -7971 4441 -7921
rect 4501 -7971 4511 -7911
rect 4111 -7981 4511 -7971
rect 4567 -7561 4967 -7551
rect 4567 -7621 4577 -7561
rect 4637 -7611 4897 -7561
rect 4637 -7621 4647 -7611
rect 4567 -7631 4647 -7621
rect 4887 -7621 4897 -7611
rect 4957 -7621 4967 -7561
rect 4887 -7631 4967 -7621
rect 4567 -7901 4627 -7631
rect 4897 -7641 4967 -7631
rect 4707 -7691 4737 -7671
rect 4687 -7731 4737 -7691
rect 4797 -7691 4827 -7671
rect 4797 -7731 4847 -7691
rect 4687 -7801 4847 -7731
rect 4687 -7841 4737 -7801
rect 4707 -7861 4737 -7841
rect 4797 -7841 4847 -7801
rect 4797 -7861 4827 -7841
rect 4907 -7901 4967 -7641
rect 4567 -7911 4647 -7901
rect 4567 -7971 4577 -7911
rect 4637 -7921 4647 -7911
rect 4887 -7911 4967 -7901
rect 4887 -7921 4897 -7911
rect 4637 -7971 4897 -7921
rect 4957 -7971 4967 -7911
rect 4567 -7981 4967 -7971
rect 5023 -7561 5423 -7551
rect 5023 -7621 5033 -7561
rect 5093 -7611 5353 -7561
rect 5093 -7621 5103 -7611
rect 5023 -7631 5103 -7621
rect 5343 -7621 5353 -7611
rect 5413 -7621 5423 -7561
rect 5343 -7631 5423 -7621
rect 5023 -7901 5083 -7631
rect 5353 -7641 5423 -7631
rect 5163 -7691 5193 -7671
rect 5143 -7731 5193 -7691
rect 5253 -7691 5283 -7671
rect 5253 -7731 5303 -7691
rect 5143 -7801 5303 -7731
rect 5143 -7841 5193 -7801
rect 5163 -7861 5193 -7841
rect 5253 -7841 5303 -7801
rect 5253 -7861 5283 -7841
rect 5363 -7901 5423 -7641
rect 5023 -7911 5103 -7901
rect 5023 -7971 5033 -7911
rect 5093 -7921 5103 -7911
rect 5343 -7911 5423 -7901
rect 5343 -7921 5353 -7911
rect 5093 -7971 5353 -7921
rect 5413 -7971 5423 -7911
rect 5023 -7981 5423 -7971
rect 5481 -7561 5881 -7551
rect 5481 -7621 5491 -7561
rect 5551 -7611 5811 -7561
rect 5551 -7621 5561 -7611
rect 5481 -7631 5561 -7621
rect 5801 -7621 5811 -7611
rect 5871 -7621 5881 -7561
rect 5801 -7631 5881 -7621
rect 5481 -7901 5541 -7631
rect 5811 -7641 5881 -7631
rect 5621 -7691 5651 -7671
rect 5601 -7731 5651 -7691
rect 5711 -7691 5741 -7671
rect 5711 -7731 5761 -7691
rect 5601 -7801 5761 -7731
rect 5601 -7841 5651 -7801
rect 5621 -7861 5651 -7841
rect 5711 -7841 5761 -7801
rect 5711 -7861 5741 -7841
rect 5821 -7901 5881 -7641
rect 5481 -7911 5561 -7901
rect 5481 -7971 5491 -7911
rect 5551 -7921 5561 -7911
rect 5801 -7911 5881 -7901
rect 5801 -7921 5811 -7911
rect 5551 -7971 5811 -7921
rect 5871 -7971 5881 -7911
rect 5481 -7981 5881 -7971
rect 5937 -7561 6337 -7551
rect 5937 -7621 5947 -7561
rect 6007 -7611 6267 -7561
rect 6007 -7621 6017 -7611
rect 5937 -7631 6017 -7621
rect 6257 -7621 6267 -7611
rect 6327 -7621 6337 -7561
rect 6257 -7631 6337 -7621
rect 5937 -7901 5997 -7631
rect 6267 -7641 6337 -7631
rect 6077 -7691 6107 -7671
rect 6057 -7731 6107 -7691
rect 6167 -7691 6197 -7671
rect 6167 -7731 6217 -7691
rect 6057 -7801 6217 -7731
rect 6057 -7841 6107 -7801
rect 6077 -7861 6107 -7841
rect 6167 -7841 6217 -7801
rect 6167 -7861 6197 -7841
rect 6277 -7901 6337 -7641
rect 5937 -7911 6017 -7901
rect 5937 -7971 5947 -7911
rect 6007 -7921 6017 -7911
rect 6257 -7911 6337 -7901
rect 6257 -7921 6267 -7911
rect 6007 -7971 6267 -7921
rect 6327 -7971 6337 -7911
rect 5937 -7981 6337 -7971
rect 6393 -7561 6793 -7551
rect 6393 -7621 6403 -7561
rect 6463 -7611 6723 -7561
rect 6463 -7621 6473 -7611
rect 6393 -7631 6473 -7621
rect 6713 -7621 6723 -7611
rect 6783 -7621 6793 -7561
rect 6713 -7631 6793 -7621
rect 6393 -7901 6453 -7631
rect 6723 -7641 6793 -7631
rect 6533 -7691 6563 -7671
rect 6513 -7731 6563 -7691
rect 6623 -7691 6653 -7671
rect 6623 -7731 6673 -7691
rect 6513 -7801 6673 -7731
rect 6513 -7841 6563 -7801
rect 6533 -7861 6563 -7841
rect 6623 -7841 6673 -7801
rect 6623 -7861 6653 -7841
rect 6733 -7901 6793 -7641
rect 6393 -7911 6473 -7901
rect 6393 -7971 6403 -7911
rect 6463 -7921 6473 -7911
rect 6713 -7911 6793 -7901
rect 6713 -7921 6723 -7911
rect 6463 -7971 6723 -7921
rect 6783 -7971 6793 -7911
rect 6393 -7981 6793 -7971
rect 6851 -7561 7251 -7551
rect 6851 -7621 6861 -7561
rect 6921 -7611 7181 -7561
rect 6921 -7621 6931 -7611
rect 6851 -7631 6931 -7621
rect 7171 -7621 7181 -7611
rect 7241 -7621 7251 -7561
rect 7171 -7631 7251 -7621
rect 6851 -7901 6911 -7631
rect 7181 -7641 7251 -7631
rect 6991 -7691 7021 -7671
rect 6971 -7731 7021 -7691
rect 7081 -7691 7111 -7671
rect 7081 -7731 7131 -7691
rect 6971 -7801 7131 -7731
rect 6971 -7841 7021 -7801
rect 6991 -7861 7021 -7841
rect 7081 -7841 7131 -7801
rect 7081 -7861 7111 -7841
rect 7191 -7901 7251 -7641
rect 6851 -7911 6931 -7901
rect 6851 -7971 6861 -7911
rect 6921 -7921 6931 -7911
rect 7171 -7911 7251 -7901
rect 7171 -7921 7181 -7911
rect 6921 -7971 7181 -7921
rect 7241 -7971 7251 -7911
rect 6851 -7981 7251 -7971
rect 7307 -7561 7707 -7551
rect 7307 -7621 7317 -7561
rect 7377 -7611 7637 -7561
rect 7377 -7621 7387 -7611
rect 7307 -7631 7387 -7621
rect 7627 -7621 7637 -7611
rect 7697 -7621 7707 -7561
rect 7627 -7631 7707 -7621
rect 7307 -7901 7367 -7631
rect 7637 -7641 7707 -7631
rect 7447 -7691 7477 -7671
rect 7427 -7731 7477 -7691
rect 7537 -7691 7567 -7671
rect 7537 -7731 7587 -7691
rect 7427 -7801 7587 -7731
rect 7427 -7841 7477 -7801
rect 7447 -7861 7477 -7841
rect 7537 -7841 7587 -7801
rect 7537 -7861 7567 -7841
rect 7647 -7901 7707 -7641
rect 7307 -7911 7387 -7901
rect 7307 -7971 7317 -7911
rect 7377 -7921 7387 -7911
rect 7627 -7911 7707 -7901
rect 7627 -7921 7637 -7911
rect 7377 -7971 7637 -7921
rect 7697 -7971 7707 -7911
rect 7307 -7981 7707 -7971
rect 7763 -7561 8163 -7551
rect 7763 -7621 7773 -7561
rect 7833 -7611 8093 -7561
rect 7833 -7621 7843 -7611
rect 7763 -7631 7843 -7621
rect 8083 -7621 8093 -7611
rect 8153 -7621 8163 -7561
rect 8083 -7631 8163 -7621
rect 7763 -7901 7823 -7631
rect 8093 -7641 8163 -7631
rect 7903 -7691 7933 -7671
rect 7883 -7731 7933 -7691
rect 7993 -7691 8023 -7671
rect 7993 -7731 8043 -7691
rect 7883 -7801 8043 -7731
rect 7883 -7841 7933 -7801
rect 7903 -7861 7933 -7841
rect 7993 -7841 8043 -7801
rect 7993 -7861 8023 -7841
rect 8103 -7901 8163 -7641
rect 7763 -7911 7843 -7901
rect 7763 -7971 7773 -7911
rect 7833 -7921 7843 -7911
rect 8083 -7911 8163 -7901
rect 8083 -7921 8093 -7911
rect 7833 -7971 8093 -7921
rect 8153 -7971 8163 -7911
rect 7763 -7981 8163 -7971
rect 8237 -7561 8637 -7551
rect 8237 -7621 8247 -7561
rect 8307 -7611 8567 -7561
rect 8307 -7621 8317 -7611
rect 8237 -7631 8317 -7621
rect 8557 -7621 8567 -7611
rect 8627 -7621 8637 -7561
rect 8557 -7631 8637 -7621
rect 8237 -7901 8297 -7631
rect 8567 -7641 8637 -7631
rect 8377 -7691 8407 -7671
rect 8357 -7731 8407 -7691
rect 8467 -7691 8497 -7671
rect 8467 -7731 8517 -7691
rect 8357 -7801 8517 -7731
rect 8357 -7841 8407 -7801
rect 8377 -7861 8407 -7841
rect 8467 -7841 8517 -7801
rect 8467 -7861 8497 -7841
rect 8577 -7901 8637 -7641
rect 8237 -7911 8317 -7901
rect 8237 -7971 8247 -7911
rect 8307 -7921 8317 -7911
rect 8557 -7911 8637 -7901
rect 8557 -7921 8567 -7911
rect 8307 -7971 8567 -7921
rect 8627 -7971 8637 -7911
rect 8237 -7981 8637 -7971
rect 8693 -7561 9093 -7551
rect 8693 -7621 8703 -7561
rect 8763 -7611 9023 -7561
rect 8763 -7621 8773 -7611
rect 8693 -7631 8773 -7621
rect 9013 -7621 9023 -7611
rect 9083 -7621 9093 -7561
rect 9013 -7631 9093 -7621
rect 8693 -7901 8753 -7631
rect 9023 -7641 9093 -7631
rect 8833 -7691 8863 -7671
rect 8813 -7731 8863 -7691
rect 8923 -7691 8953 -7671
rect 8923 -7731 8973 -7691
rect 8813 -7801 8973 -7731
rect 8813 -7841 8863 -7801
rect 8833 -7861 8863 -7841
rect 8923 -7841 8973 -7801
rect 8923 -7861 8953 -7841
rect 9033 -7901 9093 -7641
rect 8693 -7911 8773 -7901
rect 8693 -7971 8703 -7911
rect 8763 -7921 8773 -7911
rect 9013 -7911 9093 -7901
rect 9013 -7921 9023 -7911
rect 8763 -7971 9023 -7921
rect 9083 -7971 9093 -7911
rect 8693 -7981 9093 -7971
rect 9151 -7561 9551 -7551
rect 9151 -7621 9161 -7561
rect 9221 -7611 9481 -7561
rect 9221 -7621 9231 -7611
rect 9151 -7631 9231 -7621
rect 9471 -7621 9481 -7611
rect 9541 -7621 9551 -7561
rect 9471 -7631 9551 -7621
rect 9151 -7901 9211 -7631
rect 9481 -7641 9551 -7631
rect 9291 -7691 9321 -7671
rect 9271 -7731 9321 -7691
rect 9381 -7691 9411 -7671
rect 9381 -7731 9431 -7691
rect 9271 -7801 9431 -7731
rect 9271 -7841 9321 -7801
rect 9291 -7861 9321 -7841
rect 9381 -7841 9431 -7801
rect 9381 -7861 9411 -7841
rect 9491 -7901 9551 -7641
rect 9151 -7911 9231 -7901
rect 9151 -7971 9161 -7911
rect 9221 -7921 9231 -7911
rect 9471 -7911 9551 -7901
rect 9471 -7921 9481 -7911
rect 9221 -7971 9481 -7921
rect 9541 -7971 9551 -7911
rect 9151 -7981 9551 -7971
rect 9607 -7561 10007 -7551
rect 9607 -7621 9617 -7561
rect 9677 -7611 9937 -7561
rect 9677 -7621 9687 -7611
rect 9607 -7631 9687 -7621
rect 9927 -7621 9937 -7611
rect 9997 -7621 10007 -7561
rect 9927 -7631 10007 -7621
rect 9607 -7901 9667 -7631
rect 9937 -7641 10007 -7631
rect 9747 -7691 9777 -7671
rect 9727 -7731 9777 -7691
rect 9837 -7691 9867 -7671
rect 9837 -7731 9887 -7691
rect 9727 -7801 9887 -7731
rect 9727 -7841 9777 -7801
rect 9747 -7861 9777 -7841
rect 9837 -7841 9887 -7801
rect 9837 -7861 9867 -7841
rect 9947 -7901 10007 -7641
rect 9607 -7911 9687 -7901
rect 9607 -7971 9617 -7911
rect 9677 -7921 9687 -7911
rect 9927 -7911 10007 -7901
rect 9927 -7921 9937 -7911
rect 9677 -7971 9937 -7921
rect 9997 -7971 10007 -7911
rect 9607 -7981 10007 -7971
rect 10063 -7561 10463 -7551
rect 10063 -7621 10073 -7561
rect 10133 -7611 10393 -7561
rect 10133 -7621 10143 -7611
rect 10063 -7631 10143 -7621
rect 10383 -7621 10393 -7611
rect 10453 -7621 10463 -7561
rect 10383 -7631 10463 -7621
rect 10063 -7901 10123 -7631
rect 10393 -7641 10463 -7631
rect 10203 -7691 10233 -7671
rect 10183 -7731 10233 -7691
rect 10293 -7691 10323 -7671
rect 10293 -7731 10343 -7691
rect 10183 -7801 10343 -7731
rect 10183 -7841 10233 -7801
rect 10203 -7861 10233 -7841
rect 10293 -7841 10343 -7801
rect 10293 -7861 10323 -7841
rect 10403 -7901 10463 -7641
rect 10063 -7911 10143 -7901
rect 10063 -7971 10073 -7911
rect 10133 -7921 10143 -7911
rect 10383 -7911 10463 -7901
rect 10383 -7921 10393 -7911
rect 10133 -7971 10393 -7921
rect 10453 -7971 10463 -7911
rect 10063 -7981 10463 -7971
rect 10521 -7561 10921 -7551
rect 10521 -7621 10531 -7561
rect 10591 -7611 10851 -7561
rect 10591 -7621 10601 -7611
rect 10521 -7631 10601 -7621
rect 10841 -7621 10851 -7611
rect 10911 -7621 10921 -7561
rect 10841 -7631 10921 -7621
rect 10521 -7901 10581 -7631
rect 10851 -7641 10921 -7631
rect 10661 -7691 10691 -7671
rect 10641 -7731 10691 -7691
rect 10751 -7691 10781 -7671
rect 10751 -7731 10801 -7691
rect 10641 -7801 10801 -7731
rect 10641 -7841 10691 -7801
rect 10661 -7861 10691 -7841
rect 10751 -7841 10801 -7801
rect 10751 -7861 10781 -7841
rect 10861 -7901 10921 -7641
rect 10521 -7911 10601 -7901
rect 10521 -7971 10531 -7911
rect 10591 -7921 10601 -7911
rect 10841 -7911 10921 -7901
rect 10841 -7921 10851 -7911
rect 10591 -7971 10851 -7921
rect 10911 -7971 10921 -7911
rect 10521 -7981 10921 -7971
rect 10977 -7561 11377 -7551
rect 10977 -7621 10987 -7561
rect 11047 -7611 11307 -7561
rect 11047 -7621 11057 -7611
rect 10977 -7631 11057 -7621
rect 11297 -7621 11307 -7611
rect 11367 -7621 11377 -7561
rect 11297 -7631 11377 -7621
rect 10977 -7901 11037 -7631
rect 11307 -7641 11377 -7631
rect 11117 -7691 11147 -7671
rect 11097 -7731 11147 -7691
rect 11207 -7691 11237 -7671
rect 11207 -7731 11257 -7691
rect 11097 -7801 11257 -7731
rect 11097 -7841 11147 -7801
rect 11117 -7861 11147 -7841
rect 11207 -7841 11257 -7801
rect 11207 -7861 11237 -7841
rect 11317 -7901 11377 -7641
rect 10977 -7911 11057 -7901
rect 10977 -7971 10987 -7911
rect 11047 -7921 11057 -7911
rect 11297 -7911 11377 -7901
rect 11297 -7921 11307 -7911
rect 11047 -7971 11307 -7921
rect 11367 -7971 11377 -7911
rect 10977 -7981 11377 -7971
rect 11433 -7561 11833 -7551
rect 11433 -7621 11443 -7561
rect 11503 -7611 11763 -7561
rect 11503 -7621 11513 -7611
rect 11433 -7631 11513 -7621
rect 11753 -7621 11763 -7611
rect 11823 -7621 11833 -7561
rect 11753 -7631 11833 -7621
rect 11433 -7901 11493 -7631
rect 11763 -7641 11833 -7631
rect 11573 -7691 11603 -7671
rect 11553 -7731 11603 -7691
rect 11663 -7691 11693 -7671
rect 11663 -7731 11713 -7691
rect 11553 -7801 11713 -7731
rect 11553 -7841 11603 -7801
rect 11573 -7861 11603 -7841
rect 11663 -7841 11713 -7801
rect 11663 -7861 11693 -7841
rect 11773 -7901 11833 -7641
rect 11433 -7911 11513 -7901
rect 11433 -7971 11443 -7911
rect 11503 -7921 11513 -7911
rect 11753 -7911 11833 -7901
rect 11753 -7921 11763 -7911
rect 11503 -7971 11763 -7921
rect 11823 -7971 11833 -7911
rect 11433 -7981 11833 -7971
rect 11891 -7561 12291 -7551
rect 11891 -7621 11901 -7561
rect 11961 -7611 12221 -7561
rect 11961 -7621 11971 -7611
rect 11891 -7631 11971 -7621
rect 12211 -7621 12221 -7611
rect 12281 -7621 12291 -7561
rect 12211 -7631 12291 -7621
rect 11891 -7901 11951 -7631
rect 12221 -7641 12291 -7631
rect 12031 -7691 12061 -7671
rect 12011 -7731 12061 -7691
rect 12121 -7691 12151 -7671
rect 12121 -7731 12171 -7691
rect 12011 -7801 12171 -7731
rect 12011 -7841 12061 -7801
rect 12031 -7861 12061 -7841
rect 12121 -7841 12171 -7801
rect 12121 -7861 12151 -7841
rect 12231 -7901 12291 -7641
rect 11891 -7911 11971 -7901
rect 11891 -7971 11901 -7911
rect 11961 -7921 11971 -7911
rect 12211 -7911 12291 -7901
rect 12211 -7921 12221 -7911
rect 11961 -7971 12221 -7921
rect 12281 -7971 12291 -7911
rect 11891 -7981 12291 -7971
rect 12347 -7561 12747 -7551
rect 12347 -7621 12357 -7561
rect 12417 -7611 12677 -7561
rect 12417 -7621 12427 -7611
rect 12347 -7631 12427 -7621
rect 12667 -7621 12677 -7611
rect 12737 -7621 12747 -7561
rect 12667 -7631 12747 -7621
rect 12347 -7901 12407 -7631
rect 12677 -7641 12747 -7631
rect 12487 -7691 12517 -7671
rect 12467 -7731 12517 -7691
rect 12577 -7691 12607 -7671
rect 12577 -7731 12627 -7691
rect 12467 -7801 12627 -7731
rect 12467 -7841 12517 -7801
rect 12487 -7861 12517 -7841
rect 12577 -7841 12627 -7801
rect 12577 -7861 12607 -7841
rect 12687 -7901 12747 -7641
rect 12347 -7911 12427 -7901
rect 12347 -7971 12357 -7911
rect 12417 -7921 12427 -7911
rect 12667 -7911 12747 -7901
rect 12667 -7921 12677 -7911
rect 12417 -7971 12677 -7921
rect 12737 -7971 12747 -7911
rect 12347 -7981 12747 -7971
rect 12803 -7561 13203 -7551
rect 12803 -7621 12813 -7561
rect 12873 -7611 13133 -7561
rect 12873 -7621 12883 -7611
rect 12803 -7631 12883 -7621
rect 13123 -7621 13133 -7611
rect 13193 -7621 13203 -7561
rect 13123 -7631 13203 -7621
rect 12803 -7901 12863 -7631
rect 13133 -7641 13203 -7631
rect 12943 -7691 12973 -7671
rect 12923 -7731 12973 -7691
rect 13033 -7691 13063 -7671
rect 13033 -7731 13083 -7691
rect 12923 -7801 13083 -7731
rect 12923 -7841 12973 -7801
rect 12943 -7861 12973 -7841
rect 13033 -7841 13083 -7801
rect 13033 -7861 13063 -7841
rect 13143 -7901 13203 -7641
rect 12803 -7911 12883 -7901
rect 12803 -7971 12813 -7911
rect 12873 -7921 12883 -7911
rect 13123 -7911 13203 -7901
rect 13123 -7921 13133 -7911
rect 12873 -7971 13133 -7921
rect 13193 -7971 13203 -7911
rect 12803 -7981 13203 -7971
rect 13261 -7561 13661 -7551
rect 13261 -7621 13271 -7561
rect 13331 -7611 13591 -7561
rect 13331 -7621 13341 -7611
rect 13261 -7631 13341 -7621
rect 13581 -7621 13591 -7611
rect 13651 -7621 13661 -7561
rect 13581 -7631 13661 -7621
rect 13261 -7901 13321 -7631
rect 13591 -7641 13661 -7631
rect 13401 -7691 13431 -7671
rect 13381 -7731 13431 -7691
rect 13491 -7691 13521 -7671
rect 13491 -7731 13541 -7691
rect 13381 -7801 13541 -7731
rect 13381 -7841 13431 -7801
rect 13401 -7861 13431 -7841
rect 13491 -7841 13541 -7801
rect 13491 -7861 13521 -7841
rect 13601 -7901 13661 -7641
rect 13261 -7911 13341 -7901
rect 13261 -7971 13271 -7911
rect 13331 -7921 13341 -7911
rect 13581 -7911 13661 -7901
rect 13581 -7921 13591 -7911
rect 13331 -7971 13591 -7921
rect 13651 -7971 13661 -7911
rect 13261 -7981 13661 -7971
rect 13717 -7561 14117 -7551
rect 13717 -7621 13727 -7561
rect 13787 -7611 14047 -7561
rect 13787 -7621 13797 -7611
rect 13717 -7631 13797 -7621
rect 14037 -7621 14047 -7611
rect 14107 -7621 14117 -7561
rect 14037 -7631 14117 -7621
rect 13717 -7901 13777 -7631
rect 14047 -7641 14117 -7631
rect 13857 -7691 13887 -7671
rect 13837 -7731 13887 -7691
rect 13947 -7691 13977 -7671
rect 13947 -7731 13997 -7691
rect 13837 -7801 13997 -7731
rect 13837 -7841 13887 -7801
rect 13857 -7861 13887 -7841
rect 13947 -7841 13997 -7801
rect 13947 -7861 13977 -7841
rect 14057 -7901 14117 -7641
rect 13717 -7911 13797 -7901
rect 13717 -7971 13727 -7911
rect 13787 -7921 13797 -7911
rect 14037 -7911 14117 -7901
rect 14037 -7921 14047 -7911
rect 13787 -7971 14047 -7921
rect 14107 -7971 14117 -7911
rect 13717 -7981 14117 -7971
rect 14173 -7561 14573 -7551
rect 14173 -7621 14183 -7561
rect 14243 -7611 14503 -7561
rect 14243 -7621 14253 -7611
rect 14173 -7631 14253 -7621
rect 14493 -7621 14503 -7611
rect 14563 -7621 14573 -7561
rect 14493 -7631 14573 -7621
rect 14173 -7901 14233 -7631
rect 14503 -7641 14573 -7631
rect 14313 -7691 14343 -7671
rect 14293 -7731 14343 -7691
rect 14403 -7691 14433 -7671
rect 14403 -7731 14453 -7691
rect 14293 -7801 14453 -7731
rect 14293 -7841 14343 -7801
rect 14313 -7861 14343 -7841
rect 14403 -7841 14453 -7801
rect 14403 -7861 14433 -7841
rect 14513 -7901 14573 -7641
rect 14173 -7911 14253 -7901
rect 14173 -7971 14183 -7911
rect 14243 -7921 14253 -7911
rect 14493 -7911 14573 -7901
rect 14493 -7921 14503 -7911
rect 14243 -7971 14503 -7921
rect 14563 -7971 14573 -7911
rect 14173 -7981 14573 -7971
rect 14631 -7561 15031 -7551
rect 14631 -7621 14641 -7561
rect 14701 -7611 14961 -7561
rect 14701 -7621 14711 -7611
rect 14631 -7631 14711 -7621
rect 14951 -7621 14961 -7611
rect 15021 -7621 15031 -7561
rect 14951 -7631 15031 -7621
rect 14631 -7901 14691 -7631
rect 14961 -7641 15031 -7631
rect 14771 -7691 14801 -7671
rect 14751 -7731 14801 -7691
rect 14861 -7691 14891 -7671
rect 14861 -7731 14911 -7691
rect 14751 -7801 14911 -7731
rect 14751 -7841 14801 -7801
rect 14771 -7861 14801 -7841
rect 14861 -7841 14911 -7801
rect 14861 -7861 14891 -7841
rect 14971 -7901 15031 -7641
rect 14631 -7911 14711 -7901
rect 14631 -7971 14641 -7911
rect 14701 -7921 14711 -7911
rect 14951 -7911 15031 -7901
rect 14951 -7921 14961 -7911
rect 14701 -7971 14961 -7921
rect 15021 -7971 15031 -7911
rect 14631 -7981 15031 -7971
rect 15087 -7561 15487 -7551
rect 15087 -7621 15097 -7561
rect 15157 -7611 15417 -7561
rect 15157 -7621 15167 -7611
rect 15087 -7631 15167 -7621
rect 15407 -7621 15417 -7611
rect 15477 -7621 15487 -7561
rect 15407 -7631 15487 -7621
rect 15087 -7901 15147 -7631
rect 15417 -7641 15487 -7631
rect 15227 -7691 15257 -7671
rect 15207 -7731 15257 -7691
rect 15317 -7691 15347 -7671
rect 15317 -7731 15367 -7691
rect 15207 -7801 15367 -7731
rect 15207 -7841 15257 -7801
rect 15227 -7861 15257 -7841
rect 15317 -7841 15367 -7801
rect 15317 -7861 15347 -7841
rect 15427 -7901 15487 -7641
rect 15087 -7911 15167 -7901
rect 15087 -7971 15097 -7911
rect 15157 -7921 15167 -7911
rect 15407 -7911 15487 -7901
rect 15407 -7921 15417 -7911
rect 15157 -7971 15417 -7921
rect 15477 -7971 15487 -7911
rect 15087 -7981 15487 -7971
rect 1 -8053 401 -8043
rect 1 -8113 11 -8053
rect 71 -8103 331 -8053
rect 71 -8113 81 -8103
rect 1 -8123 81 -8113
rect 321 -8113 331 -8103
rect 391 -8113 401 -8053
rect 321 -8123 401 -8113
rect 1 -8393 61 -8123
rect 331 -8133 401 -8123
rect 141 -8183 171 -8163
rect 121 -8223 171 -8183
rect 231 -8183 261 -8163
rect 231 -8223 281 -8183
rect 121 -8293 281 -8223
rect 121 -8333 171 -8293
rect 141 -8353 171 -8333
rect 231 -8333 281 -8293
rect 231 -8353 261 -8333
rect 341 -8393 401 -8133
rect 1 -8403 81 -8393
rect 1 -8463 11 -8403
rect 71 -8413 81 -8403
rect 321 -8403 401 -8393
rect 321 -8413 331 -8403
rect 71 -8463 331 -8413
rect 391 -8463 401 -8403
rect 1 -8473 401 -8463
rect 457 -8053 857 -8043
rect 457 -8113 467 -8053
rect 527 -8103 787 -8053
rect 527 -8113 537 -8103
rect 457 -8123 537 -8113
rect 777 -8113 787 -8103
rect 847 -8113 857 -8053
rect 777 -8123 857 -8113
rect 457 -8393 517 -8123
rect 787 -8133 857 -8123
rect 597 -8183 627 -8163
rect 577 -8223 627 -8183
rect 687 -8183 717 -8163
rect 687 -8223 737 -8183
rect 577 -8293 737 -8223
rect 577 -8333 627 -8293
rect 597 -8353 627 -8333
rect 687 -8333 737 -8293
rect 687 -8353 717 -8333
rect 797 -8393 857 -8133
rect 457 -8403 537 -8393
rect 457 -8463 467 -8403
rect 527 -8413 537 -8403
rect 777 -8403 857 -8393
rect 777 -8413 787 -8403
rect 527 -8463 787 -8413
rect 847 -8463 857 -8403
rect 457 -8473 857 -8463
rect 913 -8053 1313 -8043
rect 913 -8113 923 -8053
rect 983 -8103 1243 -8053
rect 983 -8113 993 -8103
rect 913 -8123 993 -8113
rect 1233 -8113 1243 -8103
rect 1303 -8113 1313 -8053
rect 1233 -8123 1313 -8113
rect 913 -8393 973 -8123
rect 1243 -8133 1313 -8123
rect 1053 -8183 1083 -8163
rect 1033 -8223 1083 -8183
rect 1143 -8183 1173 -8163
rect 1143 -8223 1193 -8183
rect 1033 -8293 1193 -8223
rect 1033 -8333 1083 -8293
rect 1053 -8353 1083 -8333
rect 1143 -8333 1193 -8293
rect 1143 -8353 1173 -8333
rect 1253 -8393 1313 -8133
rect 913 -8403 993 -8393
rect 913 -8463 923 -8403
rect 983 -8413 993 -8403
rect 1233 -8403 1313 -8393
rect 1233 -8413 1243 -8403
rect 983 -8463 1243 -8413
rect 1303 -8463 1313 -8403
rect 913 -8473 1313 -8463
rect 1371 -8053 1771 -8043
rect 1371 -8113 1381 -8053
rect 1441 -8103 1701 -8053
rect 1441 -8113 1451 -8103
rect 1371 -8123 1451 -8113
rect 1691 -8113 1701 -8103
rect 1761 -8113 1771 -8053
rect 1691 -8123 1771 -8113
rect 1371 -8393 1431 -8123
rect 1701 -8133 1771 -8123
rect 1511 -8183 1541 -8163
rect 1491 -8223 1541 -8183
rect 1601 -8183 1631 -8163
rect 1601 -8223 1651 -8183
rect 1491 -8293 1651 -8223
rect 1491 -8333 1541 -8293
rect 1511 -8353 1541 -8333
rect 1601 -8333 1651 -8293
rect 1601 -8353 1631 -8333
rect 1711 -8393 1771 -8133
rect 1371 -8403 1451 -8393
rect 1371 -8463 1381 -8403
rect 1441 -8413 1451 -8403
rect 1691 -8403 1771 -8393
rect 1691 -8413 1701 -8403
rect 1441 -8463 1701 -8413
rect 1761 -8463 1771 -8403
rect 1371 -8473 1771 -8463
rect 1827 -8053 2227 -8043
rect 1827 -8113 1837 -8053
rect 1897 -8103 2157 -8053
rect 1897 -8113 1907 -8103
rect 1827 -8123 1907 -8113
rect 2147 -8113 2157 -8103
rect 2217 -8113 2227 -8053
rect 2147 -8123 2227 -8113
rect 1827 -8393 1887 -8123
rect 2157 -8133 2227 -8123
rect 1967 -8183 1997 -8163
rect 1947 -8223 1997 -8183
rect 2057 -8183 2087 -8163
rect 2057 -8223 2107 -8183
rect 1947 -8293 2107 -8223
rect 1947 -8333 1997 -8293
rect 1967 -8353 1997 -8333
rect 2057 -8333 2107 -8293
rect 2057 -8353 2087 -8333
rect 2167 -8393 2227 -8133
rect 1827 -8403 1907 -8393
rect 1827 -8463 1837 -8403
rect 1897 -8413 1907 -8403
rect 2147 -8403 2227 -8393
rect 2147 -8413 2157 -8403
rect 1897 -8463 2157 -8413
rect 2217 -8463 2227 -8403
rect 1827 -8473 2227 -8463
rect 2283 -8053 2683 -8043
rect 2283 -8113 2293 -8053
rect 2353 -8103 2613 -8053
rect 2353 -8113 2363 -8103
rect 2283 -8123 2363 -8113
rect 2603 -8113 2613 -8103
rect 2673 -8113 2683 -8053
rect 2603 -8123 2683 -8113
rect 2283 -8393 2343 -8123
rect 2613 -8133 2683 -8123
rect 2423 -8183 2453 -8163
rect 2403 -8223 2453 -8183
rect 2513 -8183 2543 -8163
rect 2513 -8223 2563 -8183
rect 2403 -8293 2563 -8223
rect 2403 -8333 2453 -8293
rect 2423 -8353 2453 -8333
rect 2513 -8333 2563 -8293
rect 2513 -8353 2543 -8333
rect 2623 -8393 2683 -8133
rect 2283 -8403 2363 -8393
rect 2283 -8463 2293 -8403
rect 2353 -8413 2363 -8403
rect 2603 -8403 2683 -8393
rect 2603 -8413 2613 -8403
rect 2353 -8463 2613 -8413
rect 2673 -8463 2683 -8403
rect 2283 -8473 2683 -8463
rect 2741 -8053 3141 -8043
rect 2741 -8113 2751 -8053
rect 2811 -8103 3071 -8053
rect 2811 -8113 2821 -8103
rect 2741 -8123 2821 -8113
rect 3061 -8113 3071 -8103
rect 3131 -8113 3141 -8053
rect 3061 -8123 3141 -8113
rect 2741 -8393 2801 -8123
rect 3071 -8133 3141 -8123
rect 2881 -8183 2911 -8163
rect 2861 -8223 2911 -8183
rect 2971 -8183 3001 -8163
rect 2971 -8223 3021 -8183
rect 2861 -8293 3021 -8223
rect 2861 -8333 2911 -8293
rect 2881 -8353 2911 -8333
rect 2971 -8333 3021 -8293
rect 2971 -8353 3001 -8333
rect 3081 -8393 3141 -8133
rect 2741 -8403 2821 -8393
rect 2741 -8463 2751 -8403
rect 2811 -8413 2821 -8403
rect 3061 -8403 3141 -8393
rect 3061 -8413 3071 -8403
rect 2811 -8463 3071 -8413
rect 3131 -8463 3141 -8403
rect 2741 -8473 3141 -8463
rect 3197 -8053 3597 -8043
rect 3197 -8113 3207 -8053
rect 3267 -8103 3527 -8053
rect 3267 -8113 3277 -8103
rect 3197 -8123 3277 -8113
rect 3517 -8113 3527 -8103
rect 3587 -8113 3597 -8053
rect 3517 -8123 3597 -8113
rect 3197 -8393 3257 -8123
rect 3527 -8133 3597 -8123
rect 3337 -8183 3367 -8163
rect 3317 -8223 3367 -8183
rect 3427 -8183 3457 -8163
rect 3427 -8223 3477 -8183
rect 3317 -8293 3477 -8223
rect 3317 -8333 3367 -8293
rect 3337 -8353 3367 -8333
rect 3427 -8333 3477 -8293
rect 3427 -8353 3457 -8333
rect 3537 -8393 3597 -8133
rect 3197 -8403 3277 -8393
rect 3197 -8463 3207 -8403
rect 3267 -8413 3277 -8403
rect 3517 -8403 3597 -8393
rect 3517 -8413 3527 -8403
rect 3267 -8463 3527 -8413
rect 3587 -8463 3597 -8403
rect 3197 -8473 3597 -8463
rect 3653 -8053 4053 -8043
rect 3653 -8113 3663 -8053
rect 3723 -8103 3983 -8053
rect 3723 -8113 3733 -8103
rect 3653 -8123 3733 -8113
rect 3973 -8113 3983 -8103
rect 4043 -8113 4053 -8053
rect 3973 -8123 4053 -8113
rect 3653 -8393 3713 -8123
rect 3983 -8133 4053 -8123
rect 3793 -8183 3823 -8163
rect 3773 -8223 3823 -8183
rect 3883 -8183 3913 -8163
rect 3883 -8223 3933 -8183
rect 3773 -8293 3933 -8223
rect 3773 -8333 3823 -8293
rect 3793 -8353 3823 -8333
rect 3883 -8333 3933 -8293
rect 3883 -8353 3913 -8333
rect 3993 -8393 4053 -8133
rect 3653 -8403 3733 -8393
rect 3653 -8463 3663 -8403
rect 3723 -8413 3733 -8403
rect 3973 -8403 4053 -8393
rect 3973 -8413 3983 -8403
rect 3723 -8463 3983 -8413
rect 4043 -8463 4053 -8403
rect 3653 -8473 4053 -8463
rect 4111 -8053 4511 -8043
rect 4111 -8113 4121 -8053
rect 4181 -8103 4441 -8053
rect 4181 -8113 4191 -8103
rect 4111 -8123 4191 -8113
rect 4431 -8113 4441 -8103
rect 4501 -8113 4511 -8053
rect 4431 -8123 4511 -8113
rect 4111 -8393 4171 -8123
rect 4441 -8133 4511 -8123
rect 4251 -8183 4281 -8163
rect 4231 -8223 4281 -8183
rect 4341 -8183 4371 -8163
rect 4341 -8223 4391 -8183
rect 4231 -8293 4391 -8223
rect 4231 -8333 4281 -8293
rect 4251 -8353 4281 -8333
rect 4341 -8333 4391 -8293
rect 4341 -8353 4371 -8333
rect 4451 -8393 4511 -8133
rect 4111 -8403 4191 -8393
rect 4111 -8463 4121 -8403
rect 4181 -8413 4191 -8403
rect 4431 -8403 4511 -8393
rect 4431 -8413 4441 -8403
rect 4181 -8463 4441 -8413
rect 4501 -8463 4511 -8403
rect 4111 -8473 4511 -8463
rect 4567 -8053 4967 -8043
rect 4567 -8113 4577 -8053
rect 4637 -8103 4897 -8053
rect 4637 -8113 4647 -8103
rect 4567 -8123 4647 -8113
rect 4887 -8113 4897 -8103
rect 4957 -8113 4967 -8053
rect 4887 -8123 4967 -8113
rect 4567 -8393 4627 -8123
rect 4897 -8133 4967 -8123
rect 4707 -8183 4737 -8163
rect 4687 -8223 4737 -8183
rect 4797 -8183 4827 -8163
rect 4797 -8223 4847 -8183
rect 4687 -8293 4847 -8223
rect 4687 -8333 4737 -8293
rect 4707 -8353 4737 -8333
rect 4797 -8333 4847 -8293
rect 4797 -8353 4827 -8333
rect 4907 -8393 4967 -8133
rect 4567 -8403 4647 -8393
rect 4567 -8463 4577 -8403
rect 4637 -8413 4647 -8403
rect 4887 -8403 4967 -8393
rect 4887 -8413 4897 -8403
rect 4637 -8463 4897 -8413
rect 4957 -8463 4967 -8403
rect 4567 -8473 4967 -8463
rect 5023 -8053 5423 -8043
rect 5023 -8113 5033 -8053
rect 5093 -8103 5353 -8053
rect 5093 -8113 5103 -8103
rect 5023 -8123 5103 -8113
rect 5343 -8113 5353 -8103
rect 5413 -8113 5423 -8053
rect 5343 -8123 5423 -8113
rect 5023 -8393 5083 -8123
rect 5353 -8133 5423 -8123
rect 5163 -8183 5193 -8163
rect 5143 -8223 5193 -8183
rect 5253 -8183 5283 -8163
rect 5253 -8223 5303 -8183
rect 5143 -8293 5303 -8223
rect 5143 -8333 5193 -8293
rect 5163 -8353 5193 -8333
rect 5253 -8333 5303 -8293
rect 5253 -8353 5283 -8333
rect 5363 -8393 5423 -8133
rect 5023 -8403 5103 -8393
rect 5023 -8463 5033 -8403
rect 5093 -8413 5103 -8403
rect 5343 -8403 5423 -8393
rect 5343 -8413 5353 -8403
rect 5093 -8463 5353 -8413
rect 5413 -8463 5423 -8403
rect 5023 -8473 5423 -8463
rect 5481 -8053 5881 -8043
rect 5481 -8113 5491 -8053
rect 5551 -8103 5811 -8053
rect 5551 -8113 5561 -8103
rect 5481 -8123 5561 -8113
rect 5801 -8113 5811 -8103
rect 5871 -8113 5881 -8053
rect 5801 -8123 5881 -8113
rect 5481 -8393 5541 -8123
rect 5811 -8133 5881 -8123
rect 5621 -8183 5651 -8163
rect 5601 -8223 5651 -8183
rect 5711 -8183 5741 -8163
rect 5711 -8223 5761 -8183
rect 5601 -8293 5761 -8223
rect 5601 -8333 5651 -8293
rect 5621 -8353 5651 -8333
rect 5711 -8333 5761 -8293
rect 5711 -8353 5741 -8333
rect 5821 -8393 5881 -8133
rect 5481 -8403 5561 -8393
rect 5481 -8463 5491 -8403
rect 5551 -8413 5561 -8403
rect 5801 -8403 5881 -8393
rect 5801 -8413 5811 -8403
rect 5551 -8463 5811 -8413
rect 5871 -8463 5881 -8403
rect 5481 -8473 5881 -8463
rect 5937 -8053 6337 -8043
rect 5937 -8113 5947 -8053
rect 6007 -8103 6267 -8053
rect 6007 -8113 6017 -8103
rect 5937 -8123 6017 -8113
rect 6257 -8113 6267 -8103
rect 6327 -8113 6337 -8053
rect 6257 -8123 6337 -8113
rect 5937 -8393 5997 -8123
rect 6267 -8133 6337 -8123
rect 6077 -8183 6107 -8163
rect 6057 -8223 6107 -8183
rect 6167 -8183 6197 -8163
rect 6167 -8223 6217 -8183
rect 6057 -8293 6217 -8223
rect 6057 -8333 6107 -8293
rect 6077 -8353 6107 -8333
rect 6167 -8333 6217 -8293
rect 6167 -8353 6197 -8333
rect 6277 -8393 6337 -8133
rect 5937 -8403 6017 -8393
rect 5937 -8463 5947 -8403
rect 6007 -8413 6017 -8403
rect 6257 -8403 6337 -8393
rect 6257 -8413 6267 -8403
rect 6007 -8463 6267 -8413
rect 6327 -8463 6337 -8403
rect 5937 -8473 6337 -8463
rect 6393 -8053 6793 -8043
rect 6393 -8113 6403 -8053
rect 6463 -8103 6723 -8053
rect 6463 -8113 6473 -8103
rect 6393 -8123 6473 -8113
rect 6713 -8113 6723 -8103
rect 6783 -8113 6793 -8053
rect 6713 -8123 6793 -8113
rect 6393 -8393 6453 -8123
rect 6723 -8133 6793 -8123
rect 6533 -8183 6563 -8163
rect 6513 -8223 6563 -8183
rect 6623 -8183 6653 -8163
rect 6623 -8223 6673 -8183
rect 6513 -8293 6673 -8223
rect 6513 -8333 6563 -8293
rect 6533 -8353 6563 -8333
rect 6623 -8333 6673 -8293
rect 6623 -8353 6653 -8333
rect 6733 -8393 6793 -8133
rect 6393 -8403 6473 -8393
rect 6393 -8463 6403 -8403
rect 6463 -8413 6473 -8403
rect 6713 -8403 6793 -8393
rect 6713 -8413 6723 -8403
rect 6463 -8463 6723 -8413
rect 6783 -8463 6793 -8403
rect 6393 -8473 6793 -8463
rect 6851 -8053 7251 -8043
rect 6851 -8113 6861 -8053
rect 6921 -8103 7181 -8053
rect 6921 -8113 6931 -8103
rect 6851 -8123 6931 -8113
rect 7171 -8113 7181 -8103
rect 7241 -8113 7251 -8053
rect 7171 -8123 7251 -8113
rect 6851 -8393 6911 -8123
rect 7181 -8133 7251 -8123
rect 6991 -8183 7021 -8163
rect 6971 -8223 7021 -8183
rect 7081 -8183 7111 -8163
rect 7081 -8223 7131 -8183
rect 6971 -8293 7131 -8223
rect 6971 -8333 7021 -8293
rect 6991 -8353 7021 -8333
rect 7081 -8333 7131 -8293
rect 7081 -8353 7111 -8333
rect 7191 -8393 7251 -8133
rect 6851 -8403 6931 -8393
rect 6851 -8463 6861 -8403
rect 6921 -8413 6931 -8403
rect 7171 -8403 7251 -8393
rect 7171 -8413 7181 -8403
rect 6921 -8463 7181 -8413
rect 7241 -8463 7251 -8403
rect 6851 -8473 7251 -8463
rect 7307 -8053 7707 -8043
rect 7307 -8113 7317 -8053
rect 7377 -8103 7637 -8053
rect 7377 -8113 7387 -8103
rect 7307 -8123 7387 -8113
rect 7627 -8113 7637 -8103
rect 7697 -8113 7707 -8053
rect 7627 -8123 7707 -8113
rect 7307 -8393 7367 -8123
rect 7637 -8133 7707 -8123
rect 7447 -8183 7477 -8163
rect 7427 -8223 7477 -8183
rect 7537 -8183 7567 -8163
rect 7537 -8223 7587 -8183
rect 7427 -8293 7587 -8223
rect 7427 -8333 7477 -8293
rect 7447 -8353 7477 -8333
rect 7537 -8333 7587 -8293
rect 7537 -8353 7567 -8333
rect 7647 -8393 7707 -8133
rect 7307 -8403 7387 -8393
rect 7307 -8463 7317 -8403
rect 7377 -8413 7387 -8403
rect 7627 -8403 7707 -8393
rect 7627 -8413 7637 -8403
rect 7377 -8463 7637 -8413
rect 7697 -8463 7707 -8403
rect 7307 -8473 7707 -8463
rect 7763 -8053 8163 -8043
rect 7763 -8113 7773 -8053
rect 7833 -8103 8093 -8053
rect 7833 -8113 7843 -8103
rect 7763 -8123 7843 -8113
rect 8083 -8113 8093 -8103
rect 8153 -8113 8163 -8053
rect 8083 -8123 8163 -8113
rect 7763 -8393 7823 -8123
rect 8093 -8133 8163 -8123
rect 7903 -8183 7933 -8163
rect 7883 -8223 7933 -8183
rect 7993 -8183 8023 -8163
rect 7993 -8223 8043 -8183
rect 7883 -8293 8043 -8223
rect 7883 -8333 7933 -8293
rect 7903 -8353 7933 -8333
rect 7993 -8333 8043 -8293
rect 7993 -8353 8023 -8333
rect 8103 -8393 8163 -8133
rect 7763 -8403 7843 -8393
rect 7763 -8463 7773 -8403
rect 7833 -8413 7843 -8403
rect 8083 -8403 8163 -8393
rect 8083 -8413 8093 -8403
rect 7833 -8463 8093 -8413
rect 8153 -8463 8163 -8403
rect 7763 -8473 8163 -8463
rect 8237 -8053 8637 -8043
rect 8237 -8113 8247 -8053
rect 8307 -8103 8567 -8053
rect 8307 -8113 8317 -8103
rect 8237 -8123 8317 -8113
rect 8557 -8113 8567 -8103
rect 8627 -8113 8637 -8053
rect 8557 -8123 8637 -8113
rect 8237 -8393 8297 -8123
rect 8567 -8133 8637 -8123
rect 8377 -8183 8407 -8163
rect 8357 -8223 8407 -8183
rect 8467 -8183 8497 -8163
rect 8467 -8223 8517 -8183
rect 8357 -8293 8517 -8223
rect 8357 -8333 8407 -8293
rect 8377 -8353 8407 -8333
rect 8467 -8333 8517 -8293
rect 8467 -8353 8497 -8333
rect 8577 -8393 8637 -8133
rect 8237 -8403 8317 -8393
rect 8237 -8463 8247 -8403
rect 8307 -8413 8317 -8403
rect 8557 -8403 8637 -8393
rect 8557 -8413 8567 -8403
rect 8307 -8463 8567 -8413
rect 8627 -8463 8637 -8403
rect 8237 -8473 8637 -8463
rect 8693 -8053 9093 -8043
rect 8693 -8113 8703 -8053
rect 8763 -8103 9023 -8053
rect 8763 -8113 8773 -8103
rect 8693 -8123 8773 -8113
rect 9013 -8113 9023 -8103
rect 9083 -8113 9093 -8053
rect 9013 -8123 9093 -8113
rect 8693 -8393 8753 -8123
rect 9023 -8133 9093 -8123
rect 8833 -8183 8863 -8163
rect 8813 -8223 8863 -8183
rect 8923 -8183 8953 -8163
rect 8923 -8223 8973 -8183
rect 8813 -8293 8973 -8223
rect 8813 -8333 8863 -8293
rect 8833 -8353 8863 -8333
rect 8923 -8333 8973 -8293
rect 8923 -8353 8953 -8333
rect 9033 -8393 9093 -8133
rect 8693 -8403 8773 -8393
rect 8693 -8463 8703 -8403
rect 8763 -8413 8773 -8403
rect 9013 -8403 9093 -8393
rect 9013 -8413 9023 -8403
rect 8763 -8463 9023 -8413
rect 9083 -8463 9093 -8403
rect 8693 -8473 9093 -8463
rect 9151 -8053 9551 -8043
rect 9151 -8113 9161 -8053
rect 9221 -8103 9481 -8053
rect 9221 -8113 9231 -8103
rect 9151 -8123 9231 -8113
rect 9471 -8113 9481 -8103
rect 9541 -8113 9551 -8053
rect 9471 -8123 9551 -8113
rect 9151 -8393 9211 -8123
rect 9481 -8133 9551 -8123
rect 9291 -8183 9321 -8163
rect 9271 -8223 9321 -8183
rect 9381 -8183 9411 -8163
rect 9381 -8223 9431 -8183
rect 9271 -8293 9431 -8223
rect 9271 -8333 9321 -8293
rect 9291 -8353 9321 -8333
rect 9381 -8333 9431 -8293
rect 9381 -8353 9411 -8333
rect 9491 -8393 9551 -8133
rect 9151 -8403 9231 -8393
rect 9151 -8463 9161 -8403
rect 9221 -8413 9231 -8403
rect 9471 -8403 9551 -8393
rect 9471 -8413 9481 -8403
rect 9221 -8463 9481 -8413
rect 9541 -8463 9551 -8403
rect 9151 -8473 9551 -8463
rect 9607 -8053 10007 -8043
rect 9607 -8113 9617 -8053
rect 9677 -8103 9937 -8053
rect 9677 -8113 9687 -8103
rect 9607 -8123 9687 -8113
rect 9927 -8113 9937 -8103
rect 9997 -8113 10007 -8053
rect 9927 -8123 10007 -8113
rect 9607 -8393 9667 -8123
rect 9937 -8133 10007 -8123
rect 9747 -8183 9777 -8163
rect 9727 -8223 9777 -8183
rect 9837 -8183 9867 -8163
rect 9837 -8223 9887 -8183
rect 9727 -8293 9887 -8223
rect 9727 -8333 9777 -8293
rect 9747 -8353 9777 -8333
rect 9837 -8333 9887 -8293
rect 9837 -8353 9867 -8333
rect 9947 -8393 10007 -8133
rect 9607 -8403 9687 -8393
rect 9607 -8463 9617 -8403
rect 9677 -8413 9687 -8403
rect 9927 -8403 10007 -8393
rect 9927 -8413 9937 -8403
rect 9677 -8463 9937 -8413
rect 9997 -8463 10007 -8403
rect 9607 -8473 10007 -8463
rect 10063 -8053 10463 -8043
rect 10063 -8113 10073 -8053
rect 10133 -8103 10393 -8053
rect 10133 -8113 10143 -8103
rect 10063 -8123 10143 -8113
rect 10383 -8113 10393 -8103
rect 10453 -8113 10463 -8053
rect 10383 -8123 10463 -8113
rect 10063 -8393 10123 -8123
rect 10393 -8133 10463 -8123
rect 10203 -8183 10233 -8163
rect 10183 -8223 10233 -8183
rect 10293 -8183 10323 -8163
rect 10293 -8223 10343 -8183
rect 10183 -8293 10343 -8223
rect 10183 -8333 10233 -8293
rect 10203 -8353 10233 -8333
rect 10293 -8333 10343 -8293
rect 10293 -8353 10323 -8333
rect 10403 -8393 10463 -8133
rect 10063 -8403 10143 -8393
rect 10063 -8463 10073 -8403
rect 10133 -8413 10143 -8403
rect 10383 -8403 10463 -8393
rect 10383 -8413 10393 -8403
rect 10133 -8463 10393 -8413
rect 10453 -8463 10463 -8403
rect 10063 -8473 10463 -8463
rect 10521 -8053 10921 -8043
rect 10521 -8113 10531 -8053
rect 10591 -8103 10851 -8053
rect 10591 -8113 10601 -8103
rect 10521 -8123 10601 -8113
rect 10841 -8113 10851 -8103
rect 10911 -8113 10921 -8053
rect 10841 -8123 10921 -8113
rect 10521 -8393 10581 -8123
rect 10851 -8133 10921 -8123
rect 10661 -8183 10691 -8163
rect 10641 -8223 10691 -8183
rect 10751 -8183 10781 -8163
rect 10751 -8223 10801 -8183
rect 10641 -8293 10801 -8223
rect 10641 -8333 10691 -8293
rect 10661 -8353 10691 -8333
rect 10751 -8333 10801 -8293
rect 10751 -8353 10781 -8333
rect 10861 -8393 10921 -8133
rect 10521 -8403 10601 -8393
rect 10521 -8463 10531 -8403
rect 10591 -8413 10601 -8403
rect 10841 -8403 10921 -8393
rect 10841 -8413 10851 -8403
rect 10591 -8463 10851 -8413
rect 10911 -8463 10921 -8403
rect 10521 -8473 10921 -8463
rect 10977 -8053 11377 -8043
rect 10977 -8113 10987 -8053
rect 11047 -8103 11307 -8053
rect 11047 -8113 11057 -8103
rect 10977 -8123 11057 -8113
rect 11297 -8113 11307 -8103
rect 11367 -8113 11377 -8053
rect 11297 -8123 11377 -8113
rect 10977 -8393 11037 -8123
rect 11307 -8133 11377 -8123
rect 11117 -8183 11147 -8163
rect 11097 -8223 11147 -8183
rect 11207 -8183 11237 -8163
rect 11207 -8223 11257 -8183
rect 11097 -8293 11257 -8223
rect 11097 -8333 11147 -8293
rect 11117 -8353 11147 -8333
rect 11207 -8333 11257 -8293
rect 11207 -8353 11237 -8333
rect 11317 -8393 11377 -8133
rect 10977 -8403 11057 -8393
rect 10977 -8463 10987 -8403
rect 11047 -8413 11057 -8403
rect 11297 -8403 11377 -8393
rect 11297 -8413 11307 -8403
rect 11047 -8463 11307 -8413
rect 11367 -8463 11377 -8403
rect 10977 -8473 11377 -8463
rect 11433 -8053 11833 -8043
rect 11433 -8113 11443 -8053
rect 11503 -8103 11763 -8053
rect 11503 -8113 11513 -8103
rect 11433 -8123 11513 -8113
rect 11753 -8113 11763 -8103
rect 11823 -8113 11833 -8053
rect 11753 -8123 11833 -8113
rect 11433 -8393 11493 -8123
rect 11763 -8133 11833 -8123
rect 11573 -8183 11603 -8163
rect 11553 -8223 11603 -8183
rect 11663 -8183 11693 -8163
rect 11663 -8223 11713 -8183
rect 11553 -8293 11713 -8223
rect 11553 -8333 11603 -8293
rect 11573 -8353 11603 -8333
rect 11663 -8333 11713 -8293
rect 11663 -8353 11693 -8333
rect 11773 -8393 11833 -8133
rect 11433 -8403 11513 -8393
rect 11433 -8463 11443 -8403
rect 11503 -8413 11513 -8403
rect 11753 -8403 11833 -8393
rect 11753 -8413 11763 -8403
rect 11503 -8463 11763 -8413
rect 11823 -8463 11833 -8403
rect 11433 -8473 11833 -8463
rect 11891 -8053 12291 -8043
rect 11891 -8113 11901 -8053
rect 11961 -8103 12221 -8053
rect 11961 -8113 11971 -8103
rect 11891 -8123 11971 -8113
rect 12211 -8113 12221 -8103
rect 12281 -8113 12291 -8053
rect 12211 -8123 12291 -8113
rect 11891 -8393 11951 -8123
rect 12221 -8133 12291 -8123
rect 12031 -8183 12061 -8163
rect 12011 -8223 12061 -8183
rect 12121 -8183 12151 -8163
rect 12121 -8223 12171 -8183
rect 12011 -8293 12171 -8223
rect 12011 -8333 12061 -8293
rect 12031 -8353 12061 -8333
rect 12121 -8333 12171 -8293
rect 12121 -8353 12151 -8333
rect 12231 -8393 12291 -8133
rect 11891 -8403 11971 -8393
rect 11891 -8463 11901 -8403
rect 11961 -8413 11971 -8403
rect 12211 -8403 12291 -8393
rect 12211 -8413 12221 -8403
rect 11961 -8463 12221 -8413
rect 12281 -8463 12291 -8403
rect 11891 -8473 12291 -8463
rect 12347 -8053 12747 -8043
rect 12347 -8113 12357 -8053
rect 12417 -8103 12677 -8053
rect 12417 -8113 12427 -8103
rect 12347 -8123 12427 -8113
rect 12667 -8113 12677 -8103
rect 12737 -8113 12747 -8053
rect 12667 -8123 12747 -8113
rect 12347 -8393 12407 -8123
rect 12677 -8133 12747 -8123
rect 12487 -8183 12517 -8163
rect 12467 -8223 12517 -8183
rect 12577 -8183 12607 -8163
rect 12577 -8223 12627 -8183
rect 12467 -8293 12627 -8223
rect 12467 -8333 12517 -8293
rect 12487 -8353 12517 -8333
rect 12577 -8333 12627 -8293
rect 12577 -8353 12607 -8333
rect 12687 -8393 12747 -8133
rect 12347 -8403 12427 -8393
rect 12347 -8463 12357 -8403
rect 12417 -8413 12427 -8403
rect 12667 -8403 12747 -8393
rect 12667 -8413 12677 -8403
rect 12417 -8463 12677 -8413
rect 12737 -8463 12747 -8403
rect 12347 -8473 12747 -8463
rect 12803 -8053 13203 -8043
rect 12803 -8113 12813 -8053
rect 12873 -8103 13133 -8053
rect 12873 -8113 12883 -8103
rect 12803 -8123 12883 -8113
rect 13123 -8113 13133 -8103
rect 13193 -8113 13203 -8053
rect 13123 -8123 13203 -8113
rect 12803 -8393 12863 -8123
rect 13133 -8133 13203 -8123
rect 12943 -8183 12973 -8163
rect 12923 -8223 12973 -8183
rect 13033 -8183 13063 -8163
rect 13033 -8223 13083 -8183
rect 12923 -8293 13083 -8223
rect 12923 -8333 12973 -8293
rect 12943 -8353 12973 -8333
rect 13033 -8333 13083 -8293
rect 13033 -8353 13063 -8333
rect 13143 -8393 13203 -8133
rect 12803 -8403 12883 -8393
rect 12803 -8463 12813 -8403
rect 12873 -8413 12883 -8403
rect 13123 -8403 13203 -8393
rect 13123 -8413 13133 -8403
rect 12873 -8463 13133 -8413
rect 13193 -8463 13203 -8403
rect 12803 -8473 13203 -8463
rect 13261 -8053 13661 -8043
rect 13261 -8113 13271 -8053
rect 13331 -8103 13591 -8053
rect 13331 -8113 13341 -8103
rect 13261 -8123 13341 -8113
rect 13581 -8113 13591 -8103
rect 13651 -8113 13661 -8053
rect 13581 -8123 13661 -8113
rect 13261 -8393 13321 -8123
rect 13591 -8133 13661 -8123
rect 13401 -8183 13431 -8163
rect 13381 -8223 13431 -8183
rect 13491 -8183 13521 -8163
rect 13491 -8223 13541 -8183
rect 13381 -8293 13541 -8223
rect 13381 -8333 13431 -8293
rect 13401 -8353 13431 -8333
rect 13491 -8333 13541 -8293
rect 13491 -8353 13521 -8333
rect 13601 -8393 13661 -8133
rect 13261 -8403 13341 -8393
rect 13261 -8463 13271 -8403
rect 13331 -8413 13341 -8403
rect 13581 -8403 13661 -8393
rect 13581 -8413 13591 -8403
rect 13331 -8463 13591 -8413
rect 13651 -8463 13661 -8403
rect 13261 -8473 13661 -8463
rect 13717 -8053 14117 -8043
rect 13717 -8113 13727 -8053
rect 13787 -8103 14047 -8053
rect 13787 -8113 13797 -8103
rect 13717 -8123 13797 -8113
rect 14037 -8113 14047 -8103
rect 14107 -8113 14117 -8053
rect 14037 -8123 14117 -8113
rect 13717 -8393 13777 -8123
rect 14047 -8133 14117 -8123
rect 13857 -8183 13887 -8163
rect 13837 -8223 13887 -8183
rect 13947 -8183 13977 -8163
rect 13947 -8223 13997 -8183
rect 13837 -8293 13997 -8223
rect 13837 -8333 13887 -8293
rect 13857 -8353 13887 -8333
rect 13947 -8333 13997 -8293
rect 13947 -8353 13977 -8333
rect 14057 -8393 14117 -8133
rect 13717 -8403 13797 -8393
rect 13717 -8463 13727 -8403
rect 13787 -8413 13797 -8403
rect 14037 -8403 14117 -8393
rect 14037 -8413 14047 -8403
rect 13787 -8463 14047 -8413
rect 14107 -8463 14117 -8403
rect 13717 -8473 14117 -8463
rect 14173 -8053 14573 -8043
rect 14173 -8113 14183 -8053
rect 14243 -8103 14503 -8053
rect 14243 -8113 14253 -8103
rect 14173 -8123 14253 -8113
rect 14493 -8113 14503 -8103
rect 14563 -8113 14573 -8053
rect 14493 -8123 14573 -8113
rect 14173 -8393 14233 -8123
rect 14503 -8133 14573 -8123
rect 14313 -8183 14343 -8163
rect 14293 -8223 14343 -8183
rect 14403 -8183 14433 -8163
rect 14403 -8223 14453 -8183
rect 14293 -8293 14453 -8223
rect 14293 -8333 14343 -8293
rect 14313 -8353 14343 -8333
rect 14403 -8333 14453 -8293
rect 14403 -8353 14433 -8333
rect 14513 -8393 14573 -8133
rect 14173 -8403 14253 -8393
rect 14173 -8463 14183 -8403
rect 14243 -8413 14253 -8403
rect 14493 -8403 14573 -8393
rect 14493 -8413 14503 -8403
rect 14243 -8463 14503 -8413
rect 14563 -8463 14573 -8403
rect 14173 -8473 14573 -8463
rect 14631 -8053 15031 -8043
rect 14631 -8113 14641 -8053
rect 14701 -8103 14961 -8053
rect 14701 -8113 14711 -8103
rect 14631 -8123 14711 -8113
rect 14951 -8113 14961 -8103
rect 15021 -8113 15031 -8053
rect 14951 -8123 15031 -8113
rect 14631 -8393 14691 -8123
rect 14961 -8133 15031 -8123
rect 14771 -8183 14801 -8163
rect 14751 -8223 14801 -8183
rect 14861 -8183 14891 -8163
rect 14861 -8223 14911 -8183
rect 14751 -8293 14911 -8223
rect 14751 -8333 14801 -8293
rect 14771 -8353 14801 -8333
rect 14861 -8333 14911 -8293
rect 14861 -8353 14891 -8333
rect 14971 -8393 15031 -8133
rect 14631 -8403 14711 -8393
rect 14631 -8463 14641 -8403
rect 14701 -8413 14711 -8403
rect 14951 -8403 15031 -8393
rect 14951 -8413 14961 -8403
rect 14701 -8463 14961 -8413
rect 15021 -8463 15031 -8403
rect 14631 -8473 15031 -8463
rect 15087 -8053 15487 -8043
rect 15087 -8113 15097 -8053
rect 15157 -8103 15417 -8053
rect 15157 -8113 15167 -8103
rect 15087 -8123 15167 -8113
rect 15407 -8113 15417 -8103
rect 15477 -8113 15487 -8053
rect 15407 -8123 15487 -8113
rect 15087 -8393 15147 -8123
rect 15417 -8133 15487 -8123
rect 15227 -8183 15257 -8163
rect 15207 -8223 15257 -8183
rect 15317 -8183 15347 -8163
rect 15317 -8223 15367 -8183
rect 15207 -8293 15367 -8223
rect 15207 -8333 15257 -8293
rect 15227 -8353 15257 -8333
rect 15317 -8333 15367 -8293
rect 15317 -8353 15347 -8333
rect 15427 -8393 15487 -8133
rect 15087 -8403 15167 -8393
rect 15087 -8463 15097 -8403
rect 15157 -8413 15167 -8403
rect 15407 -8403 15487 -8393
rect 15407 -8413 15417 -8403
rect 15157 -8463 15417 -8413
rect 15477 -8463 15487 -8403
rect 15087 -8473 15487 -8463
rect 1 -8547 401 -8537
rect 1 -8607 11 -8547
rect 71 -8597 331 -8547
rect 71 -8607 81 -8597
rect 1 -8617 81 -8607
rect 321 -8607 331 -8597
rect 391 -8607 401 -8547
rect 321 -8617 401 -8607
rect 1 -8887 61 -8617
rect 331 -8627 401 -8617
rect 141 -8677 171 -8657
rect 121 -8717 171 -8677
rect 231 -8677 261 -8657
rect 231 -8717 281 -8677
rect 121 -8787 281 -8717
rect 121 -8827 171 -8787
rect 141 -8847 171 -8827
rect 231 -8827 281 -8787
rect 231 -8847 261 -8827
rect 341 -8887 401 -8627
rect 1 -8897 81 -8887
rect 1 -8957 11 -8897
rect 71 -8907 81 -8897
rect 321 -8897 401 -8887
rect 321 -8907 331 -8897
rect 71 -8957 331 -8907
rect 391 -8957 401 -8897
rect 1 -8967 401 -8957
rect 457 -8547 857 -8537
rect 457 -8607 467 -8547
rect 527 -8597 787 -8547
rect 527 -8607 537 -8597
rect 457 -8617 537 -8607
rect 777 -8607 787 -8597
rect 847 -8607 857 -8547
rect 777 -8617 857 -8607
rect 457 -8887 517 -8617
rect 787 -8627 857 -8617
rect 597 -8677 627 -8657
rect 577 -8717 627 -8677
rect 687 -8677 717 -8657
rect 687 -8717 737 -8677
rect 577 -8787 737 -8717
rect 577 -8827 627 -8787
rect 597 -8847 627 -8827
rect 687 -8827 737 -8787
rect 687 -8847 717 -8827
rect 797 -8887 857 -8627
rect 457 -8897 537 -8887
rect 457 -8957 467 -8897
rect 527 -8907 537 -8897
rect 777 -8897 857 -8887
rect 777 -8907 787 -8897
rect 527 -8957 787 -8907
rect 847 -8957 857 -8897
rect 457 -8967 857 -8957
rect 913 -8547 1313 -8537
rect 913 -8607 923 -8547
rect 983 -8597 1243 -8547
rect 983 -8607 993 -8597
rect 913 -8617 993 -8607
rect 1233 -8607 1243 -8597
rect 1303 -8607 1313 -8547
rect 1233 -8617 1313 -8607
rect 913 -8887 973 -8617
rect 1243 -8627 1313 -8617
rect 1053 -8677 1083 -8657
rect 1033 -8717 1083 -8677
rect 1143 -8677 1173 -8657
rect 1143 -8717 1193 -8677
rect 1033 -8787 1193 -8717
rect 1033 -8827 1083 -8787
rect 1053 -8847 1083 -8827
rect 1143 -8827 1193 -8787
rect 1143 -8847 1173 -8827
rect 1253 -8887 1313 -8627
rect 913 -8897 993 -8887
rect 913 -8957 923 -8897
rect 983 -8907 993 -8897
rect 1233 -8897 1313 -8887
rect 1233 -8907 1243 -8897
rect 983 -8957 1243 -8907
rect 1303 -8957 1313 -8897
rect 913 -8967 1313 -8957
rect 1371 -8547 1771 -8537
rect 1371 -8607 1381 -8547
rect 1441 -8597 1701 -8547
rect 1441 -8607 1451 -8597
rect 1371 -8617 1451 -8607
rect 1691 -8607 1701 -8597
rect 1761 -8607 1771 -8547
rect 1691 -8617 1771 -8607
rect 1371 -8887 1431 -8617
rect 1701 -8627 1771 -8617
rect 1511 -8677 1541 -8657
rect 1491 -8717 1541 -8677
rect 1601 -8677 1631 -8657
rect 1601 -8717 1651 -8677
rect 1491 -8787 1651 -8717
rect 1491 -8827 1541 -8787
rect 1511 -8847 1541 -8827
rect 1601 -8827 1651 -8787
rect 1601 -8847 1631 -8827
rect 1711 -8887 1771 -8627
rect 1371 -8897 1451 -8887
rect 1371 -8957 1381 -8897
rect 1441 -8907 1451 -8897
rect 1691 -8897 1771 -8887
rect 1691 -8907 1701 -8897
rect 1441 -8957 1701 -8907
rect 1761 -8957 1771 -8897
rect 1371 -8967 1771 -8957
rect 1827 -8547 2227 -8537
rect 1827 -8607 1837 -8547
rect 1897 -8597 2157 -8547
rect 1897 -8607 1907 -8597
rect 1827 -8617 1907 -8607
rect 2147 -8607 2157 -8597
rect 2217 -8607 2227 -8547
rect 2147 -8617 2227 -8607
rect 1827 -8887 1887 -8617
rect 2157 -8627 2227 -8617
rect 1967 -8677 1997 -8657
rect 1947 -8717 1997 -8677
rect 2057 -8677 2087 -8657
rect 2057 -8717 2107 -8677
rect 1947 -8787 2107 -8717
rect 1947 -8827 1997 -8787
rect 1967 -8847 1997 -8827
rect 2057 -8827 2107 -8787
rect 2057 -8847 2087 -8827
rect 2167 -8887 2227 -8627
rect 1827 -8897 1907 -8887
rect 1827 -8957 1837 -8897
rect 1897 -8907 1907 -8897
rect 2147 -8897 2227 -8887
rect 2147 -8907 2157 -8897
rect 1897 -8957 2157 -8907
rect 2217 -8957 2227 -8897
rect 1827 -8967 2227 -8957
rect 2283 -8547 2683 -8537
rect 2283 -8607 2293 -8547
rect 2353 -8597 2613 -8547
rect 2353 -8607 2363 -8597
rect 2283 -8617 2363 -8607
rect 2603 -8607 2613 -8597
rect 2673 -8607 2683 -8547
rect 2603 -8617 2683 -8607
rect 2283 -8887 2343 -8617
rect 2613 -8627 2683 -8617
rect 2423 -8677 2453 -8657
rect 2403 -8717 2453 -8677
rect 2513 -8677 2543 -8657
rect 2513 -8717 2563 -8677
rect 2403 -8787 2563 -8717
rect 2403 -8827 2453 -8787
rect 2423 -8847 2453 -8827
rect 2513 -8827 2563 -8787
rect 2513 -8847 2543 -8827
rect 2623 -8887 2683 -8627
rect 2283 -8897 2363 -8887
rect 2283 -8957 2293 -8897
rect 2353 -8907 2363 -8897
rect 2603 -8897 2683 -8887
rect 2603 -8907 2613 -8897
rect 2353 -8957 2613 -8907
rect 2673 -8957 2683 -8897
rect 2283 -8967 2683 -8957
rect 2741 -8547 3141 -8537
rect 2741 -8607 2751 -8547
rect 2811 -8597 3071 -8547
rect 2811 -8607 2821 -8597
rect 2741 -8617 2821 -8607
rect 3061 -8607 3071 -8597
rect 3131 -8607 3141 -8547
rect 3061 -8617 3141 -8607
rect 2741 -8887 2801 -8617
rect 3071 -8627 3141 -8617
rect 2881 -8677 2911 -8657
rect 2861 -8717 2911 -8677
rect 2971 -8677 3001 -8657
rect 2971 -8717 3021 -8677
rect 2861 -8787 3021 -8717
rect 2861 -8827 2911 -8787
rect 2881 -8847 2911 -8827
rect 2971 -8827 3021 -8787
rect 2971 -8847 3001 -8827
rect 3081 -8887 3141 -8627
rect 2741 -8897 2821 -8887
rect 2741 -8957 2751 -8897
rect 2811 -8907 2821 -8897
rect 3061 -8897 3141 -8887
rect 3061 -8907 3071 -8897
rect 2811 -8957 3071 -8907
rect 3131 -8957 3141 -8897
rect 2741 -8967 3141 -8957
rect 3197 -8547 3597 -8537
rect 3197 -8607 3207 -8547
rect 3267 -8597 3527 -8547
rect 3267 -8607 3277 -8597
rect 3197 -8617 3277 -8607
rect 3517 -8607 3527 -8597
rect 3587 -8607 3597 -8547
rect 3517 -8617 3597 -8607
rect 3197 -8887 3257 -8617
rect 3527 -8627 3597 -8617
rect 3337 -8677 3367 -8657
rect 3317 -8717 3367 -8677
rect 3427 -8677 3457 -8657
rect 3427 -8717 3477 -8677
rect 3317 -8787 3477 -8717
rect 3317 -8827 3367 -8787
rect 3337 -8847 3367 -8827
rect 3427 -8827 3477 -8787
rect 3427 -8847 3457 -8827
rect 3537 -8887 3597 -8627
rect 3197 -8897 3277 -8887
rect 3197 -8957 3207 -8897
rect 3267 -8907 3277 -8897
rect 3517 -8897 3597 -8887
rect 3517 -8907 3527 -8897
rect 3267 -8957 3527 -8907
rect 3587 -8957 3597 -8897
rect 3197 -8967 3597 -8957
rect 3653 -8547 4053 -8537
rect 3653 -8607 3663 -8547
rect 3723 -8597 3983 -8547
rect 3723 -8607 3733 -8597
rect 3653 -8617 3733 -8607
rect 3973 -8607 3983 -8597
rect 4043 -8607 4053 -8547
rect 3973 -8617 4053 -8607
rect 3653 -8887 3713 -8617
rect 3983 -8627 4053 -8617
rect 3793 -8677 3823 -8657
rect 3773 -8717 3823 -8677
rect 3883 -8677 3913 -8657
rect 3883 -8717 3933 -8677
rect 3773 -8787 3933 -8717
rect 3773 -8827 3823 -8787
rect 3793 -8847 3823 -8827
rect 3883 -8827 3933 -8787
rect 3883 -8847 3913 -8827
rect 3993 -8887 4053 -8627
rect 3653 -8897 3733 -8887
rect 3653 -8957 3663 -8897
rect 3723 -8907 3733 -8897
rect 3973 -8897 4053 -8887
rect 3973 -8907 3983 -8897
rect 3723 -8957 3983 -8907
rect 4043 -8957 4053 -8897
rect 3653 -8967 4053 -8957
rect 4111 -8547 4511 -8537
rect 4111 -8607 4121 -8547
rect 4181 -8597 4441 -8547
rect 4181 -8607 4191 -8597
rect 4111 -8617 4191 -8607
rect 4431 -8607 4441 -8597
rect 4501 -8607 4511 -8547
rect 4431 -8617 4511 -8607
rect 4111 -8887 4171 -8617
rect 4441 -8627 4511 -8617
rect 4251 -8677 4281 -8657
rect 4231 -8717 4281 -8677
rect 4341 -8677 4371 -8657
rect 4341 -8717 4391 -8677
rect 4231 -8787 4391 -8717
rect 4231 -8827 4281 -8787
rect 4251 -8847 4281 -8827
rect 4341 -8827 4391 -8787
rect 4341 -8847 4371 -8827
rect 4451 -8887 4511 -8627
rect 4111 -8897 4191 -8887
rect 4111 -8957 4121 -8897
rect 4181 -8907 4191 -8897
rect 4431 -8897 4511 -8887
rect 4431 -8907 4441 -8897
rect 4181 -8957 4441 -8907
rect 4501 -8957 4511 -8897
rect 4111 -8967 4511 -8957
rect 4567 -8547 4967 -8537
rect 4567 -8607 4577 -8547
rect 4637 -8597 4897 -8547
rect 4637 -8607 4647 -8597
rect 4567 -8617 4647 -8607
rect 4887 -8607 4897 -8597
rect 4957 -8607 4967 -8547
rect 4887 -8617 4967 -8607
rect 4567 -8887 4627 -8617
rect 4897 -8627 4967 -8617
rect 4707 -8677 4737 -8657
rect 4687 -8717 4737 -8677
rect 4797 -8677 4827 -8657
rect 4797 -8717 4847 -8677
rect 4687 -8787 4847 -8717
rect 4687 -8827 4737 -8787
rect 4707 -8847 4737 -8827
rect 4797 -8827 4847 -8787
rect 4797 -8847 4827 -8827
rect 4907 -8887 4967 -8627
rect 4567 -8897 4647 -8887
rect 4567 -8957 4577 -8897
rect 4637 -8907 4647 -8897
rect 4887 -8897 4967 -8887
rect 4887 -8907 4897 -8897
rect 4637 -8957 4897 -8907
rect 4957 -8957 4967 -8897
rect 4567 -8967 4967 -8957
rect 5023 -8547 5423 -8537
rect 5023 -8607 5033 -8547
rect 5093 -8597 5353 -8547
rect 5093 -8607 5103 -8597
rect 5023 -8617 5103 -8607
rect 5343 -8607 5353 -8597
rect 5413 -8607 5423 -8547
rect 5343 -8617 5423 -8607
rect 5023 -8887 5083 -8617
rect 5353 -8627 5423 -8617
rect 5163 -8677 5193 -8657
rect 5143 -8717 5193 -8677
rect 5253 -8677 5283 -8657
rect 5253 -8717 5303 -8677
rect 5143 -8787 5303 -8717
rect 5143 -8827 5193 -8787
rect 5163 -8847 5193 -8827
rect 5253 -8827 5303 -8787
rect 5253 -8847 5283 -8827
rect 5363 -8887 5423 -8627
rect 5023 -8897 5103 -8887
rect 5023 -8957 5033 -8897
rect 5093 -8907 5103 -8897
rect 5343 -8897 5423 -8887
rect 5343 -8907 5353 -8897
rect 5093 -8957 5353 -8907
rect 5413 -8957 5423 -8897
rect 5023 -8967 5423 -8957
rect 5481 -8547 5881 -8537
rect 5481 -8607 5491 -8547
rect 5551 -8597 5811 -8547
rect 5551 -8607 5561 -8597
rect 5481 -8617 5561 -8607
rect 5801 -8607 5811 -8597
rect 5871 -8607 5881 -8547
rect 5801 -8617 5881 -8607
rect 5481 -8887 5541 -8617
rect 5811 -8627 5881 -8617
rect 5621 -8677 5651 -8657
rect 5601 -8717 5651 -8677
rect 5711 -8677 5741 -8657
rect 5711 -8717 5761 -8677
rect 5601 -8787 5761 -8717
rect 5601 -8827 5651 -8787
rect 5621 -8847 5651 -8827
rect 5711 -8827 5761 -8787
rect 5711 -8847 5741 -8827
rect 5821 -8887 5881 -8627
rect 5481 -8897 5561 -8887
rect 5481 -8957 5491 -8897
rect 5551 -8907 5561 -8897
rect 5801 -8897 5881 -8887
rect 5801 -8907 5811 -8897
rect 5551 -8957 5811 -8907
rect 5871 -8957 5881 -8897
rect 5481 -8967 5881 -8957
rect 5937 -8547 6337 -8537
rect 5937 -8607 5947 -8547
rect 6007 -8597 6267 -8547
rect 6007 -8607 6017 -8597
rect 5937 -8617 6017 -8607
rect 6257 -8607 6267 -8597
rect 6327 -8607 6337 -8547
rect 6257 -8617 6337 -8607
rect 5937 -8887 5997 -8617
rect 6267 -8627 6337 -8617
rect 6077 -8677 6107 -8657
rect 6057 -8717 6107 -8677
rect 6167 -8677 6197 -8657
rect 6167 -8717 6217 -8677
rect 6057 -8787 6217 -8717
rect 6057 -8827 6107 -8787
rect 6077 -8847 6107 -8827
rect 6167 -8827 6217 -8787
rect 6167 -8847 6197 -8827
rect 6277 -8887 6337 -8627
rect 5937 -8897 6017 -8887
rect 5937 -8957 5947 -8897
rect 6007 -8907 6017 -8897
rect 6257 -8897 6337 -8887
rect 6257 -8907 6267 -8897
rect 6007 -8957 6267 -8907
rect 6327 -8957 6337 -8897
rect 5937 -8967 6337 -8957
rect 6393 -8547 6793 -8537
rect 6393 -8607 6403 -8547
rect 6463 -8597 6723 -8547
rect 6463 -8607 6473 -8597
rect 6393 -8617 6473 -8607
rect 6713 -8607 6723 -8597
rect 6783 -8607 6793 -8547
rect 6713 -8617 6793 -8607
rect 6393 -8887 6453 -8617
rect 6723 -8627 6793 -8617
rect 6533 -8677 6563 -8657
rect 6513 -8717 6563 -8677
rect 6623 -8677 6653 -8657
rect 6623 -8717 6673 -8677
rect 6513 -8787 6673 -8717
rect 6513 -8827 6563 -8787
rect 6533 -8847 6563 -8827
rect 6623 -8827 6673 -8787
rect 6623 -8847 6653 -8827
rect 6733 -8887 6793 -8627
rect 6393 -8897 6473 -8887
rect 6393 -8957 6403 -8897
rect 6463 -8907 6473 -8897
rect 6713 -8897 6793 -8887
rect 6713 -8907 6723 -8897
rect 6463 -8957 6723 -8907
rect 6783 -8957 6793 -8897
rect 6393 -8967 6793 -8957
rect 6851 -8547 7251 -8537
rect 6851 -8607 6861 -8547
rect 6921 -8597 7181 -8547
rect 6921 -8607 6931 -8597
rect 6851 -8617 6931 -8607
rect 7171 -8607 7181 -8597
rect 7241 -8607 7251 -8547
rect 7171 -8617 7251 -8607
rect 6851 -8887 6911 -8617
rect 7181 -8627 7251 -8617
rect 6991 -8677 7021 -8657
rect 6971 -8717 7021 -8677
rect 7081 -8677 7111 -8657
rect 7081 -8717 7131 -8677
rect 6971 -8787 7131 -8717
rect 6971 -8827 7021 -8787
rect 6991 -8847 7021 -8827
rect 7081 -8827 7131 -8787
rect 7081 -8847 7111 -8827
rect 7191 -8887 7251 -8627
rect 6851 -8897 6931 -8887
rect 6851 -8957 6861 -8897
rect 6921 -8907 6931 -8897
rect 7171 -8897 7251 -8887
rect 7171 -8907 7181 -8897
rect 6921 -8957 7181 -8907
rect 7241 -8957 7251 -8897
rect 6851 -8967 7251 -8957
rect 7307 -8547 7707 -8537
rect 7307 -8607 7317 -8547
rect 7377 -8597 7637 -8547
rect 7377 -8607 7387 -8597
rect 7307 -8617 7387 -8607
rect 7627 -8607 7637 -8597
rect 7697 -8607 7707 -8547
rect 7627 -8617 7707 -8607
rect 7307 -8887 7367 -8617
rect 7637 -8627 7707 -8617
rect 7447 -8677 7477 -8657
rect 7427 -8717 7477 -8677
rect 7537 -8677 7567 -8657
rect 7537 -8717 7587 -8677
rect 7427 -8787 7587 -8717
rect 7427 -8827 7477 -8787
rect 7447 -8847 7477 -8827
rect 7537 -8827 7587 -8787
rect 7537 -8847 7567 -8827
rect 7647 -8887 7707 -8627
rect 7307 -8897 7387 -8887
rect 7307 -8957 7317 -8897
rect 7377 -8907 7387 -8897
rect 7627 -8897 7707 -8887
rect 7627 -8907 7637 -8897
rect 7377 -8957 7637 -8907
rect 7697 -8957 7707 -8897
rect 7307 -8967 7707 -8957
rect 7763 -8547 8163 -8537
rect 7763 -8607 7773 -8547
rect 7833 -8597 8093 -8547
rect 7833 -8607 7843 -8597
rect 7763 -8617 7843 -8607
rect 8083 -8607 8093 -8597
rect 8153 -8607 8163 -8547
rect 8083 -8617 8163 -8607
rect 7763 -8887 7823 -8617
rect 8093 -8627 8163 -8617
rect 7903 -8677 7933 -8657
rect 7883 -8717 7933 -8677
rect 7993 -8677 8023 -8657
rect 7993 -8717 8043 -8677
rect 7883 -8787 8043 -8717
rect 7883 -8827 7933 -8787
rect 7903 -8847 7933 -8827
rect 7993 -8827 8043 -8787
rect 7993 -8847 8023 -8827
rect 8103 -8887 8163 -8627
rect 7763 -8897 7843 -8887
rect 7763 -8957 7773 -8897
rect 7833 -8907 7843 -8897
rect 8083 -8897 8163 -8887
rect 8083 -8907 8093 -8897
rect 7833 -8957 8093 -8907
rect 8153 -8957 8163 -8897
rect 7763 -8967 8163 -8957
rect 8237 -8547 8637 -8537
rect 8237 -8607 8247 -8547
rect 8307 -8597 8567 -8547
rect 8307 -8607 8317 -8597
rect 8237 -8617 8317 -8607
rect 8557 -8607 8567 -8597
rect 8627 -8607 8637 -8547
rect 8557 -8617 8637 -8607
rect 8237 -8887 8297 -8617
rect 8567 -8627 8637 -8617
rect 8377 -8677 8407 -8657
rect 8357 -8717 8407 -8677
rect 8467 -8677 8497 -8657
rect 8467 -8717 8517 -8677
rect 8357 -8787 8517 -8717
rect 8357 -8827 8407 -8787
rect 8377 -8847 8407 -8827
rect 8467 -8827 8517 -8787
rect 8467 -8847 8497 -8827
rect 8577 -8887 8637 -8627
rect 8237 -8897 8317 -8887
rect 8237 -8957 8247 -8897
rect 8307 -8907 8317 -8897
rect 8557 -8897 8637 -8887
rect 8557 -8907 8567 -8897
rect 8307 -8957 8567 -8907
rect 8627 -8957 8637 -8897
rect 8237 -8967 8637 -8957
rect 8693 -8547 9093 -8537
rect 8693 -8607 8703 -8547
rect 8763 -8597 9023 -8547
rect 8763 -8607 8773 -8597
rect 8693 -8617 8773 -8607
rect 9013 -8607 9023 -8597
rect 9083 -8607 9093 -8547
rect 9013 -8617 9093 -8607
rect 8693 -8887 8753 -8617
rect 9023 -8627 9093 -8617
rect 8833 -8677 8863 -8657
rect 8813 -8717 8863 -8677
rect 8923 -8677 8953 -8657
rect 8923 -8717 8973 -8677
rect 8813 -8787 8973 -8717
rect 8813 -8827 8863 -8787
rect 8833 -8847 8863 -8827
rect 8923 -8827 8973 -8787
rect 8923 -8847 8953 -8827
rect 9033 -8887 9093 -8627
rect 8693 -8897 8773 -8887
rect 8693 -8957 8703 -8897
rect 8763 -8907 8773 -8897
rect 9013 -8897 9093 -8887
rect 9013 -8907 9023 -8897
rect 8763 -8957 9023 -8907
rect 9083 -8957 9093 -8897
rect 8693 -8967 9093 -8957
rect 9151 -8547 9551 -8537
rect 9151 -8607 9161 -8547
rect 9221 -8597 9481 -8547
rect 9221 -8607 9231 -8597
rect 9151 -8617 9231 -8607
rect 9471 -8607 9481 -8597
rect 9541 -8607 9551 -8547
rect 9471 -8617 9551 -8607
rect 9151 -8887 9211 -8617
rect 9481 -8627 9551 -8617
rect 9291 -8677 9321 -8657
rect 9271 -8717 9321 -8677
rect 9381 -8677 9411 -8657
rect 9381 -8717 9431 -8677
rect 9271 -8787 9431 -8717
rect 9271 -8827 9321 -8787
rect 9291 -8847 9321 -8827
rect 9381 -8827 9431 -8787
rect 9381 -8847 9411 -8827
rect 9491 -8887 9551 -8627
rect 9151 -8897 9231 -8887
rect 9151 -8957 9161 -8897
rect 9221 -8907 9231 -8897
rect 9471 -8897 9551 -8887
rect 9471 -8907 9481 -8897
rect 9221 -8957 9481 -8907
rect 9541 -8957 9551 -8897
rect 9151 -8967 9551 -8957
rect 9607 -8547 10007 -8537
rect 9607 -8607 9617 -8547
rect 9677 -8597 9937 -8547
rect 9677 -8607 9687 -8597
rect 9607 -8617 9687 -8607
rect 9927 -8607 9937 -8597
rect 9997 -8607 10007 -8547
rect 9927 -8617 10007 -8607
rect 9607 -8887 9667 -8617
rect 9937 -8627 10007 -8617
rect 9747 -8677 9777 -8657
rect 9727 -8717 9777 -8677
rect 9837 -8677 9867 -8657
rect 9837 -8717 9887 -8677
rect 9727 -8787 9887 -8717
rect 9727 -8827 9777 -8787
rect 9747 -8847 9777 -8827
rect 9837 -8827 9887 -8787
rect 9837 -8847 9867 -8827
rect 9947 -8887 10007 -8627
rect 9607 -8897 9687 -8887
rect 9607 -8957 9617 -8897
rect 9677 -8907 9687 -8897
rect 9927 -8897 10007 -8887
rect 9927 -8907 9937 -8897
rect 9677 -8957 9937 -8907
rect 9997 -8957 10007 -8897
rect 9607 -8967 10007 -8957
rect 10063 -8547 10463 -8537
rect 10063 -8607 10073 -8547
rect 10133 -8597 10393 -8547
rect 10133 -8607 10143 -8597
rect 10063 -8617 10143 -8607
rect 10383 -8607 10393 -8597
rect 10453 -8607 10463 -8547
rect 10383 -8617 10463 -8607
rect 10063 -8887 10123 -8617
rect 10393 -8627 10463 -8617
rect 10203 -8677 10233 -8657
rect 10183 -8717 10233 -8677
rect 10293 -8677 10323 -8657
rect 10293 -8717 10343 -8677
rect 10183 -8787 10343 -8717
rect 10183 -8827 10233 -8787
rect 10203 -8847 10233 -8827
rect 10293 -8827 10343 -8787
rect 10293 -8847 10323 -8827
rect 10403 -8887 10463 -8627
rect 10063 -8897 10143 -8887
rect 10063 -8957 10073 -8897
rect 10133 -8907 10143 -8897
rect 10383 -8897 10463 -8887
rect 10383 -8907 10393 -8897
rect 10133 -8957 10393 -8907
rect 10453 -8957 10463 -8897
rect 10063 -8967 10463 -8957
rect 10521 -8547 10921 -8537
rect 10521 -8607 10531 -8547
rect 10591 -8597 10851 -8547
rect 10591 -8607 10601 -8597
rect 10521 -8617 10601 -8607
rect 10841 -8607 10851 -8597
rect 10911 -8607 10921 -8547
rect 10841 -8617 10921 -8607
rect 10521 -8887 10581 -8617
rect 10851 -8627 10921 -8617
rect 10661 -8677 10691 -8657
rect 10641 -8717 10691 -8677
rect 10751 -8677 10781 -8657
rect 10751 -8717 10801 -8677
rect 10641 -8787 10801 -8717
rect 10641 -8827 10691 -8787
rect 10661 -8847 10691 -8827
rect 10751 -8827 10801 -8787
rect 10751 -8847 10781 -8827
rect 10861 -8887 10921 -8627
rect 10521 -8897 10601 -8887
rect 10521 -8957 10531 -8897
rect 10591 -8907 10601 -8897
rect 10841 -8897 10921 -8887
rect 10841 -8907 10851 -8897
rect 10591 -8957 10851 -8907
rect 10911 -8957 10921 -8897
rect 10521 -8967 10921 -8957
rect 10977 -8547 11377 -8537
rect 10977 -8607 10987 -8547
rect 11047 -8597 11307 -8547
rect 11047 -8607 11057 -8597
rect 10977 -8617 11057 -8607
rect 11297 -8607 11307 -8597
rect 11367 -8607 11377 -8547
rect 11297 -8617 11377 -8607
rect 10977 -8887 11037 -8617
rect 11307 -8627 11377 -8617
rect 11117 -8677 11147 -8657
rect 11097 -8717 11147 -8677
rect 11207 -8677 11237 -8657
rect 11207 -8717 11257 -8677
rect 11097 -8787 11257 -8717
rect 11097 -8827 11147 -8787
rect 11117 -8847 11147 -8827
rect 11207 -8827 11257 -8787
rect 11207 -8847 11237 -8827
rect 11317 -8887 11377 -8627
rect 10977 -8897 11057 -8887
rect 10977 -8957 10987 -8897
rect 11047 -8907 11057 -8897
rect 11297 -8897 11377 -8887
rect 11297 -8907 11307 -8897
rect 11047 -8957 11307 -8907
rect 11367 -8957 11377 -8897
rect 10977 -8967 11377 -8957
rect 11433 -8547 11833 -8537
rect 11433 -8607 11443 -8547
rect 11503 -8597 11763 -8547
rect 11503 -8607 11513 -8597
rect 11433 -8617 11513 -8607
rect 11753 -8607 11763 -8597
rect 11823 -8607 11833 -8547
rect 11753 -8617 11833 -8607
rect 11433 -8887 11493 -8617
rect 11763 -8627 11833 -8617
rect 11573 -8677 11603 -8657
rect 11553 -8717 11603 -8677
rect 11663 -8677 11693 -8657
rect 11663 -8717 11713 -8677
rect 11553 -8787 11713 -8717
rect 11553 -8827 11603 -8787
rect 11573 -8847 11603 -8827
rect 11663 -8827 11713 -8787
rect 11663 -8847 11693 -8827
rect 11773 -8887 11833 -8627
rect 11433 -8897 11513 -8887
rect 11433 -8957 11443 -8897
rect 11503 -8907 11513 -8897
rect 11753 -8897 11833 -8887
rect 11753 -8907 11763 -8897
rect 11503 -8957 11763 -8907
rect 11823 -8957 11833 -8897
rect 11433 -8967 11833 -8957
rect 11891 -8547 12291 -8537
rect 11891 -8607 11901 -8547
rect 11961 -8597 12221 -8547
rect 11961 -8607 11971 -8597
rect 11891 -8617 11971 -8607
rect 12211 -8607 12221 -8597
rect 12281 -8607 12291 -8547
rect 12211 -8617 12291 -8607
rect 11891 -8887 11951 -8617
rect 12221 -8627 12291 -8617
rect 12031 -8677 12061 -8657
rect 12011 -8717 12061 -8677
rect 12121 -8677 12151 -8657
rect 12121 -8717 12171 -8677
rect 12011 -8787 12171 -8717
rect 12011 -8827 12061 -8787
rect 12031 -8847 12061 -8827
rect 12121 -8827 12171 -8787
rect 12121 -8847 12151 -8827
rect 12231 -8887 12291 -8627
rect 11891 -8897 11971 -8887
rect 11891 -8957 11901 -8897
rect 11961 -8907 11971 -8897
rect 12211 -8897 12291 -8887
rect 12211 -8907 12221 -8897
rect 11961 -8957 12221 -8907
rect 12281 -8957 12291 -8897
rect 11891 -8967 12291 -8957
rect 12347 -8547 12747 -8537
rect 12347 -8607 12357 -8547
rect 12417 -8597 12677 -8547
rect 12417 -8607 12427 -8597
rect 12347 -8617 12427 -8607
rect 12667 -8607 12677 -8597
rect 12737 -8607 12747 -8547
rect 12667 -8617 12747 -8607
rect 12347 -8887 12407 -8617
rect 12677 -8627 12747 -8617
rect 12487 -8677 12517 -8657
rect 12467 -8717 12517 -8677
rect 12577 -8677 12607 -8657
rect 12577 -8717 12627 -8677
rect 12467 -8787 12627 -8717
rect 12467 -8827 12517 -8787
rect 12487 -8847 12517 -8827
rect 12577 -8827 12627 -8787
rect 12577 -8847 12607 -8827
rect 12687 -8887 12747 -8627
rect 12347 -8897 12427 -8887
rect 12347 -8957 12357 -8897
rect 12417 -8907 12427 -8897
rect 12667 -8897 12747 -8887
rect 12667 -8907 12677 -8897
rect 12417 -8957 12677 -8907
rect 12737 -8957 12747 -8897
rect 12347 -8967 12747 -8957
rect 12803 -8547 13203 -8537
rect 12803 -8607 12813 -8547
rect 12873 -8597 13133 -8547
rect 12873 -8607 12883 -8597
rect 12803 -8617 12883 -8607
rect 13123 -8607 13133 -8597
rect 13193 -8607 13203 -8547
rect 13123 -8617 13203 -8607
rect 12803 -8887 12863 -8617
rect 13133 -8627 13203 -8617
rect 12943 -8677 12973 -8657
rect 12923 -8717 12973 -8677
rect 13033 -8677 13063 -8657
rect 13033 -8717 13083 -8677
rect 12923 -8787 13083 -8717
rect 12923 -8827 12973 -8787
rect 12943 -8847 12973 -8827
rect 13033 -8827 13083 -8787
rect 13033 -8847 13063 -8827
rect 13143 -8887 13203 -8627
rect 12803 -8897 12883 -8887
rect 12803 -8957 12813 -8897
rect 12873 -8907 12883 -8897
rect 13123 -8897 13203 -8887
rect 13123 -8907 13133 -8897
rect 12873 -8957 13133 -8907
rect 13193 -8957 13203 -8897
rect 12803 -8967 13203 -8957
rect 13261 -8547 13661 -8537
rect 13261 -8607 13271 -8547
rect 13331 -8597 13591 -8547
rect 13331 -8607 13341 -8597
rect 13261 -8617 13341 -8607
rect 13581 -8607 13591 -8597
rect 13651 -8607 13661 -8547
rect 13581 -8617 13661 -8607
rect 13261 -8887 13321 -8617
rect 13591 -8627 13661 -8617
rect 13401 -8677 13431 -8657
rect 13381 -8717 13431 -8677
rect 13491 -8677 13521 -8657
rect 13491 -8717 13541 -8677
rect 13381 -8787 13541 -8717
rect 13381 -8827 13431 -8787
rect 13401 -8847 13431 -8827
rect 13491 -8827 13541 -8787
rect 13491 -8847 13521 -8827
rect 13601 -8887 13661 -8627
rect 13261 -8897 13341 -8887
rect 13261 -8957 13271 -8897
rect 13331 -8907 13341 -8897
rect 13581 -8897 13661 -8887
rect 13581 -8907 13591 -8897
rect 13331 -8957 13591 -8907
rect 13651 -8957 13661 -8897
rect 13261 -8967 13661 -8957
rect 13717 -8547 14117 -8537
rect 13717 -8607 13727 -8547
rect 13787 -8597 14047 -8547
rect 13787 -8607 13797 -8597
rect 13717 -8617 13797 -8607
rect 14037 -8607 14047 -8597
rect 14107 -8607 14117 -8547
rect 14037 -8617 14117 -8607
rect 13717 -8887 13777 -8617
rect 14047 -8627 14117 -8617
rect 13857 -8677 13887 -8657
rect 13837 -8717 13887 -8677
rect 13947 -8677 13977 -8657
rect 13947 -8717 13997 -8677
rect 13837 -8787 13997 -8717
rect 13837 -8827 13887 -8787
rect 13857 -8847 13887 -8827
rect 13947 -8827 13997 -8787
rect 13947 -8847 13977 -8827
rect 14057 -8887 14117 -8627
rect 13717 -8897 13797 -8887
rect 13717 -8957 13727 -8897
rect 13787 -8907 13797 -8897
rect 14037 -8897 14117 -8887
rect 14037 -8907 14047 -8897
rect 13787 -8957 14047 -8907
rect 14107 -8957 14117 -8897
rect 13717 -8967 14117 -8957
rect 14173 -8547 14573 -8537
rect 14173 -8607 14183 -8547
rect 14243 -8597 14503 -8547
rect 14243 -8607 14253 -8597
rect 14173 -8617 14253 -8607
rect 14493 -8607 14503 -8597
rect 14563 -8607 14573 -8547
rect 14493 -8617 14573 -8607
rect 14173 -8887 14233 -8617
rect 14503 -8627 14573 -8617
rect 14313 -8677 14343 -8657
rect 14293 -8717 14343 -8677
rect 14403 -8677 14433 -8657
rect 14403 -8717 14453 -8677
rect 14293 -8787 14453 -8717
rect 14293 -8827 14343 -8787
rect 14313 -8847 14343 -8827
rect 14403 -8827 14453 -8787
rect 14403 -8847 14433 -8827
rect 14513 -8887 14573 -8627
rect 14173 -8897 14253 -8887
rect 14173 -8957 14183 -8897
rect 14243 -8907 14253 -8897
rect 14493 -8897 14573 -8887
rect 14493 -8907 14503 -8897
rect 14243 -8957 14503 -8907
rect 14563 -8957 14573 -8897
rect 14173 -8967 14573 -8957
rect 14631 -8547 15031 -8537
rect 14631 -8607 14641 -8547
rect 14701 -8597 14961 -8547
rect 14701 -8607 14711 -8597
rect 14631 -8617 14711 -8607
rect 14951 -8607 14961 -8597
rect 15021 -8607 15031 -8547
rect 14951 -8617 15031 -8607
rect 14631 -8887 14691 -8617
rect 14961 -8627 15031 -8617
rect 14771 -8677 14801 -8657
rect 14751 -8717 14801 -8677
rect 14861 -8677 14891 -8657
rect 14861 -8717 14911 -8677
rect 14751 -8787 14911 -8717
rect 14751 -8827 14801 -8787
rect 14771 -8847 14801 -8827
rect 14861 -8827 14911 -8787
rect 14861 -8847 14891 -8827
rect 14971 -8887 15031 -8627
rect 14631 -8897 14711 -8887
rect 14631 -8957 14641 -8897
rect 14701 -8907 14711 -8897
rect 14951 -8897 15031 -8887
rect 14951 -8907 14961 -8897
rect 14701 -8957 14961 -8907
rect 15021 -8957 15031 -8897
rect 14631 -8967 15031 -8957
rect 15087 -8547 15487 -8537
rect 15087 -8607 15097 -8547
rect 15157 -8597 15417 -8547
rect 15157 -8607 15167 -8597
rect 15087 -8617 15167 -8607
rect 15407 -8607 15417 -8597
rect 15477 -8607 15487 -8547
rect 15407 -8617 15487 -8607
rect 15087 -8887 15147 -8617
rect 15417 -8627 15487 -8617
rect 15227 -8677 15257 -8657
rect 15207 -8717 15257 -8677
rect 15317 -8677 15347 -8657
rect 15317 -8717 15367 -8677
rect 15207 -8787 15367 -8717
rect 15207 -8827 15257 -8787
rect 15227 -8847 15257 -8827
rect 15317 -8827 15367 -8787
rect 15317 -8847 15347 -8827
rect 15427 -8887 15487 -8627
rect 15087 -8897 15167 -8887
rect 15087 -8957 15097 -8897
rect 15157 -8907 15167 -8897
rect 15407 -8897 15487 -8887
rect 15407 -8907 15417 -8897
rect 15157 -8957 15417 -8907
rect 15477 -8957 15487 -8897
rect 15087 -8967 15487 -8957
rect 1 -9049 401 -9039
rect 1 -9109 11 -9049
rect 71 -9099 331 -9049
rect 71 -9109 81 -9099
rect 1 -9119 81 -9109
rect 321 -9109 331 -9099
rect 391 -9109 401 -9049
rect 321 -9119 401 -9109
rect 1 -9389 61 -9119
rect 331 -9129 401 -9119
rect 141 -9179 171 -9159
rect 121 -9219 171 -9179
rect 231 -9179 261 -9159
rect 231 -9219 281 -9179
rect 121 -9289 281 -9219
rect 121 -9329 171 -9289
rect 141 -9349 171 -9329
rect 231 -9329 281 -9289
rect 231 -9349 261 -9329
rect 341 -9389 401 -9129
rect 1 -9399 81 -9389
rect 1 -9459 11 -9399
rect 71 -9409 81 -9399
rect 321 -9399 401 -9389
rect 321 -9409 331 -9399
rect 71 -9459 331 -9409
rect 391 -9459 401 -9399
rect 1 -9469 401 -9459
rect 457 -9049 857 -9039
rect 457 -9109 467 -9049
rect 527 -9099 787 -9049
rect 527 -9109 537 -9099
rect 457 -9119 537 -9109
rect 777 -9109 787 -9099
rect 847 -9109 857 -9049
rect 777 -9119 857 -9109
rect 457 -9389 517 -9119
rect 787 -9129 857 -9119
rect 597 -9179 627 -9159
rect 577 -9219 627 -9179
rect 687 -9179 717 -9159
rect 687 -9219 737 -9179
rect 577 -9289 737 -9219
rect 577 -9329 627 -9289
rect 597 -9349 627 -9329
rect 687 -9329 737 -9289
rect 687 -9349 717 -9329
rect 797 -9389 857 -9129
rect 457 -9399 537 -9389
rect 457 -9459 467 -9399
rect 527 -9409 537 -9399
rect 777 -9399 857 -9389
rect 777 -9409 787 -9399
rect 527 -9459 787 -9409
rect 847 -9459 857 -9399
rect 457 -9469 857 -9459
rect 913 -9049 1313 -9039
rect 913 -9109 923 -9049
rect 983 -9099 1243 -9049
rect 983 -9109 993 -9099
rect 913 -9119 993 -9109
rect 1233 -9109 1243 -9099
rect 1303 -9109 1313 -9049
rect 1233 -9119 1313 -9109
rect 913 -9389 973 -9119
rect 1243 -9129 1313 -9119
rect 1053 -9179 1083 -9159
rect 1033 -9219 1083 -9179
rect 1143 -9179 1173 -9159
rect 1143 -9219 1193 -9179
rect 1033 -9289 1193 -9219
rect 1033 -9329 1083 -9289
rect 1053 -9349 1083 -9329
rect 1143 -9329 1193 -9289
rect 1143 -9349 1173 -9329
rect 1253 -9389 1313 -9129
rect 913 -9399 993 -9389
rect 913 -9459 923 -9399
rect 983 -9409 993 -9399
rect 1233 -9399 1313 -9389
rect 1233 -9409 1243 -9399
rect 983 -9459 1243 -9409
rect 1303 -9459 1313 -9399
rect 913 -9469 1313 -9459
rect 1371 -9049 1771 -9039
rect 1371 -9109 1381 -9049
rect 1441 -9099 1701 -9049
rect 1441 -9109 1451 -9099
rect 1371 -9119 1451 -9109
rect 1691 -9109 1701 -9099
rect 1761 -9109 1771 -9049
rect 1691 -9119 1771 -9109
rect 1371 -9389 1431 -9119
rect 1701 -9129 1771 -9119
rect 1511 -9179 1541 -9159
rect 1491 -9219 1541 -9179
rect 1601 -9179 1631 -9159
rect 1601 -9219 1651 -9179
rect 1491 -9289 1651 -9219
rect 1491 -9329 1541 -9289
rect 1511 -9349 1541 -9329
rect 1601 -9329 1651 -9289
rect 1601 -9349 1631 -9329
rect 1711 -9389 1771 -9129
rect 1371 -9399 1451 -9389
rect 1371 -9459 1381 -9399
rect 1441 -9409 1451 -9399
rect 1691 -9399 1771 -9389
rect 1691 -9409 1701 -9399
rect 1441 -9459 1701 -9409
rect 1761 -9459 1771 -9399
rect 1371 -9469 1771 -9459
rect 1827 -9049 2227 -9039
rect 1827 -9109 1837 -9049
rect 1897 -9099 2157 -9049
rect 1897 -9109 1907 -9099
rect 1827 -9119 1907 -9109
rect 2147 -9109 2157 -9099
rect 2217 -9109 2227 -9049
rect 2147 -9119 2227 -9109
rect 1827 -9389 1887 -9119
rect 2157 -9129 2227 -9119
rect 1967 -9179 1997 -9159
rect 1947 -9219 1997 -9179
rect 2057 -9179 2087 -9159
rect 2057 -9219 2107 -9179
rect 1947 -9289 2107 -9219
rect 1947 -9329 1997 -9289
rect 1967 -9349 1997 -9329
rect 2057 -9329 2107 -9289
rect 2057 -9349 2087 -9329
rect 2167 -9389 2227 -9129
rect 1827 -9399 1907 -9389
rect 1827 -9459 1837 -9399
rect 1897 -9409 1907 -9399
rect 2147 -9399 2227 -9389
rect 2147 -9409 2157 -9399
rect 1897 -9459 2157 -9409
rect 2217 -9459 2227 -9399
rect 1827 -9469 2227 -9459
rect 2283 -9049 2683 -9039
rect 2283 -9109 2293 -9049
rect 2353 -9099 2613 -9049
rect 2353 -9109 2363 -9099
rect 2283 -9119 2363 -9109
rect 2603 -9109 2613 -9099
rect 2673 -9109 2683 -9049
rect 2603 -9119 2683 -9109
rect 2283 -9389 2343 -9119
rect 2613 -9129 2683 -9119
rect 2423 -9179 2453 -9159
rect 2403 -9219 2453 -9179
rect 2513 -9179 2543 -9159
rect 2513 -9219 2563 -9179
rect 2403 -9289 2563 -9219
rect 2403 -9329 2453 -9289
rect 2423 -9349 2453 -9329
rect 2513 -9329 2563 -9289
rect 2513 -9349 2543 -9329
rect 2623 -9389 2683 -9129
rect 2283 -9399 2363 -9389
rect 2283 -9459 2293 -9399
rect 2353 -9409 2363 -9399
rect 2603 -9399 2683 -9389
rect 2603 -9409 2613 -9399
rect 2353 -9459 2613 -9409
rect 2673 -9459 2683 -9399
rect 2283 -9469 2683 -9459
rect 2741 -9049 3141 -9039
rect 2741 -9109 2751 -9049
rect 2811 -9099 3071 -9049
rect 2811 -9109 2821 -9099
rect 2741 -9119 2821 -9109
rect 3061 -9109 3071 -9099
rect 3131 -9109 3141 -9049
rect 3061 -9119 3141 -9109
rect 2741 -9389 2801 -9119
rect 3071 -9129 3141 -9119
rect 2881 -9179 2911 -9159
rect 2861 -9219 2911 -9179
rect 2971 -9179 3001 -9159
rect 2971 -9219 3021 -9179
rect 2861 -9289 3021 -9219
rect 2861 -9329 2911 -9289
rect 2881 -9349 2911 -9329
rect 2971 -9329 3021 -9289
rect 2971 -9349 3001 -9329
rect 3081 -9389 3141 -9129
rect 2741 -9399 2821 -9389
rect 2741 -9459 2751 -9399
rect 2811 -9409 2821 -9399
rect 3061 -9399 3141 -9389
rect 3061 -9409 3071 -9399
rect 2811 -9459 3071 -9409
rect 3131 -9459 3141 -9399
rect 2741 -9469 3141 -9459
rect 3197 -9049 3597 -9039
rect 3197 -9109 3207 -9049
rect 3267 -9099 3527 -9049
rect 3267 -9109 3277 -9099
rect 3197 -9119 3277 -9109
rect 3517 -9109 3527 -9099
rect 3587 -9109 3597 -9049
rect 3517 -9119 3597 -9109
rect 3197 -9389 3257 -9119
rect 3527 -9129 3597 -9119
rect 3337 -9179 3367 -9159
rect 3317 -9219 3367 -9179
rect 3427 -9179 3457 -9159
rect 3427 -9219 3477 -9179
rect 3317 -9289 3477 -9219
rect 3317 -9329 3367 -9289
rect 3337 -9349 3367 -9329
rect 3427 -9329 3477 -9289
rect 3427 -9349 3457 -9329
rect 3537 -9389 3597 -9129
rect 3197 -9399 3277 -9389
rect 3197 -9459 3207 -9399
rect 3267 -9409 3277 -9399
rect 3517 -9399 3597 -9389
rect 3517 -9409 3527 -9399
rect 3267 -9459 3527 -9409
rect 3587 -9459 3597 -9399
rect 3197 -9469 3597 -9459
rect 3653 -9049 4053 -9039
rect 3653 -9109 3663 -9049
rect 3723 -9099 3983 -9049
rect 3723 -9109 3733 -9099
rect 3653 -9119 3733 -9109
rect 3973 -9109 3983 -9099
rect 4043 -9109 4053 -9049
rect 3973 -9119 4053 -9109
rect 3653 -9389 3713 -9119
rect 3983 -9129 4053 -9119
rect 3793 -9179 3823 -9159
rect 3773 -9219 3823 -9179
rect 3883 -9179 3913 -9159
rect 3883 -9219 3933 -9179
rect 3773 -9289 3933 -9219
rect 3773 -9329 3823 -9289
rect 3793 -9349 3823 -9329
rect 3883 -9329 3933 -9289
rect 3883 -9349 3913 -9329
rect 3993 -9389 4053 -9129
rect 3653 -9399 3733 -9389
rect 3653 -9459 3663 -9399
rect 3723 -9409 3733 -9399
rect 3973 -9399 4053 -9389
rect 3973 -9409 3983 -9399
rect 3723 -9459 3983 -9409
rect 4043 -9459 4053 -9399
rect 3653 -9469 4053 -9459
rect 4111 -9049 4511 -9039
rect 4111 -9109 4121 -9049
rect 4181 -9099 4441 -9049
rect 4181 -9109 4191 -9099
rect 4111 -9119 4191 -9109
rect 4431 -9109 4441 -9099
rect 4501 -9109 4511 -9049
rect 4431 -9119 4511 -9109
rect 4111 -9389 4171 -9119
rect 4441 -9129 4511 -9119
rect 4251 -9179 4281 -9159
rect 4231 -9219 4281 -9179
rect 4341 -9179 4371 -9159
rect 4341 -9219 4391 -9179
rect 4231 -9289 4391 -9219
rect 4231 -9329 4281 -9289
rect 4251 -9349 4281 -9329
rect 4341 -9329 4391 -9289
rect 4341 -9349 4371 -9329
rect 4451 -9389 4511 -9129
rect 4111 -9399 4191 -9389
rect 4111 -9459 4121 -9399
rect 4181 -9409 4191 -9399
rect 4431 -9399 4511 -9389
rect 4431 -9409 4441 -9399
rect 4181 -9459 4441 -9409
rect 4501 -9459 4511 -9399
rect 4111 -9469 4511 -9459
rect 4567 -9049 4967 -9039
rect 4567 -9109 4577 -9049
rect 4637 -9099 4897 -9049
rect 4637 -9109 4647 -9099
rect 4567 -9119 4647 -9109
rect 4887 -9109 4897 -9099
rect 4957 -9109 4967 -9049
rect 4887 -9119 4967 -9109
rect 4567 -9389 4627 -9119
rect 4897 -9129 4967 -9119
rect 4707 -9179 4737 -9159
rect 4687 -9219 4737 -9179
rect 4797 -9179 4827 -9159
rect 4797 -9219 4847 -9179
rect 4687 -9289 4847 -9219
rect 4687 -9329 4737 -9289
rect 4707 -9349 4737 -9329
rect 4797 -9329 4847 -9289
rect 4797 -9349 4827 -9329
rect 4907 -9389 4967 -9129
rect 4567 -9399 4647 -9389
rect 4567 -9459 4577 -9399
rect 4637 -9409 4647 -9399
rect 4887 -9399 4967 -9389
rect 4887 -9409 4897 -9399
rect 4637 -9459 4897 -9409
rect 4957 -9459 4967 -9399
rect 4567 -9469 4967 -9459
rect 5023 -9049 5423 -9039
rect 5023 -9109 5033 -9049
rect 5093 -9099 5353 -9049
rect 5093 -9109 5103 -9099
rect 5023 -9119 5103 -9109
rect 5343 -9109 5353 -9099
rect 5413 -9109 5423 -9049
rect 5343 -9119 5423 -9109
rect 5023 -9389 5083 -9119
rect 5353 -9129 5423 -9119
rect 5163 -9179 5193 -9159
rect 5143 -9219 5193 -9179
rect 5253 -9179 5283 -9159
rect 5253 -9219 5303 -9179
rect 5143 -9289 5303 -9219
rect 5143 -9329 5193 -9289
rect 5163 -9349 5193 -9329
rect 5253 -9329 5303 -9289
rect 5253 -9349 5283 -9329
rect 5363 -9389 5423 -9129
rect 5023 -9399 5103 -9389
rect 5023 -9459 5033 -9399
rect 5093 -9409 5103 -9399
rect 5343 -9399 5423 -9389
rect 5343 -9409 5353 -9399
rect 5093 -9459 5353 -9409
rect 5413 -9459 5423 -9399
rect 5023 -9469 5423 -9459
rect 5481 -9049 5881 -9039
rect 5481 -9109 5491 -9049
rect 5551 -9099 5811 -9049
rect 5551 -9109 5561 -9099
rect 5481 -9119 5561 -9109
rect 5801 -9109 5811 -9099
rect 5871 -9109 5881 -9049
rect 5801 -9119 5881 -9109
rect 5481 -9389 5541 -9119
rect 5811 -9129 5881 -9119
rect 5621 -9179 5651 -9159
rect 5601 -9219 5651 -9179
rect 5711 -9179 5741 -9159
rect 5711 -9219 5761 -9179
rect 5601 -9289 5761 -9219
rect 5601 -9329 5651 -9289
rect 5621 -9349 5651 -9329
rect 5711 -9329 5761 -9289
rect 5711 -9349 5741 -9329
rect 5821 -9389 5881 -9129
rect 5481 -9399 5561 -9389
rect 5481 -9459 5491 -9399
rect 5551 -9409 5561 -9399
rect 5801 -9399 5881 -9389
rect 5801 -9409 5811 -9399
rect 5551 -9459 5811 -9409
rect 5871 -9459 5881 -9399
rect 5481 -9469 5881 -9459
rect 5937 -9049 6337 -9039
rect 5937 -9109 5947 -9049
rect 6007 -9099 6267 -9049
rect 6007 -9109 6017 -9099
rect 5937 -9119 6017 -9109
rect 6257 -9109 6267 -9099
rect 6327 -9109 6337 -9049
rect 6257 -9119 6337 -9109
rect 5937 -9389 5997 -9119
rect 6267 -9129 6337 -9119
rect 6077 -9179 6107 -9159
rect 6057 -9219 6107 -9179
rect 6167 -9179 6197 -9159
rect 6167 -9219 6217 -9179
rect 6057 -9289 6217 -9219
rect 6057 -9329 6107 -9289
rect 6077 -9349 6107 -9329
rect 6167 -9329 6217 -9289
rect 6167 -9349 6197 -9329
rect 6277 -9389 6337 -9129
rect 5937 -9399 6017 -9389
rect 5937 -9459 5947 -9399
rect 6007 -9409 6017 -9399
rect 6257 -9399 6337 -9389
rect 6257 -9409 6267 -9399
rect 6007 -9459 6267 -9409
rect 6327 -9459 6337 -9399
rect 5937 -9469 6337 -9459
rect 6393 -9049 6793 -9039
rect 6393 -9109 6403 -9049
rect 6463 -9099 6723 -9049
rect 6463 -9109 6473 -9099
rect 6393 -9119 6473 -9109
rect 6713 -9109 6723 -9099
rect 6783 -9109 6793 -9049
rect 6713 -9119 6793 -9109
rect 6393 -9389 6453 -9119
rect 6723 -9129 6793 -9119
rect 6533 -9179 6563 -9159
rect 6513 -9219 6563 -9179
rect 6623 -9179 6653 -9159
rect 6623 -9219 6673 -9179
rect 6513 -9289 6673 -9219
rect 6513 -9329 6563 -9289
rect 6533 -9349 6563 -9329
rect 6623 -9329 6673 -9289
rect 6623 -9349 6653 -9329
rect 6733 -9389 6793 -9129
rect 6393 -9399 6473 -9389
rect 6393 -9459 6403 -9399
rect 6463 -9409 6473 -9399
rect 6713 -9399 6793 -9389
rect 6713 -9409 6723 -9399
rect 6463 -9459 6723 -9409
rect 6783 -9459 6793 -9399
rect 6393 -9469 6793 -9459
rect 6851 -9049 7251 -9039
rect 6851 -9109 6861 -9049
rect 6921 -9099 7181 -9049
rect 6921 -9109 6931 -9099
rect 6851 -9119 6931 -9109
rect 7171 -9109 7181 -9099
rect 7241 -9109 7251 -9049
rect 7171 -9119 7251 -9109
rect 6851 -9389 6911 -9119
rect 7181 -9129 7251 -9119
rect 6991 -9179 7021 -9159
rect 6971 -9219 7021 -9179
rect 7081 -9179 7111 -9159
rect 7081 -9219 7131 -9179
rect 6971 -9289 7131 -9219
rect 6971 -9329 7021 -9289
rect 6991 -9349 7021 -9329
rect 7081 -9329 7131 -9289
rect 7081 -9349 7111 -9329
rect 7191 -9389 7251 -9129
rect 6851 -9399 6931 -9389
rect 6851 -9459 6861 -9399
rect 6921 -9409 6931 -9399
rect 7171 -9399 7251 -9389
rect 7171 -9409 7181 -9399
rect 6921 -9459 7181 -9409
rect 7241 -9459 7251 -9399
rect 6851 -9469 7251 -9459
rect 7307 -9049 7707 -9039
rect 7307 -9109 7317 -9049
rect 7377 -9099 7637 -9049
rect 7377 -9109 7387 -9099
rect 7307 -9119 7387 -9109
rect 7627 -9109 7637 -9099
rect 7697 -9109 7707 -9049
rect 7627 -9119 7707 -9109
rect 7307 -9389 7367 -9119
rect 7637 -9129 7707 -9119
rect 7447 -9179 7477 -9159
rect 7427 -9219 7477 -9179
rect 7537 -9179 7567 -9159
rect 7537 -9219 7587 -9179
rect 7427 -9289 7587 -9219
rect 7427 -9329 7477 -9289
rect 7447 -9349 7477 -9329
rect 7537 -9329 7587 -9289
rect 7537 -9349 7567 -9329
rect 7647 -9389 7707 -9129
rect 7307 -9399 7387 -9389
rect 7307 -9459 7317 -9399
rect 7377 -9409 7387 -9399
rect 7627 -9399 7707 -9389
rect 7627 -9409 7637 -9399
rect 7377 -9459 7637 -9409
rect 7697 -9459 7707 -9399
rect 7307 -9469 7707 -9459
rect 7763 -9049 8163 -9039
rect 7763 -9109 7773 -9049
rect 7833 -9099 8093 -9049
rect 7833 -9109 7843 -9099
rect 7763 -9119 7843 -9109
rect 8083 -9109 8093 -9099
rect 8153 -9109 8163 -9049
rect 8083 -9119 8163 -9109
rect 7763 -9389 7823 -9119
rect 8093 -9129 8163 -9119
rect 7903 -9179 7933 -9159
rect 7883 -9219 7933 -9179
rect 7993 -9179 8023 -9159
rect 7993 -9219 8043 -9179
rect 7883 -9289 8043 -9219
rect 7883 -9329 7933 -9289
rect 7903 -9349 7933 -9329
rect 7993 -9329 8043 -9289
rect 7993 -9349 8023 -9329
rect 8103 -9389 8163 -9129
rect 7763 -9399 7843 -9389
rect 7763 -9459 7773 -9399
rect 7833 -9409 7843 -9399
rect 8083 -9399 8163 -9389
rect 8083 -9409 8093 -9399
rect 7833 -9459 8093 -9409
rect 8153 -9459 8163 -9399
rect 7763 -9469 8163 -9459
rect 8237 -9049 8637 -9039
rect 8237 -9109 8247 -9049
rect 8307 -9099 8567 -9049
rect 8307 -9109 8317 -9099
rect 8237 -9119 8317 -9109
rect 8557 -9109 8567 -9099
rect 8627 -9109 8637 -9049
rect 8557 -9119 8637 -9109
rect 8237 -9389 8297 -9119
rect 8567 -9129 8637 -9119
rect 8377 -9179 8407 -9159
rect 8357 -9219 8407 -9179
rect 8467 -9179 8497 -9159
rect 8467 -9219 8517 -9179
rect 8357 -9289 8517 -9219
rect 8357 -9329 8407 -9289
rect 8377 -9349 8407 -9329
rect 8467 -9329 8517 -9289
rect 8467 -9349 8497 -9329
rect 8577 -9389 8637 -9129
rect 8237 -9399 8317 -9389
rect 8237 -9459 8247 -9399
rect 8307 -9409 8317 -9399
rect 8557 -9399 8637 -9389
rect 8557 -9409 8567 -9399
rect 8307 -9459 8567 -9409
rect 8627 -9459 8637 -9399
rect 8237 -9469 8637 -9459
rect 8693 -9049 9093 -9039
rect 8693 -9109 8703 -9049
rect 8763 -9099 9023 -9049
rect 8763 -9109 8773 -9099
rect 8693 -9119 8773 -9109
rect 9013 -9109 9023 -9099
rect 9083 -9109 9093 -9049
rect 9013 -9119 9093 -9109
rect 8693 -9389 8753 -9119
rect 9023 -9129 9093 -9119
rect 8833 -9179 8863 -9159
rect 8813 -9219 8863 -9179
rect 8923 -9179 8953 -9159
rect 8923 -9219 8973 -9179
rect 8813 -9289 8973 -9219
rect 8813 -9329 8863 -9289
rect 8833 -9349 8863 -9329
rect 8923 -9329 8973 -9289
rect 8923 -9349 8953 -9329
rect 9033 -9389 9093 -9129
rect 8693 -9399 8773 -9389
rect 8693 -9459 8703 -9399
rect 8763 -9409 8773 -9399
rect 9013 -9399 9093 -9389
rect 9013 -9409 9023 -9399
rect 8763 -9459 9023 -9409
rect 9083 -9459 9093 -9399
rect 8693 -9469 9093 -9459
rect 9151 -9049 9551 -9039
rect 9151 -9109 9161 -9049
rect 9221 -9099 9481 -9049
rect 9221 -9109 9231 -9099
rect 9151 -9119 9231 -9109
rect 9471 -9109 9481 -9099
rect 9541 -9109 9551 -9049
rect 9471 -9119 9551 -9109
rect 9151 -9389 9211 -9119
rect 9481 -9129 9551 -9119
rect 9291 -9179 9321 -9159
rect 9271 -9219 9321 -9179
rect 9381 -9179 9411 -9159
rect 9381 -9219 9431 -9179
rect 9271 -9289 9431 -9219
rect 9271 -9329 9321 -9289
rect 9291 -9349 9321 -9329
rect 9381 -9329 9431 -9289
rect 9381 -9349 9411 -9329
rect 9491 -9389 9551 -9129
rect 9151 -9399 9231 -9389
rect 9151 -9459 9161 -9399
rect 9221 -9409 9231 -9399
rect 9471 -9399 9551 -9389
rect 9471 -9409 9481 -9399
rect 9221 -9459 9481 -9409
rect 9541 -9459 9551 -9399
rect 9151 -9469 9551 -9459
rect 9607 -9049 10007 -9039
rect 9607 -9109 9617 -9049
rect 9677 -9099 9937 -9049
rect 9677 -9109 9687 -9099
rect 9607 -9119 9687 -9109
rect 9927 -9109 9937 -9099
rect 9997 -9109 10007 -9049
rect 9927 -9119 10007 -9109
rect 9607 -9389 9667 -9119
rect 9937 -9129 10007 -9119
rect 9747 -9179 9777 -9159
rect 9727 -9219 9777 -9179
rect 9837 -9179 9867 -9159
rect 9837 -9219 9887 -9179
rect 9727 -9289 9887 -9219
rect 9727 -9329 9777 -9289
rect 9747 -9349 9777 -9329
rect 9837 -9329 9887 -9289
rect 9837 -9349 9867 -9329
rect 9947 -9389 10007 -9129
rect 9607 -9399 9687 -9389
rect 9607 -9459 9617 -9399
rect 9677 -9409 9687 -9399
rect 9927 -9399 10007 -9389
rect 9927 -9409 9937 -9399
rect 9677 -9459 9937 -9409
rect 9997 -9459 10007 -9399
rect 9607 -9469 10007 -9459
rect 10063 -9049 10463 -9039
rect 10063 -9109 10073 -9049
rect 10133 -9099 10393 -9049
rect 10133 -9109 10143 -9099
rect 10063 -9119 10143 -9109
rect 10383 -9109 10393 -9099
rect 10453 -9109 10463 -9049
rect 10383 -9119 10463 -9109
rect 10063 -9389 10123 -9119
rect 10393 -9129 10463 -9119
rect 10203 -9179 10233 -9159
rect 10183 -9219 10233 -9179
rect 10293 -9179 10323 -9159
rect 10293 -9219 10343 -9179
rect 10183 -9289 10343 -9219
rect 10183 -9329 10233 -9289
rect 10203 -9349 10233 -9329
rect 10293 -9329 10343 -9289
rect 10293 -9349 10323 -9329
rect 10403 -9389 10463 -9129
rect 10063 -9399 10143 -9389
rect 10063 -9459 10073 -9399
rect 10133 -9409 10143 -9399
rect 10383 -9399 10463 -9389
rect 10383 -9409 10393 -9399
rect 10133 -9459 10393 -9409
rect 10453 -9459 10463 -9399
rect 10063 -9469 10463 -9459
rect 10521 -9049 10921 -9039
rect 10521 -9109 10531 -9049
rect 10591 -9099 10851 -9049
rect 10591 -9109 10601 -9099
rect 10521 -9119 10601 -9109
rect 10841 -9109 10851 -9099
rect 10911 -9109 10921 -9049
rect 10841 -9119 10921 -9109
rect 10521 -9389 10581 -9119
rect 10851 -9129 10921 -9119
rect 10661 -9179 10691 -9159
rect 10641 -9219 10691 -9179
rect 10751 -9179 10781 -9159
rect 10751 -9219 10801 -9179
rect 10641 -9289 10801 -9219
rect 10641 -9329 10691 -9289
rect 10661 -9349 10691 -9329
rect 10751 -9329 10801 -9289
rect 10751 -9349 10781 -9329
rect 10861 -9389 10921 -9129
rect 10521 -9399 10601 -9389
rect 10521 -9459 10531 -9399
rect 10591 -9409 10601 -9399
rect 10841 -9399 10921 -9389
rect 10841 -9409 10851 -9399
rect 10591 -9459 10851 -9409
rect 10911 -9459 10921 -9399
rect 10521 -9469 10921 -9459
rect 10977 -9049 11377 -9039
rect 10977 -9109 10987 -9049
rect 11047 -9099 11307 -9049
rect 11047 -9109 11057 -9099
rect 10977 -9119 11057 -9109
rect 11297 -9109 11307 -9099
rect 11367 -9109 11377 -9049
rect 11297 -9119 11377 -9109
rect 10977 -9389 11037 -9119
rect 11307 -9129 11377 -9119
rect 11117 -9179 11147 -9159
rect 11097 -9219 11147 -9179
rect 11207 -9179 11237 -9159
rect 11207 -9219 11257 -9179
rect 11097 -9289 11257 -9219
rect 11097 -9329 11147 -9289
rect 11117 -9349 11147 -9329
rect 11207 -9329 11257 -9289
rect 11207 -9349 11237 -9329
rect 11317 -9389 11377 -9129
rect 10977 -9399 11057 -9389
rect 10977 -9459 10987 -9399
rect 11047 -9409 11057 -9399
rect 11297 -9399 11377 -9389
rect 11297 -9409 11307 -9399
rect 11047 -9459 11307 -9409
rect 11367 -9459 11377 -9399
rect 10977 -9469 11377 -9459
rect 11433 -9049 11833 -9039
rect 11433 -9109 11443 -9049
rect 11503 -9099 11763 -9049
rect 11503 -9109 11513 -9099
rect 11433 -9119 11513 -9109
rect 11753 -9109 11763 -9099
rect 11823 -9109 11833 -9049
rect 11753 -9119 11833 -9109
rect 11433 -9389 11493 -9119
rect 11763 -9129 11833 -9119
rect 11573 -9179 11603 -9159
rect 11553 -9219 11603 -9179
rect 11663 -9179 11693 -9159
rect 11663 -9219 11713 -9179
rect 11553 -9289 11713 -9219
rect 11553 -9329 11603 -9289
rect 11573 -9349 11603 -9329
rect 11663 -9329 11713 -9289
rect 11663 -9349 11693 -9329
rect 11773 -9389 11833 -9129
rect 11433 -9399 11513 -9389
rect 11433 -9459 11443 -9399
rect 11503 -9409 11513 -9399
rect 11753 -9399 11833 -9389
rect 11753 -9409 11763 -9399
rect 11503 -9459 11763 -9409
rect 11823 -9459 11833 -9399
rect 11433 -9469 11833 -9459
rect 11891 -9049 12291 -9039
rect 11891 -9109 11901 -9049
rect 11961 -9099 12221 -9049
rect 11961 -9109 11971 -9099
rect 11891 -9119 11971 -9109
rect 12211 -9109 12221 -9099
rect 12281 -9109 12291 -9049
rect 12211 -9119 12291 -9109
rect 11891 -9389 11951 -9119
rect 12221 -9129 12291 -9119
rect 12031 -9179 12061 -9159
rect 12011 -9219 12061 -9179
rect 12121 -9179 12151 -9159
rect 12121 -9219 12171 -9179
rect 12011 -9289 12171 -9219
rect 12011 -9329 12061 -9289
rect 12031 -9349 12061 -9329
rect 12121 -9329 12171 -9289
rect 12121 -9349 12151 -9329
rect 12231 -9389 12291 -9129
rect 11891 -9399 11971 -9389
rect 11891 -9459 11901 -9399
rect 11961 -9409 11971 -9399
rect 12211 -9399 12291 -9389
rect 12211 -9409 12221 -9399
rect 11961 -9459 12221 -9409
rect 12281 -9459 12291 -9399
rect 11891 -9469 12291 -9459
rect 12347 -9049 12747 -9039
rect 12347 -9109 12357 -9049
rect 12417 -9099 12677 -9049
rect 12417 -9109 12427 -9099
rect 12347 -9119 12427 -9109
rect 12667 -9109 12677 -9099
rect 12737 -9109 12747 -9049
rect 12667 -9119 12747 -9109
rect 12347 -9389 12407 -9119
rect 12677 -9129 12747 -9119
rect 12487 -9179 12517 -9159
rect 12467 -9219 12517 -9179
rect 12577 -9179 12607 -9159
rect 12577 -9219 12627 -9179
rect 12467 -9289 12627 -9219
rect 12467 -9329 12517 -9289
rect 12487 -9349 12517 -9329
rect 12577 -9329 12627 -9289
rect 12577 -9349 12607 -9329
rect 12687 -9389 12747 -9129
rect 12347 -9399 12427 -9389
rect 12347 -9459 12357 -9399
rect 12417 -9409 12427 -9399
rect 12667 -9399 12747 -9389
rect 12667 -9409 12677 -9399
rect 12417 -9459 12677 -9409
rect 12737 -9459 12747 -9399
rect 12347 -9469 12747 -9459
rect 12803 -9049 13203 -9039
rect 12803 -9109 12813 -9049
rect 12873 -9099 13133 -9049
rect 12873 -9109 12883 -9099
rect 12803 -9119 12883 -9109
rect 13123 -9109 13133 -9099
rect 13193 -9109 13203 -9049
rect 13123 -9119 13203 -9109
rect 12803 -9389 12863 -9119
rect 13133 -9129 13203 -9119
rect 12943 -9179 12973 -9159
rect 12923 -9219 12973 -9179
rect 13033 -9179 13063 -9159
rect 13033 -9219 13083 -9179
rect 12923 -9289 13083 -9219
rect 12923 -9329 12973 -9289
rect 12943 -9349 12973 -9329
rect 13033 -9329 13083 -9289
rect 13033 -9349 13063 -9329
rect 13143 -9389 13203 -9129
rect 12803 -9399 12883 -9389
rect 12803 -9459 12813 -9399
rect 12873 -9409 12883 -9399
rect 13123 -9399 13203 -9389
rect 13123 -9409 13133 -9399
rect 12873 -9459 13133 -9409
rect 13193 -9459 13203 -9399
rect 12803 -9469 13203 -9459
rect 13261 -9049 13661 -9039
rect 13261 -9109 13271 -9049
rect 13331 -9099 13591 -9049
rect 13331 -9109 13341 -9099
rect 13261 -9119 13341 -9109
rect 13581 -9109 13591 -9099
rect 13651 -9109 13661 -9049
rect 13581 -9119 13661 -9109
rect 13261 -9389 13321 -9119
rect 13591 -9129 13661 -9119
rect 13401 -9179 13431 -9159
rect 13381 -9219 13431 -9179
rect 13491 -9179 13521 -9159
rect 13491 -9219 13541 -9179
rect 13381 -9289 13541 -9219
rect 13381 -9329 13431 -9289
rect 13401 -9349 13431 -9329
rect 13491 -9329 13541 -9289
rect 13491 -9349 13521 -9329
rect 13601 -9389 13661 -9129
rect 13261 -9399 13341 -9389
rect 13261 -9459 13271 -9399
rect 13331 -9409 13341 -9399
rect 13581 -9399 13661 -9389
rect 13581 -9409 13591 -9399
rect 13331 -9459 13591 -9409
rect 13651 -9459 13661 -9399
rect 13261 -9469 13661 -9459
rect 13717 -9049 14117 -9039
rect 13717 -9109 13727 -9049
rect 13787 -9099 14047 -9049
rect 13787 -9109 13797 -9099
rect 13717 -9119 13797 -9109
rect 14037 -9109 14047 -9099
rect 14107 -9109 14117 -9049
rect 14037 -9119 14117 -9109
rect 13717 -9389 13777 -9119
rect 14047 -9129 14117 -9119
rect 13857 -9179 13887 -9159
rect 13837 -9219 13887 -9179
rect 13947 -9179 13977 -9159
rect 13947 -9219 13997 -9179
rect 13837 -9289 13997 -9219
rect 13837 -9329 13887 -9289
rect 13857 -9349 13887 -9329
rect 13947 -9329 13997 -9289
rect 13947 -9349 13977 -9329
rect 14057 -9389 14117 -9129
rect 13717 -9399 13797 -9389
rect 13717 -9459 13727 -9399
rect 13787 -9409 13797 -9399
rect 14037 -9399 14117 -9389
rect 14037 -9409 14047 -9399
rect 13787 -9459 14047 -9409
rect 14107 -9459 14117 -9399
rect 13717 -9469 14117 -9459
rect 14173 -9049 14573 -9039
rect 14173 -9109 14183 -9049
rect 14243 -9099 14503 -9049
rect 14243 -9109 14253 -9099
rect 14173 -9119 14253 -9109
rect 14493 -9109 14503 -9099
rect 14563 -9109 14573 -9049
rect 14493 -9119 14573 -9109
rect 14173 -9389 14233 -9119
rect 14503 -9129 14573 -9119
rect 14313 -9179 14343 -9159
rect 14293 -9219 14343 -9179
rect 14403 -9179 14433 -9159
rect 14403 -9219 14453 -9179
rect 14293 -9289 14453 -9219
rect 14293 -9329 14343 -9289
rect 14313 -9349 14343 -9329
rect 14403 -9329 14453 -9289
rect 14403 -9349 14433 -9329
rect 14513 -9389 14573 -9129
rect 14173 -9399 14253 -9389
rect 14173 -9459 14183 -9399
rect 14243 -9409 14253 -9399
rect 14493 -9399 14573 -9389
rect 14493 -9409 14503 -9399
rect 14243 -9459 14503 -9409
rect 14563 -9459 14573 -9399
rect 14173 -9469 14573 -9459
rect 14631 -9049 15031 -9039
rect 14631 -9109 14641 -9049
rect 14701 -9099 14961 -9049
rect 14701 -9109 14711 -9099
rect 14631 -9119 14711 -9109
rect 14951 -9109 14961 -9099
rect 15021 -9109 15031 -9049
rect 14951 -9119 15031 -9109
rect 14631 -9389 14691 -9119
rect 14961 -9129 15031 -9119
rect 14771 -9179 14801 -9159
rect 14751 -9219 14801 -9179
rect 14861 -9179 14891 -9159
rect 14861 -9219 14911 -9179
rect 14751 -9289 14911 -9219
rect 14751 -9329 14801 -9289
rect 14771 -9349 14801 -9329
rect 14861 -9329 14911 -9289
rect 14861 -9349 14891 -9329
rect 14971 -9389 15031 -9129
rect 14631 -9399 14711 -9389
rect 14631 -9459 14641 -9399
rect 14701 -9409 14711 -9399
rect 14951 -9399 15031 -9389
rect 14951 -9409 14961 -9399
rect 14701 -9459 14961 -9409
rect 15021 -9459 15031 -9399
rect 14631 -9469 15031 -9459
rect 15087 -9049 15487 -9039
rect 15087 -9109 15097 -9049
rect 15157 -9099 15417 -9049
rect 15157 -9109 15167 -9099
rect 15087 -9119 15167 -9109
rect 15407 -9109 15417 -9099
rect 15477 -9109 15487 -9049
rect 15407 -9119 15487 -9109
rect 15087 -9389 15147 -9119
rect 15417 -9129 15487 -9119
rect 15227 -9179 15257 -9159
rect 15207 -9219 15257 -9179
rect 15317 -9179 15347 -9159
rect 15317 -9219 15367 -9179
rect 15207 -9289 15367 -9219
rect 15207 -9329 15257 -9289
rect 15227 -9349 15257 -9329
rect 15317 -9329 15367 -9289
rect 15317 -9349 15347 -9329
rect 15427 -9389 15487 -9129
rect 15087 -9399 15167 -9389
rect 15087 -9459 15097 -9399
rect 15157 -9409 15167 -9399
rect 15407 -9399 15487 -9389
rect 15407 -9409 15417 -9399
rect 15157 -9459 15417 -9409
rect 15477 -9459 15487 -9399
rect 15087 -9469 15487 -9459
rect 1 -9541 401 -9531
rect 1 -9601 11 -9541
rect 71 -9591 331 -9541
rect 71 -9601 81 -9591
rect 1 -9611 81 -9601
rect 321 -9601 331 -9591
rect 391 -9601 401 -9541
rect 321 -9611 401 -9601
rect 1 -9881 61 -9611
rect 331 -9621 401 -9611
rect 141 -9671 171 -9651
rect 121 -9711 171 -9671
rect 231 -9671 261 -9651
rect 231 -9711 281 -9671
rect 121 -9781 281 -9711
rect 121 -9821 171 -9781
rect 141 -9841 171 -9821
rect 231 -9821 281 -9781
rect 231 -9841 261 -9821
rect 341 -9881 401 -9621
rect 1 -9891 81 -9881
rect 1 -9951 11 -9891
rect 71 -9901 81 -9891
rect 321 -9891 401 -9881
rect 321 -9901 331 -9891
rect 71 -9951 331 -9901
rect 391 -9951 401 -9891
rect 1 -9961 401 -9951
rect 457 -9541 857 -9531
rect 457 -9601 467 -9541
rect 527 -9591 787 -9541
rect 527 -9601 537 -9591
rect 457 -9611 537 -9601
rect 777 -9601 787 -9591
rect 847 -9601 857 -9541
rect 777 -9611 857 -9601
rect 457 -9881 517 -9611
rect 787 -9621 857 -9611
rect 597 -9671 627 -9651
rect 577 -9711 627 -9671
rect 687 -9671 717 -9651
rect 687 -9711 737 -9671
rect 577 -9781 737 -9711
rect 577 -9821 627 -9781
rect 597 -9841 627 -9821
rect 687 -9821 737 -9781
rect 687 -9841 717 -9821
rect 797 -9881 857 -9621
rect 457 -9891 537 -9881
rect 457 -9951 467 -9891
rect 527 -9901 537 -9891
rect 777 -9891 857 -9881
rect 777 -9901 787 -9891
rect 527 -9951 787 -9901
rect 847 -9951 857 -9891
rect 457 -9961 857 -9951
rect 913 -9541 1313 -9531
rect 913 -9601 923 -9541
rect 983 -9591 1243 -9541
rect 983 -9601 993 -9591
rect 913 -9611 993 -9601
rect 1233 -9601 1243 -9591
rect 1303 -9601 1313 -9541
rect 1233 -9611 1313 -9601
rect 913 -9881 973 -9611
rect 1243 -9621 1313 -9611
rect 1053 -9671 1083 -9651
rect 1033 -9711 1083 -9671
rect 1143 -9671 1173 -9651
rect 1143 -9711 1193 -9671
rect 1033 -9781 1193 -9711
rect 1033 -9821 1083 -9781
rect 1053 -9841 1083 -9821
rect 1143 -9821 1193 -9781
rect 1143 -9841 1173 -9821
rect 1253 -9881 1313 -9621
rect 913 -9891 993 -9881
rect 913 -9951 923 -9891
rect 983 -9901 993 -9891
rect 1233 -9891 1313 -9881
rect 1233 -9901 1243 -9891
rect 983 -9951 1243 -9901
rect 1303 -9951 1313 -9891
rect 913 -9961 1313 -9951
rect 1371 -9541 1771 -9531
rect 1371 -9601 1381 -9541
rect 1441 -9591 1701 -9541
rect 1441 -9601 1451 -9591
rect 1371 -9611 1451 -9601
rect 1691 -9601 1701 -9591
rect 1761 -9601 1771 -9541
rect 1691 -9611 1771 -9601
rect 1371 -9881 1431 -9611
rect 1701 -9621 1771 -9611
rect 1511 -9671 1541 -9651
rect 1491 -9711 1541 -9671
rect 1601 -9671 1631 -9651
rect 1601 -9711 1651 -9671
rect 1491 -9781 1651 -9711
rect 1491 -9821 1541 -9781
rect 1511 -9841 1541 -9821
rect 1601 -9821 1651 -9781
rect 1601 -9841 1631 -9821
rect 1711 -9881 1771 -9621
rect 1371 -9891 1451 -9881
rect 1371 -9951 1381 -9891
rect 1441 -9901 1451 -9891
rect 1691 -9891 1771 -9881
rect 1691 -9901 1701 -9891
rect 1441 -9951 1701 -9901
rect 1761 -9951 1771 -9891
rect 1371 -9961 1771 -9951
rect 1827 -9541 2227 -9531
rect 1827 -9601 1837 -9541
rect 1897 -9591 2157 -9541
rect 1897 -9601 1907 -9591
rect 1827 -9611 1907 -9601
rect 2147 -9601 2157 -9591
rect 2217 -9601 2227 -9541
rect 2147 -9611 2227 -9601
rect 1827 -9881 1887 -9611
rect 2157 -9621 2227 -9611
rect 1967 -9671 1997 -9651
rect 1947 -9711 1997 -9671
rect 2057 -9671 2087 -9651
rect 2057 -9711 2107 -9671
rect 1947 -9781 2107 -9711
rect 1947 -9821 1997 -9781
rect 1967 -9841 1997 -9821
rect 2057 -9821 2107 -9781
rect 2057 -9841 2087 -9821
rect 2167 -9881 2227 -9621
rect 1827 -9891 1907 -9881
rect 1827 -9951 1837 -9891
rect 1897 -9901 1907 -9891
rect 2147 -9891 2227 -9881
rect 2147 -9901 2157 -9891
rect 1897 -9951 2157 -9901
rect 2217 -9951 2227 -9891
rect 1827 -9961 2227 -9951
rect 2283 -9541 2683 -9531
rect 2283 -9601 2293 -9541
rect 2353 -9591 2613 -9541
rect 2353 -9601 2363 -9591
rect 2283 -9611 2363 -9601
rect 2603 -9601 2613 -9591
rect 2673 -9601 2683 -9541
rect 2603 -9611 2683 -9601
rect 2283 -9881 2343 -9611
rect 2613 -9621 2683 -9611
rect 2423 -9671 2453 -9651
rect 2403 -9711 2453 -9671
rect 2513 -9671 2543 -9651
rect 2513 -9711 2563 -9671
rect 2403 -9781 2563 -9711
rect 2403 -9821 2453 -9781
rect 2423 -9841 2453 -9821
rect 2513 -9821 2563 -9781
rect 2513 -9841 2543 -9821
rect 2623 -9881 2683 -9621
rect 2283 -9891 2363 -9881
rect 2283 -9951 2293 -9891
rect 2353 -9901 2363 -9891
rect 2603 -9891 2683 -9881
rect 2603 -9901 2613 -9891
rect 2353 -9951 2613 -9901
rect 2673 -9951 2683 -9891
rect 2283 -9961 2683 -9951
rect 2741 -9541 3141 -9531
rect 2741 -9601 2751 -9541
rect 2811 -9591 3071 -9541
rect 2811 -9601 2821 -9591
rect 2741 -9611 2821 -9601
rect 3061 -9601 3071 -9591
rect 3131 -9601 3141 -9541
rect 3061 -9611 3141 -9601
rect 2741 -9881 2801 -9611
rect 3071 -9621 3141 -9611
rect 2881 -9671 2911 -9651
rect 2861 -9711 2911 -9671
rect 2971 -9671 3001 -9651
rect 2971 -9711 3021 -9671
rect 2861 -9781 3021 -9711
rect 2861 -9821 2911 -9781
rect 2881 -9841 2911 -9821
rect 2971 -9821 3021 -9781
rect 2971 -9841 3001 -9821
rect 3081 -9881 3141 -9621
rect 2741 -9891 2821 -9881
rect 2741 -9951 2751 -9891
rect 2811 -9901 2821 -9891
rect 3061 -9891 3141 -9881
rect 3061 -9901 3071 -9891
rect 2811 -9951 3071 -9901
rect 3131 -9951 3141 -9891
rect 2741 -9961 3141 -9951
rect 3197 -9541 3597 -9531
rect 3197 -9601 3207 -9541
rect 3267 -9591 3527 -9541
rect 3267 -9601 3277 -9591
rect 3197 -9611 3277 -9601
rect 3517 -9601 3527 -9591
rect 3587 -9601 3597 -9541
rect 3517 -9611 3597 -9601
rect 3197 -9881 3257 -9611
rect 3527 -9621 3597 -9611
rect 3337 -9671 3367 -9651
rect 3317 -9711 3367 -9671
rect 3427 -9671 3457 -9651
rect 3427 -9711 3477 -9671
rect 3317 -9781 3477 -9711
rect 3317 -9821 3367 -9781
rect 3337 -9841 3367 -9821
rect 3427 -9821 3477 -9781
rect 3427 -9841 3457 -9821
rect 3537 -9881 3597 -9621
rect 3197 -9891 3277 -9881
rect 3197 -9951 3207 -9891
rect 3267 -9901 3277 -9891
rect 3517 -9891 3597 -9881
rect 3517 -9901 3527 -9891
rect 3267 -9951 3527 -9901
rect 3587 -9951 3597 -9891
rect 3197 -9961 3597 -9951
rect 3653 -9541 4053 -9531
rect 3653 -9601 3663 -9541
rect 3723 -9591 3983 -9541
rect 3723 -9601 3733 -9591
rect 3653 -9611 3733 -9601
rect 3973 -9601 3983 -9591
rect 4043 -9601 4053 -9541
rect 3973 -9611 4053 -9601
rect 3653 -9881 3713 -9611
rect 3983 -9621 4053 -9611
rect 3793 -9671 3823 -9651
rect 3773 -9711 3823 -9671
rect 3883 -9671 3913 -9651
rect 3883 -9711 3933 -9671
rect 3773 -9781 3933 -9711
rect 3773 -9821 3823 -9781
rect 3793 -9841 3823 -9821
rect 3883 -9821 3933 -9781
rect 3883 -9841 3913 -9821
rect 3993 -9881 4053 -9621
rect 3653 -9891 3733 -9881
rect 3653 -9951 3663 -9891
rect 3723 -9901 3733 -9891
rect 3973 -9891 4053 -9881
rect 3973 -9901 3983 -9891
rect 3723 -9951 3983 -9901
rect 4043 -9951 4053 -9891
rect 3653 -9961 4053 -9951
rect 4111 -9541 4511 -9531
rect 4111 -9601 4121 -9541
rect 4181 -9591 4441 -9541
rect 4181 -9601 4191 -9591
rect 4111 -9611 4191 -9601
rect 4431 -9601 4441 -9591
rect 4501 -9601 4511 -9541
rect 4431 -9611 4511 -9601
rect 4111 -9881 4171 -9611
rect 4441 -9621 4511 -9611
rect 4251 -9671 4281 -9651
rect 4231 -9711 4281 -9671
rect 4341 -9671 4371 -9651
rect 4341 -9711 4391 -9671
rect 4231 -9781 4391 -9711
rect 4231 -9821 4281 -9781
rect 4251 -9841 4281 -9821
rect 4341 -9821 4391 -9781
rect 4341 -9841 4371 -9821
rect 4451 -9881 4511 -9621
rect 4111 -9891 4191 -9881
rect 4111 -9951 4121 -9891
rect 4181 -9901 4191 -9891
rect 4431 -9891 4511 -9881
rect 4431 -9901 4441 -9891
rect 4181 -9951 4441 -9901
rect 4501 -9951 4511 -9891
rect 4111 -9961 4511 -9951
rect 4567 -9541 4967 -9531
rect 4567 -9601 4577 -9541
rect 4637 -9591 4897 -9541
rect 4637 -9601 4647 -9591
rect 4567 -9611 4647 -9601
rect 4887 -9601 4897 -9591
rect 4957 -9601 4967 -9541
rect 4887 -9611 4967 -9601
rect 4567 -9881 4627 -9611
rect 4897 -9621 4967 -9611
rect 4707 -9671 4737 -9651
rect 4687 -9711 4737 -9671
rect 4797 -9671 4827 -9651
rect 4797 -9711 4847 -9671
rect 4687 -9781 4847 -9711
rect 4687 -9821 4737 -9781
rect 4707 -9841 4737 -9821
rect 4797 -9821 4847 -9781
rect 4797 -9841 4827 -9821
rect 4907 -9881 4967 -9621
rect 4567 -9891 4647 -9881
rect 4567 -9951 4577 -9891
rect 4637 -9901 4647 -9891
rect 4887 -9891 4967 -9881
rect 4887 -9901 4897 -9891
rect 4637 -9951 4897 -9901
rect 4957 -9951 4967 -9891
rect 4567 -9961 4967 -9951
rect 5023 -9541 5423 -9531
rect 5023 -9601 5033 -9541
rect 5093 -9591 5353 -9541
rect 5093 -9601 5103 -9591
rect 5023 -9611 5103 -9601
rect 5343 -9601 5353 -9591
rect 5413 -9601 5423 -9541
rect 5343 -9611 5423 -9601
rect 5023 -9881 5083 -9611
rect 5353 -9621 5423 -9611
rect 5163 -9671 5193 -9651
rect 5143 -9711 5193 -9671
rect 5253 -9671 5283 -9651
rect 5253 -9711 5303 -9671
rect 5143 -9781 5303 -9711
rect 5143 -9821 5193 -9781
rect 5163 -9841 5193 -9821
rect 5253 -9821 5303 -9781
rect 5253 -9841 5283 -9821
rect 5363 -9881 5423 -9621
rect 5023 -9891 5103 -9881
rect 5023 -9951 5033 -9891
rect 5093 -9901 5103 -9891
rect 5343 -9891 5423 -9881
rect 5343 -9901 5353 -9891
rect 5093 -9951 5353 -9901
rect 5413 -9951 5423 -9891
rect 5023 -9961 5423 -9951
rect 5481 -9541 5881 -9531
rect 5481 -9601 5491 -9541
rect 5551 -9591 5811 -9541
rect 5551 -9601 5561 -9591
rect 5481 -9611 5561 -9601
rect 5801 -9601 5811 -9591
rect 5871 -9601 5881 -9541
rect 5801 -9611 5881 -9601
rect 5481 -9881 5541 -9611
rect 5811 -9621 5881 -9611
rect 5621 -9671 5651 -9651
rect 5601 -9711 5651 -9671
rect 5711 -9671 5741 -9651
rect 5711 -9711 5761 -9671
rect 5601 -9781 5761 -9711
rect 5601 -9821 5651 -9781
rect 5621 -9841 5651 -9821
rect 5711 -9821 5761 -9781
rect 5711 -9841 5741 -9821
rect 5821 -9881 5881 -9621
rect 5481 -9891 5561 -9881
rect 5481 -9951 5491 -9891
rect 5551 -9901 5561 -9891
rect 5801 -9891 5881 -9881
rect 5801 -9901 5811 -9891
rect 5551 -9951 5811 -9901
rect 5871 -9951 5881 -9891
rect 5481 -9961 5881 -9951
rect 5937 -9541 6337 -9531
rect 5937 -9601 5947 -9541
rect 6007 -9591 6267 -9541
rect 6007 -9601 6017 -9591
rect 5937 -9611 6017 -9601
rect 6257 -9601 6267 -9591
rect 6327 -9601 6337 -9541
rect 6257 -9611 6337 -9601
rect 5937 -9881 5997 -9611
rect 6267 -9621 6337 -9611
rect 6077 -9671 6107 -9651
rect 6057 -9711 6107 -9671
rect 6167 -9671 6197 -9651
rect 6167 -9711 6217 -9671
rect 6057 -9781 6217 -9711
rect 6057 -9821 6107 -9781
rect 6077 -9841 6107 -9821
rect 6167 -9821 6217 -9781
rect 6167 -9841 6197 -9821
rect 6277 -9881 6337 -9621
rect 5937 -9891 6017 -9881
rect 5937 -9951 5947 -9891
rect 6007 -9901 6017 -9891
rect 6257 -9891 6337 -9881
rect 6257 -9901 6267 -9891
rect 6007 -9951 6267 -9901
rect 6327 -9951 6337 -9891
rect 5937 -9961 6337 -9951
rect 6393 -9541 6793 -9531
rect 6393 -9601 6403 -9541
rect 6463 -9591 6723 -9541
rect 6463 -9601 6473 -9591
rect 6393 -9611 6473 -9601
rect 6713 -9601 6723 -9591
rect 6783 -9601 6793 -9541
rect 6713 -9611 6793 -9601
rect 6393 -9881 6453 -9611
rect 6723 -9621 6793 -9611
rect 6533 -9671 6563 -9651
rect 6513 -9711 6563 -9671
rect 6623 -9671 6653 -9651
rect 6623 -9711 6673 -9671
rect 6513 -9781 6673 -9711
rect 6513 -9821 6563 -9781
rect 6533 -9841 6563 -9821
rect 6623 -9821 6673 -9781
rect 6623 -9841 6653 -9821
rect 6733 -9881 6793 -9621
rect 6393 -9891 6473 -9881
rect 6393 -9951 6403 -9891
rect 6463 -9901 6473 -9891
rect 6713 -9891 6793 -9881
rect 6713 -9901 6723 -9891
rect 6463 -9951 6723 -9901
rect 6783 -9951 6793 -9891
rect 6393 -9961 6793 -9951
rect 6851 -9541 7251 -9531
rect 6851 -9601 6861 -9541
rect 6921 -9591 7181 -9541
rect 6921 -9601 6931 -9591
rect 6851 -9611 6931 -9601
rect 7171 -9601 7181 -9591
rect 7241 -9601 7251 -9541
rect 7171 -9611 7251 -9601
rect 6851 -9881 6911 -9611
rect 7181 -9621 7251 -9611
rect 6991 -9671 7021 -9651
rect 6971 -9711 7021 -9671
rect 7081 -9671 7111 -9651
rect 7081 -9711 7131 -9671
rect 6971 -9781 7131 -9711
rect 6971 -9821 7021 -9781
rect 6991 -9841 7021 -9821
rect 7081 -9821 7131 -9781
rect 7081 -9841 7111 -9821
rect 7191 -9881 7251 -9621
rect 6851 -9891 6931 -9881
rect 6851 -9951 6861 -9891
rect 6921 -9901 6931 -9891
rect 7171 -9891 7251 -9881
rect 7171 -9901 7181 -9891
rect 6921 -9951 7181 -9901
rect 7241 -9951 7251 -9891
rect 6851 -9961 7251 -9951
rect 7307 -9541 7707 -9531
rect 7307 -9601 7317 -9541
rect 7377 -9591 7637 -9541
rect 7377 -9601 7387 -9591
rect 7307 -9611 7387 -9601
rect 7627 -9601 7637 -9591
rect 7697 -9601 7707 -9541
rect 7627 -9611 7707 -9601
rect 7307 -9881 7367 -9611
rect 7637 -9621 7707 -9611
rect 7447 -9671 7477 -9651
rect 7427 -9711 7477 -9671
rect 7537 -9671 7567 -9651
rect 7537 -9711 7587 -9671
rect 7427 -9781 7587 -9711
rect 7427 -9821 7477 -9781
rect 7447 -9841 7477 -9821
rect 7537 -9821 7587 -9781
rect 7537 -9841 7567 -9821
rect 7647 -9881 7707 -9621
rect 7307 -9891 7387 -9881
rect 7307 -9951 7317 -9891
rect 7377 -9901 7387 -9891
rect 7627 -9891 7707 -9881
rect 7627 -9901 7637 -9891
rect 7377 -9951 7637 -9901
rect 7697 -9951 7707 -9891
rect 7307 -9961 7707 -9951
rect 7763 -9541 8163 -9531
rect 7763 -9601 7773 -9541
rect 7833 -9591 8093 -9541
rect 7833 -9601 7843 -9591
rect 7763 -9611 7843 -9601
rect 8083 -9601 8093 -9591
rect 8153 -9601 8163 -9541
rect 8083 -9611 8163 -9601
rect 7763 -9881 7823 -9611
rect 8093 -9621 8163 -9611
rect 7903 -9671 7933 -9651
rect 7883 -9711 7933 -9671
rect 7993 -9671 8023 -9651
rect 7993 -9711 8043 -9671
rect 7883 -9781 8043 -9711
rect 7883 -9821 7933 -9781
rect 7903 -9841 7933 -9821
rect 7993 -9821 8043 -9781
rect 7993 -9841 8023 -9821
rect 8103 -9881 8163 -9621
rect 7763 -9891 7843 -9881
rect 7763 -9951 7773 -9891
rect 7833 -9901 7843 -9891
rect 8083 -9891 8163 -9881
rect 8083 -9901 8093 -9891
rect 7833 -9951 8093 -9901
rect 8153 -9951 8163 -9891
rect 7763 -9961 8163 -9951
rect 8237 -9541 8637 -9531
rect 8237 -9601 8247 -9541
rect 8307 -9591 8567 -9541
rect 8307 -9601 8317 -9591
rect 8237 -9611 8317 -9601
rect 8557 -9601 8567 -9591
rect 8627 -9601 8637 -9541
rect 8557 -9611 8637 -9601
rect 8237 -9881 8297 -9611
rect 8567 -9621 8637 -9611
rect 8377 -9671 8407 -9651
rect 8357 -9711 8407 -9671
rect 8467 -9671 8497 -9651
rect 8467 -9711 8517 -9671
rect 8357 -9781 8517 -9711
rect 8357 -9821 8407 -9781
rect 8377 -9841 8407 -9821
rect 8467 -9821 8517 -9781
rect 8467 -9841 8497 -9821
rect 8577 -9881 8637 -9621
rect 8237 -9891 8317 -9881
rect 8237 -9951 8247 -9891
rect 8307 -9901 8317 -9891
rect 8557 -9891 8637 -9881
rect 8557 -9901 8567 -9891
rect 8307 -9951 8567 -9901
rect 8627 -9951 8637 -9891
rect 8237 -9961 8637 -9951
rect 8693 -9541 9093 -9531
rect 8693 -9601 8703 -9541
rect 8763 -9591 9023 -9541
rect 8763 -9601 8773 -9591
rect 8693 -9611 8773 -9601
rect 9013 -9601 9023 -9591
rect 9083 -9601 9093 -9541
rect 9013 -9611 9093 -9601
rect 8693 -9881 8753 -9611
rect 9023 -9621 9093 -9611
rect 8833 -9671 8863 -9651
rect 8813 -9711 8863 -9671
rect 8923 -9671 8953 -9651
rect 8923 -9711 8973 -9671
rect 8813 -9781 8973 -9711
rect 8813 -9821 8863 -9781
rect 8833 -9841 8863 -9821
rect 8923 -9821 8973 -9781
rect 8923 -9841 8953 -9821
rect 9033 -9881 9093 -9621
rect 8693 -9891 8773 -9881
rect 8693 -9951 8703 -9891
rect 8763 -9901 8773 -9891
rect 9013 -9891 9093 -9881
rect 9013 -9901 9023 -9891
rect 8763 -9951 9023 -9901
rect 9083 -9951 9093 -9891
rect 8693 -9961 9093 -9951
rect 9151 -9541 9551 -9531
rect 9151 -9601 9161 -9541
rect 9221 -9591 9481 -9541
rect 9221 -9601 9231 -9591
rect 9151 -9611 9231 -9601
rect 9471 -9601 9481 -9591
rect 9541 -9601 9551 -9541
rect 9471 -9611 9551 -9601
rect 9151 -9881 9211 -9611
rect 9481 -9621 9551 -9611
rect 9291 -9671 9321 -9651
rect 9271 -9711 9321 -9671
rect 9381 -9671 9411 -9651
rect 9381 -9711 9431 -9671
rect 9271 -9781 9431 -9711
rect 9271 -9821 9321 -9781
rect 9291 -9841 9321 -9821
rect 9381 -9821 9431 -9781
rect 9381 -9841 9411 -9821
rect 9491 -9881 9551 -9621
rect 9151 -9891 9231 -9881
rect 9151 -9951 9161 -9891
rect 9221 -9901 9231 -9891
rect 9471 -9891 9551 -9881
rect 9471 -9901 9481 -9891
rect 9221 -9951 9481 -9901
rect 9541 -9951 9551 -9891
rect 9151 -9961 9551 -9951
rect 9607 -9541 10007 -9531
rect 9607 -9601 9617 -9541
rect 9677 -9591 9937 -9541
rect 9677 -9601 9687 -9591
rect 9607 -9611 9687 -9601
rect 9927 -9601 9937 -9591
rect 9997 -9601 10007 -9541
rect 9927 -9611 10007 -9601
rect 9607 -9881 9667 -9611
rect 9937 -9621 10007 -9611
rect 9747 -9671 9777 -9651
rect 9727 -9711 9777 -9671
rect 9837 -9671 9867 -9651
rect 9837 -9711 9887 -9671
rect 9727 -9781 9887 -9711
rect 9727 -9821 9777 -9781
rect 9747 -9841 9777 -9821
rect 9837 -9821 9887 -9781
rect 9837 -9841 9867 -9821
rect 9947 -9881 10007 -9621
rect 9607 -9891 9687 -9881
rect 9607 -9951 9617 -9891
rect 9677 -9901 9687 -9891
rect 9927 -9891 10007 -9881
rect 9927 -9901 9937 -9891
rect 9677 -9951 9937 -9901
rect 9997 -9951 10007 -9891
rect 9607 -9961 10007 -9951
rect 10063 -9541 10463 -9531
rect 10063 -9601 10073 -9541
rect 10133 -9591 10393 -9541
rect 10133 -9601 10143 -9591
rect 10063 -9611 10143 -9601
rect 10383 -9601 10393 -9591
rect 10453 -9601 10463 -9541
rect 10383 -9611 10463 -9601
rect 10063 -9881 10123 -9611
rect 10393 -9621 10463 -9611
rect 10203 -9671 10233 -9651
rect 10183 -9711 10233 -9671
rect 10293 -9671 10323 -9651
rect 10293 -9711 10343 -9671
rect 10183 -9781 10343 -9711
rect 10183 -9821 10233 -9781
rect 10203 -9841 10233 -9821
rect 10293 -9821 10343 -9781
rect 10293 -9841 10323 -9821
rect 10403 -9881 10463 -9621
rect 10063 -9891 10143 -9881
rect 10063 -9951 10073 -9891
rect 10133 -9901 10143 -9891
rect 10383 -9891 10463 -9881
rect 10383 -9901 10393 -9891
rect 10133 -9951 10393 -9901
rect 10453 -9951 10463 -9891
rect 10063 -9961 10463 -9951
rect 10521 -9541 10921 -9531
rect 10521 -9601 10531 -9541
rect 10591 -9591 10851 -9541
rect 10591 -9601 10601 -9591
rect 10521 -9611 10601 -9601
rect 10841 -9601 10851 -9591
rect 10911 -9601 10921 -9541
rect 10841 -9611 10921 -9601
rect 10521 -9881 10581 -9611
rect 10851 -9621 10921 -9611
rect 10661 -9671 10691 -9651
rect 10641 -9711 10691 -9671
rect 10751 -9671 10781 -9651
rect 10751 -9711 10801 -9671
rect 10641 -9781 10801 -9711
rect 10641 -9821 10691 -9781
rect 10661 -9841 10691 -9821
rect 10751 -9821 10801 -9781
rect 10751 -9841 10781 -9821
rect 10861 -9881 10921 -9621
rect 10521 -9891 10601 -9881
rect 10521 -9951 10531 -9891
rect 10591 -9901 10601 -9891
rect 10841 -9891 10921 -9881
rect 10841 -9901 10851 -9891
rect 10591 -9951 10851 -9901
rect 10911 -9951 10921 -9891
rect 10521 -9961 10921 -9951
rect 10977 -9541 11377 -9531
rect 10977 -9601 10987 -9541
rect 11047 -9591 11307 -9541
rect 11047 -9601 11057 -9591
rect 10977 -9611 11057 -9601
rect 11297 -9601 11307 -9591
rect 11367 -9601 11377 -9541
rect 11297 -9611 11377 -9601
rect 10977 -9881 11037 -9611
rect 11307 -9621 11377 -9611
rect 11117 -9671 11147 -9651
rect 11097 -9711 11147 -9671
rect 11207 -9671 11237 -9651
rect 11207 -9711 11257 -9671
rect 11097 -9781 11257 -9711
rect 11097 -9821 11147 -9781
rect 11117 -9841 11147 -9821
rect 11207 -9821 11257 -9781
rect 11207 -9841 11237 -9821
rect 11317 -9881 11377 -9621
rect 10977 -9891 11057 -9881
rect 10977 -9951 10987 -9891
rect 11047 -9901 11057 -9891
rect 11297 -9891 11377 -9881
rect 11297 -9901 11307 -9891
rect 11047 -9951 11307 -9901
rect 11367 -9951 11377 -9891
rect 10977 -9961 11377 -9951
rect 11433 -9541 11833 -9531
rect 11433 -9601 11443 -9541
rect 11503 -9591 11763 -9541
rect 11503 -9601 11513 -9591
rect 11433 -9611 11513 -9601
rect 11753 -9601 11763 -9591
rect 11823 -9601 11833 -9541
rect 11753 -9611 11833 -9601
rect 11433 -9881 11493 -9611
rect 11763 -9621 11833 -9611
rect 11573 -9671 11603 -9651
rect 11553 -9711 11603 -9671
rect 11663 -9671 11693 -9651
rect 11663 -9711 11713 -9671
rect 11553 -9781 11713 -9711
rect 11553 -9821 11603 -9781
rect 11573 -9841 11603 -9821
rect 11663 -9821 11713 -9781
rect 11663 -9841 11693 -9821
rect 11773 -9881 11833 -9621
rect 11433 -9891 11513 -9881
rect 11433 -9951 11443 -9891
rect 11503 -9901 11513 -9891
rect 11753 -9891 11833 -9881
rect 11753 -9901 11763 -9891
rect 11503 -9951 11763 -9901
rect 11823 -9951 11833 -9891
rect 11433 -9961 11833 -9951
rect 11891 -9541 12291 -9531
rect 11891 -9601 11901 -9541
rect 11961 -9591 12221 -9541
rect 11961 -9601 11971 -9591
rect 11891 -9611 11971 -9601
rect 12211 -9601 12221 -9591
rect 12281 -9601 12291 -9541
rect 12211 -9611 12291 -9601
rect 11891 -9881 11951 -9611
rect 12221 -9621 12291 -9611
rect 12031 -9671 12061 -9651
rect 12011 -9711 12061 -9671
rect 12121 -9671 12151 -9651
rect 12121 -9711 12171 -9671
rect 12011 -9781 12171 -9711
rect 12011 -9821 12061 -9781
rect 12031 -9841 12061 -9821
rect 12121 -9821 12171 -9781
rect 12121 -9841 12151 -9821
rect 12231 -9881 12291 -9621
rect 11891 -9891 11971 -9881
rect 11891 -9951 11901 -9891
rect 11961 -9901 11971 -9891
rect 12211 -9891 12291 -9881
rect 12211 -9901 12221 -9891
rect 11961 -9951 12221 -9901
rect 12281 -9951 12291 -9891
rect 11891 -9961 12291 -9951
rect 12347 -9541 12747 -9531
rect 12347 -9601 12357 -9541
rect 12417 -9591 12677 -9541
rect 12417 -9601 12427 -9591
rect 12347 -9611 12427 -9601
rect 12667 -9601 12677 -9591
rect 12737 -9601 12747 -9541
rect 12667 -9611 12747 -9601
rect 12347 -9881 12407 -9611
rect 12677 -9621 12747 -9611
rect 12487 -9671 12517 -9651
rect 12467 -9711 12517 -9671
rect 12577 -9671 12607 -9651
rect 12577 -9711 12627 -9671
rect 12467 -9781 12627 -9711
rect 12467 -9821 12517 -9781
rect 12487 -9841 12517 -9821
rect 12577 -9821 12627 -9781
rect 12577 -9841 12607 -9821
rect 12687 -9881 12747 -9621
rect 12347 -9891 12427 -9881
rect 12347 -9951 12357 -9891
rect 12417 -9901 12427 -9891
rect 12667 -9891 12747 -9881
rect 12667 -9901 12677 -9891
rect 12417 -9951 12677 -9901
rect 12737 -9951 12747 -9891
rect 12347 -9961 12747 -9951
rect 12803 -9541 13203 -9531
rect 12803 -9601 12813 -9541
rect 12873 -9591 13133 -9541
rect 12873 -9601 12883 -9591
rect 12803 -9611 12883 -9601
rect 13123 -9601 13133 -9591
rect 13193 -9601 13203 -9541
rect 13123 -9611 13203 -9601
rect 12803 -9881 12863 -9611
rect 13133 -9621 13203 -9611
rect 12943 -9671 12973 -9651
rect 12923 -9711 12973 -9671
rect 13033 -9671 13063 -9651
rect 13033 -9711 13083 -9671
rect 12923 -9781 13083 -9711
rect 12923 -9821 12973 -9781
rect 12943 -9841 12973 -9821
rect 13033 -9821 13083 -9781
rect 13033 -9841 13063 -9821
rect 13143 -9881 13203 -9621
rect 12803 -9891 12883 -9881
rect 12803 -9951 12813 -9891
rect 12873 -9901 12883 -9891
rect 13123 -9891 13203 -9881
rect 13123 -9901 13133 -9891
rect 12873 -9951 13133 -9901
rect 13193 -9951 13203 -9891
rect 12803 -9961 13203 -9951
rect 13261 -9541 13661 -9531
rect 13261 -9601 13271 -9541
rect 13331 -9591 13591 -9541
rect 13331 -9601 13341 -9591
rect 13261 -9611 13341 -9601
rect 13581 -9601 13591 -9591
rect 13651 -9601 13661 -9541
rect 13581 -9611 13661 -9601
rect 13261 -9881 13321 -9611
rect 13591 -9621 13661 -9611
rect 13401 -9671 13431 -9651
rect 13381 -9711 13431 -9671
rect 13491 -9671 13521 -9651
rect 13491 -9711 13541 -9671
rect 13381 -9781 13541 -9711
rect 13381 -9821 13431 -9781
rect 13401 -9841 13431 -9821
rect 13491 -9821 13541 -9781
rect 13491 -9841 13521 -9821
rect 13601 -9881 13661 -9621
rect 13261 -9891 13341 -9881
rect 13261 -9951 13271 -9891
rect 13331 -9901 13341 -9891
rect 13581 -9891 13661 -9881
rect 13581 -9901 13591 -9891
rect 13331 -9951 13591 -9901
rect 13651 -9951 13661 -9891
rect 13261 -9961 13661 -9951
rect 13717 -9541 14117 -9531
rect 13717 -9601 13727 -9541
rect 13787 -9591 14047 -9541
rect 13787 -9601 13797 -9591
rect 13717 -9611 13797 -9601
rect 14037 -9601 14047 -9591
rect 14107 -9601 14117 -9541
rect 14037 -9611 14117 -9601
rect 13717 -9881 13777 -9611
rect 14047 -9621 14117 -9611
rect 13857 -9671 13887 -9651
rect 13837 -9711 13887 -9671
rect 13947 -9671 13977 -9651
rect 13947 -9711 13997 -9671
rect 13837 -9781 13997 -9711
rect 13837 -9821 13887 -9781
rect 13857 -9841 13887 -9821
rect 13947 -9821 13997 -9781
rect 13947 -9841 13977 -9821
rect 14057 -9881 14117 -9621
rect 13717 -9891 13797 -9881
rect 13717 -9951 13727 -9891
rect 13787 -9901 13797 -9891
rect 14037 -9891 14117 -9881
rect 14037 -9901 14047 -9891
rect 13787 -9951 14047 -9901
rect 14107 -9951 14117 -9891
rect 13717 -9961 14117 -9951
rect 14173 -9541 14573 -9531
rect 14173 -9601 14183 -9541
rect 14243 -9591 14503 -9541
rect 14243 -9601 14253 -9591
rect 14173 -9611 14253 -9601
rect 14493 -9601 14503 -9591
rect 14563 -9601 14573 -9541
rect 14493 -9611 14573 -9601
rect 14173 -9881 14233 -9611
rect 14503 -9621 14573 -9611
rect 14313 -9671 14343 -9651
rect 14293 -9711 14343 -9671
rect 14403 -9671 14433 -9651
rect 14403 -9711 14453 -9671
rect 14293 -9781 14453 -9711
rect 14293 -9821 14343 -9781
rect 14313 -9841 14343 -9821
rect 14403 -9821 14453 -9781
rect 14403 -9841 14433 -9821
rect 14513 -9881 14573 -9621
rect 14173 -9891 14253 -9881
rect 14173 -9951 14183 -9891
rect 14243 -9901 14253 -9891
rect 14493 -9891 14573 -9881
rect 14493 -9901 14503 -9891
rect 14243 -9951 14503 -9901
rect 14563 -9951 14573 -9891
rect 14173 -9961 14573 -9951
rect 14631 -9541 15031 -9531
rect 14631 -9601 14641 -9541
rect 14701 -9591 14961 -9541
rect 14701 -9601 14711 -9591
rect 14631 -9611 14711 -9601
rect 14951 -9601 14961 -9591
rect 15021 -9601 15031 -9541
rect 14951 -9611 15031 -9601
rect 14631 -9881 14691 -9611
rect 14961 -9621 15031 -9611
rect 14771 -9671 14801 -9651
rect 14751 -9711 14801 -9671
rect 14861 -9671 14891 -9651
rect 14861 -9711 14911 -9671
rect 14751 -9781 14911 -9711
rect 14751 -9821 14801 -9781
rect 14771 -9841 14801 -9821
rect 14861 -9821 14911 -9781
rect 14861 -9841 14891 -9821
rect 14971 -9881 15031 -9621
rect 14631 -9891 14711 -9881
rect 14631 -9951 14641 -9891
rect 14701 -9901 14711 -9891
rect 14951 -9891 15031 -9881
rect 14951 -9901 14961 -9891
rect 14701 -9951 14961 -9901
rect 15021 -9951 15031 -9891
rect 14631 -9961 15031 -9951
rect 15087 -9541 15487 -9531
rect 15087 -9601 15097 -9541
rect 15157 -9591 15417 -9541
rect 15157 -9601 15167 -9591
rect 15087 -9611 15167 -9601
rect 15407 -9601 15417 -9591
rect 15477 -9601 15487 -9541
rect 15407 -9611 15487 -9601
rect 15087 -9881 15147 -9611
rect 15417 -9621 15487 -9611
rect 15227 -9671 15257 -9651
rect 15207 -9711 15257 -9671
rect 15317 -9671 15347 -9651
rect 15317 -9711 15367 -9671
rect 15207 -9781 15367 -9711
rect 15207 -9821 15257 -9781
rect 15227 -9841 15257 -9821
rect 15317 -9821 15367 -9781
rect 15317 -9841 15347 -9821
rect 15427 -9881 15487 -9621
rect 15087 -9891 15167 -9881
rect 15087 -9951 15097 -9891
rect 15157 -9901 15167 -9891
rect 15407 -9891 15487 -9881
rect 15407 -9901 15417 -9891
rect 15157 -9951 15417 -9901
rect 15477 -9951 15487 -9891
rect 15087 -9961 15487 -9951
rect 1 -10057 401 -10047
rect 1 -10117 11 -10057
rect 71 -10107 331 -10057
rect 71 -10117 81 -10107
rect 1 -10127 81 -10117
rect 321 -10117 331 -10107
rect 391 -10117 401 -10057
rect 321 -10127 401 -10117
rect 1 -10397 61 -10127
rect 331 -10137 401 -10127
rect 141 -10187 171 -10167
rect 121 -10227 171 -10187
rect 231 -10187 261 -10167
rect 231 -10227 281 -10187
rect 121 -10297 281 -10227
rect 121 -10337 171 -10297
rect 141 -10357 171 -10337
rect 231 -10337 281 -10297
rect 231 -10357 261 -10337
rect 341 -10397 401 -10137
rect 1 -10407 81 -10397
rect 1 -10467 11 -10407
rect 71 -10417 81 -10407
rect 321 -10407 401 -10397
rect 321 -10417 331 -10407
rect 71 -10467 331 -10417
rect 391 -10467 401 -10407
rect 1 -10477 401 -10467
rect 457 -10057 857 -10047
rect 457 -10117 467 -10057
rect 527 -10107 787 -10057
rect 527 -10117 537 -10107
rect 457 -10127 537 -10117
rect 777 -10117 787 -10107
rect 847 -10117 857 -10057
rect 777 -10127 857 -10117
rect 457 -10397 517 -10127
rect 787 -10137 857 -10127
rect 597 -10187 627 -10167
rect 577 -10227 627 -10187
rect 687 -10187 717 -10167
rect 687 -10227 737 -10187
rect 577 -10297 737 -10227
rect 577 -10337 627 -10297
rect 597 -10357 627 -10337
rect 687 -10337 737 -10297
rect 687 -10357 717 -10337
rect 797 -10397 857 -10137
rect 457 -10407 537 -10397
rect 457 -10467 467 -10407
rect 527 -10417 537 -10407
rect 777 -10407 857 -10397
rect 777 -10417 787 -10407
rect 527 -10467 787 -10417
rect 847 -10467 857 -10407
rect 457 -10477 857 -10467
rect 913 -10057 1313 -10047
rect 913 -10117 923 -10057
rect 983 -10107 1243 -10057
rect 983 -10117 993 -10107
rect 913 -10127 993 -10117
rect 1233 -10117 1243 -10107
rect 1303 -10117 1313 -10057
rect 1233 -10127 1313 -10117
rect 913 -10397 973 -10127
rect 1243 -10137 1313 -10127
rect 1053 -10187 1083 -10167
rect 1033 -10227 1083 -10187
rect 1143 -10187 1173 -10167
rect 1143 -10227 1193 -10187
rect 1033 -10297 1193 -10227
rect 1033 -10337 1083 -10297
rect 1053 -10357 1083 -10337
rect 1143 -10337 1193 -10297
rect 1143 -10357 1173 -10337
rect 1253 -10397 1313 -10137
rect 913 -10407 993 -10397
rect 913 -10467 923 -10407
rect 983 -10417 993 -10407
rect 1233 -10407 1313 -10397
rect 1233 -10417 1243 -10407
rect 983 -10467 1243 -10417
rect 1303 -10467 1313 -10407
rect 913 -10477 1313 -10467
rect 1371 -10057 1771 -10047
rect 1371 -10117 1381 -10057
rect 1441 -10107 1701 -10057
rect 1441 -10117 1451 -10107
rect 1371 -10127 1451 -10117
rect 1691 -10117 1701 -10107
rect 1761 -10117 1771 -10057
rect 1691 -10127 1771 -10117
rect 1371 -10397 1431 -10127
rect 1701 -10137 1771 -10127
rect 1511 -10187 1541 -10167
rect 1491 -10227 1541 -10187
rect 1601 -10187 1631 -10167
rect 1601 -10227 1651 -10187
rect 1491 -10297 1651 -10227
rect 1491 -10337 1541 -10297
rect 1511 -10357 1541 -10337
rect 1601 -10337 1651 -10297
rect 1601 -10357 1631 -10337
rect 1711 -10397 1771 -10137
rect 1371 -10407 1451 -10397
rect 1371 -10467 1381 -10407
rect 1441 -10417 1451 -10407
rect 1691 -10407 1771 -10397
rect 1691 -10417 1701 -10407
rect 1441 -10467 1701 -10417
rect 1761 -10467 1771 -10407
rect 1371 -10477 1771 -10467
rect 1827 -10057 2227 -10047
rect 1827 -10117 1837 -10057
rect 1897 -10107 2157 -10057
rect 1897 -10117 1907 -10107
rect 1827 -10127 1907 -10117
rect 2147 -10117 2157 -10107
rect 2217 -10117 2227 -10057
rect 2147 -10127 2227 -10117
rect 1827 -10397 1887 -10127
rect 2157 -10137 2227 -10127
rect 1967 -10187 1997 -10167
rect 1947 -10227 1997 -10187
rect 2057 -10187 2087 -10167
rect 2057 -10227 2107 -10187
rect 1947 -10297 2107 -10227
rect 1947 -10337 1997 -10297
rect 1967 -10357 1997 -10337
rect 2057 -10337 2107 -10297
rect 2057 -10357 2087 -10337
rect 2167 -10397 2227 -10137
rect 1827 -10407 1907 -10397
rect 1827 -10467 1837 -10407
rect 1897 -10417 1907 -10407
rect 2147 -10407 2227 -10397
rect 2147 -10417 2157 -10407
rect 1897 -10467 2157 -10417
rect 2217 -10467 2227 -10407
rect 1827 -10477 2227 -10467
rect 2283 -10057 2683 -10047
rect 2283 -10117 2293 -10057
rect 2353 -10107 2613 -10057
rect 2353 -10117 2363 -10107
rect 2283 -10127 2363 -10117
rect 2603 -10117 2613 -10107
rect 2673 -10117 2683 -10057
rect 2603 -10127 2683 -10117
rect 2283 -10397 2343 -10127
rect 2613 -10137 2683 -10127
rect 2423 -10187 2453 -10167
rect 2403 -10227 2453 -10187
rect 2513 -10187 2543 -10167
rect 2513 -10227 2563 -10187
rect 2403 -10297 2563 -10227
rect 2403 -10337 2453 -10297
rect 2423 -10357 2453 -10337
rect 2513 -10337 2563 -10297
rect 2513 -10357 2543 -10337
rect 2623 -10397 2683 -10137
rect 2283 -10407 2363 -10397
rect 2283 -10467 2293 -10407
rect 2353 -10417 2363 -10407
rect 2603 -10407 2683 -10397
rect 2603 -10417 2613 -10407
rect 2353 -10467 2613 -10417
rect 2673 -10467 2683 -10407
rect 2283 -10477 2683 -10467
rect 2741 -10057 3141 -10047
rect 2741 -10117 2751 -10057
rect 2811 -10107 3071 -10057
rect 2811 -10117 2821 -10107
rect 2741 -10127 2821 -10117
rect 3061 -10117 3071 -10107
rect 3131 -10117 3141 -10057
rect 3061 -10127 3141 -10117
rect 2741 -10397 2801 -10127
rect 3071 -10137 3141 -10127
rect 2881 -10187 2911 -10167
rect 2861 -10227 2911 -10187
rect 2971 -10187 3001 -10167
rect 2971 -10227 3021 -10187
rect 2861 -10297 3021 -10227
rect 2861 -10337 2911 -10297
rect 2881 -10357 2911 -10337
rect 2971 -10337 3021 -10297
rect 2971 -10357 3001 -10337
rect 3081 -10397 3141 -10137
rect 2741 -10407 2821 -10397
rect 2741 -10467 2751 -10407
rect 2811 -10417 2821 -10407
rect 3061 -10407 3141 -10397
rect 3061 -10417 3071 -10407
rect 2811 -10467 3071 -10417
rect 3131 -10467 3141 -10407
rect 2741 -10477 3141 -10467
rect 3197 -10057 3597 -10047
rect 3197 -10117 3207 -10057
rect 3267 -10107 3527 -10057
rect 3267 -10117 3277 -10107
rect 3197 -10127 3277 -10117
rect 3517 -10117 3527 -10107
rect 3587 -10117 3597 -10057
rect 3517 -10127 3597 -10117
rect 3197 -10397 3257 -10127
rect 3527 -10137 3597 -10127
rect 3337 -10187 3367 -10167
rect 3317 -10227 3367 -10187
rect 3427 -10187 3457 -10167
rect 3427 -10227 3477 -10187
rect 3317 -10297 3477 -10227
rect 3317 -10337 3367 -10297
rect 3337 -10357 3367 -10337
rect 3427 -10337 3477 -10297
rect 3427 -10357 3457 -10337
rect 3537 -10397 3597 -10137
rect 3197 -10407 3277 -10397
rect 3197 -10467 3207 -10407
rect 3267 -10417 3277 -10407
rect 3517 -10407 3597 -10397
rect 3517 -10417 3527 -10407
rect 3267 -10467 3527 -10417
rect 3587 -10467 3597 -10407
rect 3197 -10477 3597 -10467
rect 3653 -10057 4053 -10047
rect 3653 -10117 3663 -10057
rect 3723 -10107 3983 -10057
rect 3723 -10117 3733 -10107
rect 3653 -10127 3733 -10117
rect 3973 -10117 3983 -10107
rect 4043 -10117 4053 -10057
rect 3973 -10127 4053 -10117
rect 3653 -10397 3713 -10127
rect 3983 -10137 4053 -10127
rect 3793 -10187 3823 -10167
rect 3773 -10227 3823 -10187
rect 3883 -10187 3913 -10167
rect 3883 -10227 3933 -10187
rect 3773 -10297 3933 -10227
rect 3773 -10337 3823 -10297
rect 3793 -10357 3823 -10337
rect 3883 -10337 3933 -10297
rect 3883 -10357 3913 -10337
rect 3993 -10397 4053 -10137
rect 3653 -10407 3733 -10397
rect 3653 -10467 3663 -10407
rect 3723 -10417 3733 -10407
rect 3973 -10407 4053 -10397
rect 3973 -10417 3983 -10407
rect 3723 -10467 3983 -10417
rect 4043 -10467 4053 -10407
rect 3653 -10477 4053 -10467
rect 4111 -10057 4511 -10047
rect 4111 -10117 4121 -10057
rect 4181 -10107 4441 -10057
rect 4181 -10117 4191 -10107
rect 4111 -10127 4191 -10117
rect 4431 -10117 4441 -10107
rect 4501 -10117 4511 -10057
rect 4431 -10127 4511 -10117
rect 4111 -10397 4171 -10127
rect 4441 -10137 4511 -10127
rect 4251 -10187 4281 -10167
rect 4231 -10227 4281 -10187
rect 4341 -10187 4371 -10167
rect 4341 -10227 4391 -10187
rect 4231 -10297 4391 -10227
rect 4231 -10337 4281 -10297
rect 4251 -10357 4281 -10337
rect 4341 -10337 4391 -10297
rect 4341 -10357 4371 -10337
rect 4451 -10397 4511 -10137
rect 4111 -10407 4191 -10397
rect 4111 -10467 4121 -10407
rect 4181 -10417 4191 -10407
rect 4431 -10407 4511 -10397
rect 4431 -10417 4441 -10407
rect 4181 -10467 4441 -10417
rect 4501 -10467 4511 -10407
rect 4111 -10477 4511 -10467
rect 4567 -10057 4967 -10047
rect 4567 -10117 4577 -10057
rect 4637 -10107 4897 -10057
rect 4637 -10117 4647 -10107
rect 4567 -10127 4647 -10117
rect 4887 -10117 4897 -10107
rect 4957 -10117 4967 -10057
rect 4887 -10127 4967 -10117
rect 4567 -10397 4627 -10127
rect 4897 -10137 4967 -10127
rect 4707 -10187 4737 -10167
rect 4687 -10227 4737 -10187
rect 4797 -10187 4827 -10167
rect 4797 -10227 4847 -10187
rect 4687 -10297 4847 -10227
rect 4687 -10337 4737 -10297
rect 4707 -10357 4737 -10337
rect 4797 -10337 4847 -10297
rect 4797 -10357 4827 -10337
rect 4907 -10397 4967 -10137
rect 4567 -10407 4647 -10397
rect 4567 -10467 4577 -10407
rect 4637 -10417 4647 -10407
rect 4887 -10407 4967 -10397
rect 4887 -10417 4897 -10407
rect 4637 -10467 4897 -10417
rect 4957 -10467 4967 -10407
rect 4567 -10477 4967 -10467
rect 5023 -10057 5423 -10047
rect 5023 -10117 5033 -10057
rect 5093 -10107 5353 -10057
rect 5093 -10117 5103 -10107
rect 5023 -10127 5103 -10117
rect 5343 -10117 5353 -10107
rect 5413 -10117 5423 -10057
rect 5343 -10127 5423 -10117
rect 5023 -10397 5083 -10127
rect 5353 -10137 5423 -10127
rect 5163 -10187 5193 -10167
rect 5143 -10227 5193 -10187
rect 5253 -10187 5283 -10167
rect 5253 -10227 5303 -10187
rect 5143 -10297 5303 -10227
rect 5143 -10337 5193 -10297
rect 5163 -10357 5193 -10337
rect 5253 -10337 5303 -10297
rect 5253 -10357 5283 -10337
rect 5363 -10397 5423 -10137
rect 5023 -10407 5103 -10397
rect 5023 -10467 5033 -10407
rect 5093 -10417 5103 -10407
rect 5343 -10407 5423 -10397
rect 5343 -10417 5353 -10407
rect 5093 -10467 5353 -10417
rect 5413 -10467 5423 -10407
rect 5023 -10477 5423 -10467
rect 5481 -10057 5881 -10047
rect 5481 -10117 5491 -10057
rect 5551 -10107 5811 -10057
rect 5551 -10117 5561 -10107
rect 5481 -10127 5561 -10117
rect 5801 -10117 5811 -10107
rect 5871 -10117 5881 -10057
rect 5801 -10127 5881 -10117
rect 5481 -10397 5541 -10127
rect 5811 -10137 5881 -10127
rect 5621 -10187 5651 -10167
rect 5601 -10227 5651 -10187
rect 5711 -10187 5741 -10167
rect 5711 -10227 5761 -10187
rect 5601 -10297 5761 -10227
rect 5601 -10337 5651 -10297
rect 5621 -10357 5651 -10337
rect 5711 -10337 5761 -10297
rect 5711 -10357 5741 -10337
rect 5821 -10397 5881 -10137
rect 5481 -10407 5561 -10397
rect 5481 -10467 5491 -10407
rect 5551 -10417 5561 -10407
rect 5801 -10407 5881 -10397
rect 5801 -10417 5811 -10407
rect 5551 -10467 5811 -10417
rect 5871 -10467 5881 -10407
rect 5481 -10477 5881 -10467
rect 5937 -10057 6337 -10047
rect 5937 -10117 5947 -10057
rect 6007 -10107 6267 -10057
rect 6007 -10117 6017 -10107
rect 5937 -10127 6017 -10117
rect 6257 -10117 6267 -10107
rect 6327 -10117 6337 -10057
rect 6257 -10127 6337 -10117
rect 5937 -10397 5997 -10127
rect 6267 -10137 6337 -10127
rect 6077 -10187 6107 -10167
rect 6057 -10227 6107 -10187
rect 6167 -10187 6197 -10167
rect 6167 -10227 6217 -10187
rect 6057 -10297 6217 -10227
rect 6057 -10337 6107 -10297
rect 6077 -10357 6107 -10337
rect 6167 -10337 6217 -10297
rect 6167 -10357 6197 -10337
rect 6277 -10397 6337 -10137
rect 5937 -10407 6017 -10397
rect 5937 -10467 5947 -10407
rect 6007 -10417 6017 -10407
rect 6257 -10407 6337 -10397
rect 6257 -10417 6267 -10407
rect 6007 -10467 6267 -10417
rect 6327 -10467 6337 -10407
rect 5937 -10477 6337 -10467
rect 6393 -10057 6793 -10047
rect 6393 -10117 6403 -10057
rect 6463 -10107 6723 -10057
rect 6463 -10117 6473 -10107
rect 6393 -10127 6473 -10117
rect 6713 -10117 6723 -10107
rect 6783 -10117 6793 -10057
rect 6713 -10127 6793 -10117
rect 6393 -10397 6453 -10127
rect 6723 -10137 6793 -10127
rect 6533 -10187 6563 -10167
rect 6513 -10227 6563 -10187
rect 6623 -10187 6653 -10167
rect 6623 -10227 6673 -10187
rect 6513 -10297 6673 -10227
rect 6513 -10337 6563 -10297
rect 6533 -10357 6563 -10337
rect 6623 -10337 6673 -10297
rect 6623 -10357 6653 -10337
rect 6733 -10397 6793 -10137
rect 6393 -10407 6473 -10397
rect 6393 -10467 6403 -10407
rect 6463 -10417 6473 -10407
rect 6713 -10407 6793 -10397
rect 6713 -10417 6723 -10407
rect 6463 -10467 6723 -10417
rect 6783 -10467 6793 -10407
rect 6393 -10477 6793 -10467
rect 6851 -10057 7251 -10047
rect 6851 -10117 6861 -10057
rect 6921 -10107 7181 -10057
rect 6921 -10117 6931 -10107
rect 6851 -10127 6931 -10117
rect 7171 -10117 7181 -10107
rect 7241 -10117 7251 -10057
rect 7171 -10127 7251 -10117
rect 6851 -10397 6911 -10127
rect 7181 -10137 7251 -10127
rect 6991 -10187 7021 -10167
rect 6971 -10227 7021 -10187
rect 7081 -10187 7111 -10167
rect 7081 -10227 7131 -10187
rect 6971 -10297 7131 -10227
rect 6971 -10337 7021 -10297
rect 6991 -10357 7021 -10337
rect 7081 -10337 7131 -10297
rect 7081 -10357 7111 -10337
rect 7191 -10397 7251 -10137
rect 6851 -10407 6931 -10397
rect 6851 -10467 6861 -10407
rect 6921 -10417 6931 -10407
rect 7171 -10407 7251 -10397
rect 7171 -10417 7181 -10407
rect 6921 -10467 7181 -10417
rect 7241 -10467 7251 -10407
rect 6851 -10477 7251 -10467
rect 7307 -10057 7707 -10047
rect 7307 -10117 7317 -10057
rect 7377 -10107 7637 -10057
rect 7377 -10117 7387 -10107
rect 7307 -10127 7387 -10117
rect 7627 -10117 7637 -10107
rect 7697 -10117 7707 -10057
rect 7627 -10127 7707 -10117
rect 7307 -10397 7367 -10127
rect 7637 -10137 7707 -10127
rect 7447 -10187 7477 -10167
rect 7427 -10227 7477 -10187
rect 7537 -10187 7567 -10167
rect 7537 -10227 7587 -10187
rect 7427 -10297 7587 -10227
rect 7427 -10337 7477 -10297
rect 7447 -10357 7477 -10337
rect 7537 -10337 7587 -10297
rect 7537 -10357 7567 -10337
rect 7647 -10397 7707 -10137
rect 7307 -10407 7387 -10397
rect 7307 -10467 7317 -10407
rect 7377 -10417 7387 -10407
rect 7627 -10407 7707 -10397
rect 7627 -10417 7637 -10407
rect 7377 -10467 7637 -10417
rect 7697 -10467 7707 -10407
rect 7307 -10477 7707 -10467
rect 7763 -10057 8163 -10047
rect 7763 -10117 7773 -10057
rect 7833 -10107 8093 -10057
rect 7833 -10117 7843 -10107
rect 7763 -10127 7843 -10117
rect 8083 -10117 8093 -10107
rect 8153 -10117 8163 -10057
rect 8083 -10127 8163 -10117
rect 7763 -10397 7823 -10127
rect 8093 -10137 8163 -10127
rect 7903 -10187 7933 -10167
rect 7883 -10227 7933 -10187
rect 7993 -10187 8023 -10167
rect 7993 -10227 8043 -10187
rect 7883 -10297 8043 -10227
rect 7883 -10337 7933 -10297
rect 7903 -10357 7933 -10337
rect 7993 -10337 8043 -10297
rect 7993 -10357 8023 -10337
rect 8103 -10397 8163 -10137
rect 7763 -10407 7843 -10397
rect 7763 -10467 7773 -10407
rect 7833 -10417 7843 -10407
rect 8083 -10407 8163 -10397
rect 8083 -10417 8093 -10407
rect 7833 -10467 8093 -10417
rect 8153 -10467 8163 -10407
rect 7763 -10477 8163 -10467
rect 8237 -10057 8637 -10047
rect 8237 -10117 8247 -10057
rect 8307 -10107 8567 -10057
rect 8307 -10117 8317 -10107
rect 8237 -10127 8317 -10117
rect 8557 -10117 8567 -10107
rect 8627 -10117 8637 -10057
rect 8557 -10127 8637 -10117
rect 8237 -10397 8297 -10127
rect 8567 -10137 8637 -10127
rect 8377 -10187 8407 -10167
rect 8357 -10227 8407 -10187
rect 8467 -10187 8497 -10167
rect 8467 -10227 8517 -10187
rect 8357 -10297 8517 -10227
rect 8357 -10337 8407 -10297
rect 8377 -10357 8407 -10337
rect 8467 -10337 8517 -10297
rect 8467 -10357 8497 -10337
rect 8577 -10397 8637 -10137
rect 8237 -10407 8317 -10397
rect 8237 -10467 8247 -10407
rect 8307 -10417 8317 -10407
rect 8557 -10407 8637 -10397
rect 8557 -10417 8567 -10407
rect 8307 -10467 8567 -10417
rect 8627 -10467 8637 -10407
rect 8237 -10477 8637 -10467
rect 8693 -10057 9093 -10047
rect 8693 -10117 8703 -10057
rect 8763 -10107 9023 -10057
rect 8763 -10117 8773 -10107
rect 8693 -10127 8773 -10117
rect 9013 -10117 9023 -10107
rect 9083 -10117 9093 -10057
rect 9013 -10127 9093 -10117
rect 8693 -10397 8753 -10127
rect 9023 -10137 9093 -10127
rect 8833 -10187 8863 -10167
rect 8813 -10227 8863 -10187
rect 8923 -10187 8953 -10167
rect 8923 -10227 8973 -10187
rect 8813 -10297 8973 -10227
rect 8813 -10337 8863 -10297
rect 8833 -10357 8863 -10337
rect 8923 -10337 8973 -10297
rect 8923 -10357 8953 -10337
rect 9033 -10397 9093 -10137
rect 8693 -10407 8773 -10397
rect 8693 -10467 8703 -10407
rect 8763 -10417 8773 -10407
rect 9013 -10407 9093 -10397
rect 9013 -10417 9023 -10407
rect 8763 -10467 9023 -10417
rect 9083 -10467 9093 -10407
rect 8693 -10477 9093 -10467
rect 9151 -10057 9551 -10047
rect 9151 -10117 9161 -10057
rect 9221 -10107 9481 -10057
rect 9221 -10117 9231 -10107
rect 9151 -10127 9231 -10117
rect 9471 -10117 9481 -10107
rect 9541 -10117 9551 -10057
rect 9471 -10127 9551 -10117
rect 9151 -10397 9211 -10127
rect 9481 -10137 9551 -10127
rect 9291 -10187 9321 -10167
rect 9271 -10227 9321 -10187
rect 9381 -10187 9411 -10167
rect 9381 -10227 9431 -10187
rect 9271 -10297 9431 -10227
rect 9271 -10337 9321 -10297
rect 9291 -10357 9321 -10337
rect 9381 -10337 9431 -10297
rect 9381 -10357 9411 -10337
rect 9491 -10397 9551 -10137
rect 9151 -10407 9231 -10397
rect 9151 -10467 9161 -10407
rect 9221 -10417 9231 -10407
rect 9471 -10407 9551 -10397
rect 9471 -10417 9481 -10407
rect 9221 -10467 9481 -10417
rect 9541 -10467 9551 -10407
rect 9151 -10477 9551 -10467
rect 9607 -10057 10007 -10047
rect 9607 -10117 9617 -10057
rect 9677 -10107 9937 -10057
rect 9677 -10117 9687 -10107
rect 9607 -10127 9687 -10117
rect 9927 -10117 9937 -10107
rect 9997 -10117 10007 -10057
rect 9927 -10127 10007 -10117
rect 9607 -10397 9667 -10127
rect 9937 -10137 10007 -10127
rect 9747 -10187 9777 -10167
rect 9727 -10227 9777 -10187
rect 9837 -10187 9867 -10167
rect 9837 -10227 9887 -10187
rect 9727 -10297 9887 -10227
rect 9727 -10337 9777 -10297
rect 9747 -10357 9777 -10337
rect 9837 -10337 9887 -10297
rect 9837 -10357 9867 -10337
rect 9947 -10397 10007 -10137
rect 9607 -10407 9687 -10397
rect 9607 -10467 9617 -10407
rect 9677 -10417 9687 -10407
rect 9927 -10407 10007 -10397
rect 9927 -10417 9937 -10407
rect 9677 -10467 9937 -10417
rect 9997 -10467 10007 -10407
rect 9607 -10477 10007 -10467
rect 10063 -10057 10463 -10047
rect 10063 -10117 10073 -10057
rect 10133 -10107 10393 -10057
rect 10133 -10117 10143 -10107
rect 10063 -10127 10143 -10117
rect 10383 -10117 10393 -10107
rect 10453 -10117 10463 -10057
rect 10383 -10127 10463 -10117
rect 10063 -10397 10123 -10127
rect 10393 -10137 10463 -10127
rect 10203 -10187 10233 -10167
rect 10183 -10227 10233 -10187
rect 10293 -10187 10323 -10167
rect 10293 -10227 10343 -10187
rect 10183 -10297 10343 -10227
rect 10183 -10337 10233 -10297
rect 10203 -10357 10233 -10337
rect 10293 -10337 10343 -10297
rect 10293 -10357 10323 -10337
rect 10403 -10397 10463 -10137
rect 10063 -10407 10143 -10397
rect 10063 -10467 10073 -10407
rect 10133 -10417 10143 -10407
rect 10383 -10407 10463 -10397
rect 10383 -10417 10393 -10407
rect 10133 -10467 10393 -10417
rect 10453 -10467 10463 -10407
rect 10063 -10477 10463 -10467
rect 10521 -10057 10921 -10047
rect 10521 -10117 10531 -10057
rect 10591 -10107 10851 -10057
rect 10591 -10117 10601 -10107
rect 10521 -10127 10601 -10117
rect 10841 -10117 10851 -10107
rect 10911 -10117 10921 -10057
rect 10841 -10127 10921 -10117
rect 10521 -10397 10581 -10127
rect 10851 -10137 10921 -10127
rect 10661 -10187 10691 -10167
rect 10641 -10227 10691 -10187
rect 10751 -10187 10781 -10167
rect 10751 -10227 10801 -10187
rect 10641 -10297 10801 -10227
rect 10641 -10337 10691 -10297
rect 10661 -10357 10691 -10337
rect 10751 -10337 10801 -10297
rect 10751 -10357 10781 -10337
rect 10861 -10397 10921 -10137
rect 10521 -10407 10601 -10397
rect 10521 -10467 10531 -10407
rect 10591 -10417 10601 -10407
rect 10841 -10407 10921 -10397
rect 10841 -10417 10851 -10407
rect 10591 -10467 10851 -10417
rect 10911 -10467 10921 -10407
rect 10521 -10477 10921 -10467
rect 10977 -10057 11377 -10047
rect 10977 -10117 10987 -10057
rect 11047 -10107 11307 -10057
rect 11047 -10117 11057 -10107
rect 10977 -10127 11057 -10117
rect 11297 -10117 11307 -10107
rect 11367 -10117 11377 -10057
rect 11297 -10127 11377 -10117
rect 10977 -10397 11037 -10127
rect 11307 -10137 11377 -10127
rect 11117 -10187 11147 -10167
rect 11097 -10227 11147 -10187
rect 11207 -10187 11237 -10167
rect 11207 -10227 11257 -10187
rect 11097 -10297 11257 -10227
rect 11097 -10337 11147 -10297
rect 11117 -10357 11147 -10337
rect 11207 -10337 11257 -10297
rect 11207 -10357 11237 -10337
rect 11317 -10397 11377 -10137
rect 10977 -10407 11057 -10397
rect 10977 -10467 10987 -10407
rect 11047 -10417 11057 -10407
rect 11297 -10407 11377 -10397
rect 11297 -10417 11307 -10407
rect 11047 -10467 11307 -10417
rect 11367 -10467 11377 -10407
rect 10977 -10477 11377 -10467
rect 11433 -10057 11833 -10047
rect 11433 -10117 11443 -10057
rect 11503 -10107 11763 -10057
rect 11503 -10117 11513 -10107
rect 11433 -10127 11513 -10117
rect 11753 -10117 11763 -10107
rect 11823 -10117 11833 -10057
rect 11753 -10127 11833 -10117
rect 11433 -10397 11493 -10127
rect 11763 -10137 11833 -10127
rect 11573 -10187 11603 -10167
rect 11553 -10227 11603 -10187
rect 11663 -10187 11693 -10167
rect 11663 -10227 11713 -10187
rect 11553 -10297 11713 -10227
rect 11553 -10337 11603 -10297
rect 11573 -10357 11603 -10337
rect 11663 -10337 11713 -10297
rect 11663 -10357 11693 -10337
rect 11773 -10397 11833 -10137
rect 11433 -10407 11513 -10397
rect 11433 -10467 11443 -10407
rect 11503 -10417 11513 -10407
rect 11753 -10407 11833 -10397
rect 11753 -10417 11763 -10407
rect 11503 -10467 11763 -10417
rect 11823 -10467 11833 -10407
rect 11433 -10477 11833 -10467
rect 11891 -10057 12291 -10047
rect 11891 -10117 11901 -10057
rect 11961 -10107 12221 -10057
rect 11961 -10117 11971 -10107
rect 11891 -10127 11971 -10117
rect 12211 -10117 12221 -10107
rect 12281 -10117 12291 -10057
rect 12211 -10127 12291 -10117
rect 11891 -10397 11951 -10127
rect 12221 -10137 12291 -10127
rect 12031 -10187 12061 -10167
rect 12011 -10227 12061 -10187
rect 12121 -10187 12151 -10167
rect 12121 -10227 12171 -10187
rect 12011 -10297 12171 -10227
rect 12011 -10337 12061 -10297
rect 12031 -10357 12061 -10337
rect 12121 -10337 12171 -10297
rect 12121 -10357 12151 -10337
rect 12231 -10397 12291 -10137
rect 11891 -10407 11971 -10397
rect 11891 -10467 11901 -10407
rect 11961 -10417 11971 -10407
rect 12211 -10407 12291 -10397
rect 12211 -10417 12221 -10407
rect 11961 -10467 12221 -10417
rect 12281 -10467 12291 -10407
rect 11891 -10477 12291 -10467
rect 12347 -10057 12747 -10047
rect 12347 -10117 12357 -10057
rect 12417 -10107 12677 -10057
rect 12417 -10117 12427 -10107
rect 12347 -10127 12427 -10117
rect 12667 -10117 12677 -10107
rect 12737 -10117 12747 -10057
rect 12667 -10127 12747 -10117
rect 12347 -10397 12407 -10127
rect 12677 -10137 12747 -10127
rect 12487 -10187 12517 -10167
rect 12467 -10227 12517 -10187
rect 12577 -10187 12607 -10167
rect 12577 -10227 12627 -10187
rect 12467 -10297 12627 -10227
rect 12467 -10337 12517 -10297
rect 12487 -10357 12517 -10337
rect 12577 -10337 12627 -10297
rect 12577 -10357 12607 -10337
rect 12687 -10397 12747 -10137
rect 12347 -10407 12427 -10397
rect 12347 -10467 12357 -10407
rect 12417 -10417 12427 -10407
rect 12667 -10407 12747 -10397
rect 12667 -10417 12677 -10407
rect 12417 -10467 12677 -10417
rect 12737 -10467 12747 -10407
rect 12347 -10477 12747 -10467
rect 12803 -10057 13203 -10047
rect 12803 -10117 12813 -10057
rect 12873 -10107 13133 -10057
rect 12873 -10117 12883 -10107
rect 12803 -10127 12883 -10117
rect 13123 -10117 13133 -10107
rect 13193 -10117 13203 -10057
rect 13123 -10127 13203 -10117
rect 12803 -10397 12863 -10127
rect 13133 -10137 13203 -10127
rect 12943 -10187 12973 -10167
rect 12923 -10227 12973 -10187
rect 13033 -10187 13063 -10167
rect 13033 -10227 13083 -10187
rect 12923 -10297 13083 -10227
rect 12923 -10337 12973 -10297
rect 12943 -10357 12973 -10337
rect 13033 -10337 13083 -10297
rect 13033 -10357 13063 -10337
rect 13143 -10397 13203 -10137
rect 12803 -10407 12883 -10397
rect 12803 -10467 12813 -10407
rect 12873 -10417 12883 -10407
rect 13123 -10407 13203 -10397
rect 13123 -10417 13133 -10407
rect 12873 -10467 13133 -10417
rect 13193 -10467 13203 -10407
rect 12803 -10477 13203 -10467
rect 13261 -10057 13661 -10047
rect 13261 -10117 13271 -10057
rect 13331 -10107 13591 -10057
rect 13331 -10117 13341 -10107
rect 13261 -10127 13341 -10117
rect 13581 -10117 13591 -10107
rect 13651 -10117 13661 -10057
rect 13581 -10127 13661 -10117
rect 13261 -10397 13321 -10127
rect 13591 -10137 13661 -10127
rect 13401 -10187 13431 -10167
rect 13381 -10227 13431 -10187
rect 13491 -10187 13521 -10167
rect 13491 -10227 13541 -10187
rect 13381 -10297 13541 -10227
rect 13381 -10337 13431 -10297
rect 13401 -10357 13431 -10337
rect 13491 -10337 13541 -10297
rect 13491 -10357 13521 -10337
rect 13601 -10397 13661 -10137
rect 13261 -10407 13341 -10397
rect 13261 -10467 13271 -10407
rect 13331 -10417 13341 -10407
rect 13581 -10407 13661 -10397
rect 13581 -10417 13591 -10407
rect 13331 -10467 13591 -10417
rect 13651 -10467 13661 -10407
rect 13261 -10477 13661 -10467
rect 13717 -10057 14117 -10047
rect 13717 -10117 13727 -10057
rect 13787 -10107 14047 -10057
rect 13787 -10117 13797 -10107
rect 13717 -10127 13797 -10117
rect 14037 -10117 14047 -10107
rect 14107 -10117 14117 -10057
rect 14037 -10127 14117 -10117
rect 13717 -10397 13777 -10127
rect 14047 -10137 14117 -10127
rect 13857 -10187 13887 -10167
rect 13837 -10227 13887 -10187
rect 13947 -10187 13977 -10167
rect 13947 -10227 13997 -10187
rect 13837 -10297 13997 -10227
rect 13837 -10337 13887 -10297
rect 13857 -10357 13887 -10337
rect 13947 -10337 13997 -10297
rect 13947 -10357 13977 -10337
rect 14057 -10397 14117 -10137
rect 13717 -10407 13797 -10397
rect 13717 -10467 13727 -10407
rect 13787 -10417 13797 -10407
rect 14037 -10407 14117 -10397
rect 14037 -10417 14047 -10407
rect 13787 -10467 14047 -10417
rect 14107 -10467 14117 -10407
rect 13717 -10477 14117 -10467
rect 14173 -10057 14573 -10047
rect 14173 -10117 14183 -10057
rect 14243 -10107 14503 -10057
rect 14243 -10117 14253 -10107
rect 14173 -10127 14253 -10117
rect 14493 -10117 14503 -10107
rect 14563 -10117 14573 -10057
rect 14493 -10127 14573 -10117
rect 14173 -10397 14233 -10127
rect 14503 -10137 14573 -10127
rect 14313 -10187 14343 -10167
rect 14293 -10227 14343 -10187
rect 14403 -10187 14433 -10167
rect 14403 -10227 14453 -10187
rect 14293 -10297 14453 -10227
rect 14293 -10337 14343 -10297
rect 14313 -10357 14343 -10337
rect 14403 -10337 14453 -10297
rect 14403 -10357 14433 -10337
rect 14513 -10397 14573 -10137
rect 14173 -10407 14253 -10397
rect 14173 -10467 14183 -10407
rect 14243 -10417 14253 -10407
rect 14493 -10407 14573 -10397
rect 14493 -10417 14503 -10407
rect 14243 -10467 14503 -10417
rect 14563 -10467 14573 -10407
rect 14173 -10477 14573 -10467
rect 14631 -10057 15031 -10047
rect 14631 -10117 14641 -10057
rect 14701 -10107 14961 -10057
rect 14701 -10117 14711 -10107
rect 14631 -10127 14711 -10117
rect 14951 -10117 14961 -10107
rect 15021 -10117 15031 -10057
rect 14951 -10127 15031 -10117
rect 14631 -10397 14691 -10127
rect 14961 -10137 15031 -10127
rect 14771 -10187 14801 -10167
rect 14751 -10227 14801 -10187
rect 14861 -10187 14891 -10167
rect 14861 -10227 14911 -10187
rect 14751 -10297 14911 -10227
rect 14751 -10337 14801 -10297
rect 14771 -10357 14801 -10337
rect 14861 -10337 14911 -10297
rect 14861 -10357 14891 -10337
rect 14971 -10397 15031 -10137
rect 14631 -10407 14711 -10397
rect 14631 -10467 14641 -10407
rect 14701 -10417 14711 -10407
rect 14951 -10407 15031 -10397
rect 14951 -10417 14961 -10407
rect 14701 -10467 14961 -10417
rect 15021 -10467 15031 -10407
rect 14631 -10477 15031 -10467
rect 15087 -10057 15487 -10047
rect 15087 -10117 15097 -10057
rect 15157 -10107 15417 -10057
rect 15157 -10117 15167 -10107
rect 15087 -10127 15167 -10117
rect 15407 -10117 15417 -10107
rect 15477 -10117 15487 -10057
rect 15407 -10127 15487 -10117
rect 15087 -10397 15147 -10127
rect 15417 -10137 15487 -10127
rect 15227 -10187 15257 -10167
rect 15207 -10227 15257 -10187
rect 15317 -10187 15347 -10167
rect 15317 -10227 15367 -10187
rect 15207 -10297 15367 -10227
rect 15207 -10337 15257 -10297
rect 15227 -10357 15257 -10337
rect 15317 -10337 15367 -10297
rect 15317 -10357 15347 -10337
rect 15427 -10397 15487 -10137
rect 15087 -10407 15167 -10397
rect 15087 -10467 15097 -10407
rect 15157 -10417 15167 -10407
rect 15407 -10407 15487 -10397
rect 15407 -10417 15417 -10407
rect 15157 -10467 15417 -10417
rect 15477 -10467 15487 -10407
rect 15087 -10477 15487 -10467
rect 1 -10559 401 -10549
rect 1 -10619 11 -10559
rect 71 -10609 331 -10559
rect 71 -10619 81 -10609
rect 1 -10629 81 -10619
rect 321 -10619 331 -10609
rect 391 -10619 401 -10559
rect 321 -10629 401 -10619
rect 1 -10899 61 -10629
rect 331 -10639 401 -10629
rect 141 -10689 171 -10669
rect 121 -10729 171 -10689
rect 231 -10689 261 -10669
rect 231 -10729 281 -10689
rect 121 -10799 281 -10729
rect 121 -10839 171 -10799
rect 141 -10859 171 -10839
rect 231 -10839 281 -10799
rect 231 -10859 261 -10839
rect 341 -10899 401 -10639
rect 1 -10909 81 -10899
rect 1 -10969 11 -10909
rect 71 -10919 81 -10909
rect 321 -10909 401 -10899
rect 321 -10919 331 -10909
rect 71 -10969 331 -10919
rect 391 -10969 401 -10909
rect 1 -10979 401 -10969
rect 457 -10559 857 -10549
rect 457 -10619 467 -10559
rect 527 -10609 787 -10559
rect 527 -10619 537 -10609
rect 457 -10629 537 -10619
rect 777 -10619 787 -10609
rect 847 -10619 857 -10559
rect 777 -10629 857 -10619
rect 457 -10899 517 -10629
rect 787 -10639 857 -10629
rect 597 -10689 627 -10669
rect 577 -10729 627 -10689
rect 687 -10689 717 -10669
rect 687 -10729 737 -10689
rect 577 -10799 737 -10729
rect 577 -10839 627 -10799
rect 597 -10859 627 -10839
rect 687 -10839 737 -10799
rect 687 -10859 717 -10839
rect 797 -10899 857 -10639
rect 457 -10909 537 -10899
rect 457 -10969 467 -10909
rect 527 -10919 537 -10909
rect 777 -10909 857 -10899
rect 777 -10919 787 -10909
rect 527 -10969 787 -10919
rect 847 -10969 857 -10909
rect 457 -10979 857 -10969
rect 913 -10559 1313 -10549
rect 913 -10619 923 -10559
rect 983 -10609 1243 -10559
rect 983 -10619 993 -10609
rect 913 -10629 993 -10619
rect 1233 -10619 1243 -10609
rect 1303 -10619 1313 -10559
rect 1233 -10629 1313 -10619
rect 913 -10899 973 -10629
rect 1243 -10639 1313 -10629
rect 1053 -10689 1083 -10669
rect 1033 -10729 1083 -10689
rect 1143 -10689 1173 -10669
rect 1143 -10729 1193 -10689
rect 1033 -10799 1193 -10729
rect 1033 -10839 1083 -10799
rect 1053 -10859 1083 -10839
rect 1143 -10839 1193 -10799
rect 1143 -10859 1173 -10839
rect 1253 -10899 1313 -10639
rect 913 -10909 993 -10899
rect 913 -10969 923 -10909
rect 983 -10919 993 -10909
rect 1233 -10909 1313 -10899
rect 1233 -10919 1243 -10909
rect 983 -10969 1243 -10919
rect 1303 -10969 1313 -10909
rect 913 -10979 1313 -10969
rect 1371 -10559 1771 -10549
rect 1371 -10619 1381 -10559
rect 1441 -10609 1701 -10559
rect 1441 -10619 1451 -10609
rect 1371 -10629 1451 -10619
rect 1691 -10619 1701 -10609
rect 1761 -10619 1771 -10559
rect 1691 -10629 1771 -10619
rect 1371 -10899 1431 -10629
rect 1701 -10639 1771 -10629
rect 1511 -10689 1541 -10669
rect 1491 -10729 1541 -10689
rect 1601 -10689 1631 -10669
rect 1601 -10729 1651 -10689
rect 1491 -10799 1651 -10729
rect 1491 -10839 1541 -10799
rect 1511 -10859 1541 -10839
rect 1601 -10839 1651 -10799
rect 1601 -10859 1631 -10839
rect 1711 -10899 1771 -10639
rect 1371 -10909 1451 -10899
rect 1371 -10969 1381 -10909
rect 1441 -10919 1451 -10909
rect 1691 -10909 1771 -10899
rect 1691 -10919 1701 -10909
rect 1441 -10969 1701 -10919
rect 1761 -10969 1771 -10909
rect 1371 -10979 1771 -10969
rect 1827 -10559 2227 -10549
rect 1827 -10619 1837 -10559
rect 1897 -10609 2157 -10559
rect 1897 -10619 1907 -10609
rect 1827 -10629 1907 -10619
rect 2147 -10619 2157 -10609
rect 2217 -10619 2227 -10559
rect 2147 -10629 2227 -10619
rect 1827 -10899 1887 -10629
rect 2157 -10639 2227 -10629
rect 1967 -10689 1997 -10669
rect 1947 -10729 1997 -10689
rect 2057 -10689 2087 -10669
rect 2057 -10729 2107 -10689
rect 1947 -10799 2107 -10729
rect 1947 -10839 1997 -10799
rect 1967 -10859 1997 -10839
rect 2057 -10839 2107 -10799
rect 2057 -10859 2087 -10839
rect 2167 -10899 2227 -10639
rect 1827 -10909 1907 -10899
rect 1827 -10969 1837 -10909
rect 1897 -10919 1907 -10909
rect 2147 -10909 2227 -10899
rect 2147 -10919 2157 -10909
rect 1897 -10969 2157 -10919
rect 2217 -10969 2227 -10909
rect 1827 -10979 2227 -10969
rect 2283 -10559 2683 -10549
rect 2283 -10619 2293 -10559
rect 2353 -10609 2613 -10559
rect 2353 -10619 2363 -10609
rect 2283 -10629 2363 -10619
rect 2603 -10619 2613 -10609
rect 2673 -10619 2683 -10559
rect 2603 -10629 2683 -10619
rect 2283 -10899 2343 -10629
rect 2613 -10639 2683 -10629
rect 2423 -10689 2453 -10669
rect 2403 -10729 2453 -10689
rect 2513 -10689 2543 -10669
rect 2513 -10729 2563 -10689
rect 2403 -10799 2563 -10729
rect 2403 -10839 2453 -10799
rect 2423 -10859 2453 -10839
rect 2513 -10839 2563 -10799
rect 2513 -10859 2543 -10839
rect 2623 -10899 2683 -10639
rect 2283 -10909 2363 -10899
rect 2283 -10969 2293 -10909
rect 2353 -10919 2363 -10909
rect 2603 -10909 2683 -10899
rect 2603 -10919 2613 -10909
rect 2353 -10969 2613 -10919
rect 2673 -10969 2683 -10909
rect 2283 -10979 2683 -10969
rect 2741 -10559 3141 -10549
rect 2741 -10619 2751 -10559
rect 2811 -10609 3071 -10559
rect 2811 -10619 2821 -10609
rect 2741 -10629 2821 -10619
rect 3061 -10619 3071 -10609
rect 3131 -10619 3141 -10559
rect 3061 -10629 3141 -10619
rect 2741 -10899 2801 -10629
rect 3071 -10639 3141 -10629
rect 2881 -10689 2911 -10669
rect 2861 -10729 2911 -10689
rect 2971 -10689 3001 -10669
rect 2971 -10729 3021 -10689
rect 2861 -10799 3021 -10729
rect 2861 -10839 2911 -10799
rect 2881 -10859 2911 -10839
rect 2971 -10839 3021 -10799
rect 2971 -10859 3001 -10839
rect 3081 -10899 3141 -10639
rect 2741 -10909 2821 -10899
rect 2741 -10969 2751 -10909
rect 2811 -10919 2821 -10909
rect 3061 -10909 3141 -10899
rect 3061 -10919 3071 -10909
rect 2811 -10969 3071 -10919
rect 3131 -10969 3141 -10909
rect 2741 -10979 3141 -10969
rect 3197 -10559 3597 -10549
rect 3197 -10619 3207 -10559
rect 3267 -10609 3527 -10559
rect 3267 -10619 3277 -10609
rect 3197 -10629 3277 -10619
rect 3517 -10619 3527 -10609
rect 3587 -10619 3597 -10559
rect 3517 -10629 3597 -10619
rect 3197 -10899 3257 -10629
rect 3527 -10639 3597 -10629
rect 3337 -10689 3367 -10669
rect 3317 -10729 3367 -10689
rect 3427 -10689 3457 -10669
rect 3427 -10729 3477 -10689
rect 3317 -10799 3477 -10729
rect 3317 -10839 3367 -10799
rect 3337 -10859 3367 -10839
rect 3427 -10839 3477 -10799
rect 3427 -10859 3457 -10839
rect 3537 -10899 3597 -10639
rect 3197 -10909 3277 -10899
rect 3197 -10969 3207 -10909
rect 3267 -10919 3277 -10909
rect 3517 -10909 3597 -10899
rect 3517 -10919 3527 -10909
rect 3267 -10969 3527 -10919
rect 3587 -10969 3597 -10909
rect 3197 -10979 3597 -10969
rect 3653 -10559 4053 -10549
rect 3653 -10619 3663 -10559
rect 3723 -10609 3983 -10559
rect 3723 -10619 3733 -10609
rect 3653 -10629 3733 -10619
rect 3973 -10619 3983 -10609
rect 4043 -10619 4053 -10559
rect 3973 -10629 4053 -10619
rect 3653 -10899 3713 -10629
rect 3983 -10639 4053 -10629
rect 3793 -10689 3823 -10669
rect 3773 -10729 3823 -10689
rect 3883 -10689 3913 -10669
rect 3883 -10729 3933 -10689
rect 3773 -10799 3933 -10729
rect 3773 -10839 3823 -10799
rect 3793 -10859 3823 -10839
rect 3883 -10839 3933 -10799
rect 3883 -10859 3913 -10839
rect 3993 -10899 4053 -10639
rect 3653 -10909 3733 -10899
rect 3653 -10969 3663 -10909
rect 3723 -10919 3733 -10909
rect 3973 -10909 4053 -10899
rect 3973 -10919 3983 -10909
rect 3723 -10969 3983 -10919
rect 4043 -10969 4053 -10909
rect 3653 -10979 4053 -10969
rect 4111 -10559 4511 -10549
rect 4111 -10619 4121 -10559
rect 4181 -10609 4441 -10559
rect 4181 -10619 4191 -10609
rect 4111 -10629 4191 -10619
rect 4431 -10619 4441 -10609
rect 4501 -10619 4511 -10559
rect 4431 -10629 4511 -10619
rect 4111 -10899 4171 -10629
rect 4441 -10639 4511 -10629
rect 4251 -10689 4281 -10669
rect 4231 -10729 4281 -10689
rect 4341 -10689 4371 -10669
rect 4341 -10729 4391 -10689
rect 4231 -10799 4391 -10729
rect 4231 -10839 4281 -10799
rect 4251 -10859 4281 -10839
rect 4341 -10839 4391 -10799
rect 4341 -10859 4371 -10839
rect 4451 -10899 4511 -10639
rect 4111 -10909 4191 -10899
rect 4111 -10969 4121 -10909
rect 4181 -10919 4191 -10909
rect 4431 -10909 4511 -10899
rect 4431 -10919 4441 -10909
rect 4181 -10969 4441 -10919
rect 4501 -10969 4511 -10909
rect 4111 -10979 4511 -10969
rect 4567 -10559 4967 -10549
rect 4567 -10619 4577 -10559
rect 4637 -10609 4897 -10559
rect 4637 -10619 4647 -10609
rect 4567 -10629 4647 -10619
rect 4887 -10619 4897 -10609
rect 4957 -10619 4967 -10559
rect 4887 -10629 4967 -10619
rect 4567 -10899 4627 -10629
rect 4897 -10639 4967 -10629
rect 4707 -10689 4737 -10669
rect 4687 -10729 4737 -10689
rect 4797 -10689 4827 -10669
rect 4797 -10729 4847 -10689
rect 4687 -10799 4847 -10729
rect 4687 -10839 4737 -10799
rect 4707 -10859 4737 -10839
rect 4797 -10839 4847 -10799
rect 4797 -10859 4827 -10839
rect 4907 -10899 4967 -10639
rect 4567 -10909 4647 -10899
rect 4567 -10969 4577 -10909
rect 4637 -10919 4647 -10909
rect 4887 -10909 4967 -10899
rect 4887 -10919 4897 -10909
rect 4637 -10969 4897 -10919
rect 4957 -10969 4967 -10909
rect 4567 -10979 4967 -10969
rect 5023 -10559 5423 -10549
rect 5023 -10619 5033 -10559
rect 5093 -10609 5353 -10559
rect 5093 -10619 5103 -10609
rect 5023 -10629 5103 -10619
rect 5343 -10619 5353 -10609
rect 5413 -10619 5423 -10559
rect 5343 -10629 5423 -10619
rect 5023 -10899 5083 -10629
rect 5353 -10639 5423 -10629
rect 5163 -10689 5193 -10669
rect 5143 -10729 5193 -10689
rect 5253 -10689 5283 -10669
rect 5253 -10729 5303 -10689
rect 5143 -10799 5303 -10729
rect 5143 -10839 5193 -10799
rect 5163 -10859 5193 -10839
rect 5253 -10839 5303 -10799
rect 5253 -10859 5283 -10839
rect 5363 -10899 5423 -10639
rect 5023 -10909 5103 -10899
rect 5023 -10969 5033 -10909
rect 5093 -10919 5103 -10909
rect 5343 -10909 5423 -10899
rect 5343 -10919 5353 -10909
rect 5093 -10969 5353 -10919
rect 5413 -10969 5423 -10909
rect 5023 -10979 5423 -10969
rect 5481 -10559 5881 -10549
rect 5481 -10619 5491 -10559
rect 5551 -10609 5811 -10559
rect 5551 -10619 5561 -10609
rect 5481 -10629 5561 -10619
rect 5801 -10619 5811 -10609
rect 5871 -10619 5881 -10559
rect 5801 -10629 5881 -10619
rect 5481 -10899 5541 -10629
rect 5811 -10639 5881 -10629
rect 5621 -10689 5651 -10669
rect 5601 -10729 5651 -10689
rect 5711 -10689 5741 -10669
rect 5711 -10729 5761 -10689
rect 5601 -10799 5761 -10729
rect 5601 -10839 5651 -10799
rect 5621 -10859 5651 -10839
rect 5711 -10839 5761 -10799
rect 5711 -10859 5741 -10839
rect 5821 -10899 5881 -10639
rect 5481 -10909 5561 -10899
rect 5481 -10969 5491 -10909
rect 5551 -10919 5561 -10909
rect 5801 -10909 5881 -10899
rect 5801 -10919 5811 -10909
rect 5551 -10969 5811 -10919
rect 5871 -10969 5881 -10909
rect 5481 -10979 5881 -10969
rect 5937 -10559 6337 -10549
rect 5937 -10619 5947 -10559
rect 6007 -10609 6267 -10559
rect 6007 -10619 6017 -10609
rect 5937 -10629 6017 -10619
rect 6257 -10619 6267 -10609
rect 6327 -10619 6337 -10559
rect 6257 -10629 6337 -10619
rect 5937 -10899 5997 -10629
rect 6267 -10639 6337 -10629
rect 6077 -10689 6107 -10669
rect 6057 -10729 6107 -10689
rect 6167 -10689 6197 -10669
rect 6167 -10729 6217 -10689
rect 6057 -10799 6217 -10729
rect 6057 -10839 6107 -10799
rect 6077 -10859 6107 -10839
rect 6167 -10839 6217 -10799
rect 6167 -10859 6197 -10839
rect 6277 -10899 6337 -10639
rect 5937 -10909 6017 -10899
rect 5937 -10969 5947 -10909
rect 6007 -10919 6017 -10909
rect 6257 -10909 6337 -10899
rect 6257 -10919 6267 -10909
rect 6007 -10969 6267 -10919
rect 6327 -10969 6337 -10909
rect 5937 -10979 6337 -10969
rect 6393 -10559 6793 -10549
rect 6393 -10619 6403 -10559
rect 6463 -10609 6723 -10559
rect 6463 -10619 6473 -10609
rect 6393 -10629 6473 -10619
rect 6713 -10619 6723 -10609
rect 6783 -10619 6793 -10559
rect 6713 -10629 6793 -10619
rect 6393 -10899 6453 -10629
rect 6723 -10639 6793 -10629
rect 6533 -10689 6563 -10669
rect 6513 -10729 6563 -10689
rect 6623 -10689 6653 -10669
rect 6623 -10729 6673 -10689
rect 6513 -10799 6673 -10729
rect 6513 -10839 6563 -10799
rect 6533 -10859 6563 -10839
rect 6623 -10839 6673 -10799
rect 6623 -10859 6653 -10839
rect 6733 -10899 6793 -10639
rect 6393 -10909 6473 -10899
rect 6393 -10969 6403 -10909
rect 6463 -10919 6473 -10909
rect 6713 -10909 6793 -10899
rect 6713 -10919 6723 -10909
rect 6463 -10969 6723 -10919
rect 6783 -10969 6793 -10909
rect 6393 -10979 6793 -10969
rect 6851 -10559 7251 -10549
rect 6851 -10619 6861 -10559
rect 6921 -10609 7181 -10559
rect 6921 -10619 6931 -10609
rect 6851 -10629 6931 -10619
rect 7171 -10619 7181 -10609
rect 7241 -10619 7251 -10559
rect 7171 -10629 7251 -10619
rect 6851 -10899 6911 -10629
rect 7181 -10639 7251 -10629
rect 6991 -10689 7021 -10669
rect 6971 -10729 7021 -10689
rect 7081 -10689 7111 -10669
rect 7081 -10729 7131 -10689
rect 6971 -10799 7131 -10729
rect 6971 -10839 7021 -10799
rect 6991 -10859 7021 -10839
rect 7081 -10839 7131 -10799
rect 7081 -10859 7111 -10839
rect 7191 -10899 7251 -10639
rect 6851 -10909 6931 -10899
rect 6851 -10969 6861 -10909
rect 6921 -10919 6931 -10909
rect 7171 -10909 7251 -10899
rect 7171 -10919 7181 -10909
rect 6921 -10969 7181 -10919
rect 7241 -10969 7251 -10909
rect 6851 -10979 7251 -10969
rect 7307 -10559 7707 -10549
rect 7307 -10619 7317 -10559
rect 7377 -10609 7637 -10559
rect 7377 -10619 7387 -10609
rect 7307 -10629 7387 -10619
rect 7627 -10619 7637 -10609
rect 7697 -10619 7707 -10559
rect 7627 -10629 7707 -10619
rect 7307 -10899 7367 -10629
rect 7637 -10639 7707 -10629
rect 7447 -10689 7477 -10669
rect 7427 -10729 7477 -10689
rect 7537 -10689 7567 -10669
rect 7537 -10729 7587 -10689
rect 7427 -10799 7587 -10729
rect 7427 -10839 7477 -10799
rect 7447 -10859 7477 -10839
rect 7537 -10839 7587 -10799
rect 7537 -10859 7567 -10839
rect 7647 -10899 7707 -10639
rect 7307 -10909 7387 -10899
rect 7307 -10969 7317 -10909
rect 7377 -10919 7387 -10909
rect 7627 -10909 7707 -10899
rect 7627 -10919 7637 -10909
rect 7377 -10969 7637 -10919
rect 7697 -10969 7707 -10909
rect 7307 -10979 7707 -10969
rect 7763 -10559 8163 -10549
rect 7763 -10619 7773 -10559
rect 7833 -10609 8093 -10559
rect 7833 -10619 7843 -10609
rect 7763 -10629 7843 -10619
rect 8083 -10619 8093 -10609
rect 8153 -10619 8163 -10559
rect 8083 -10629 8163 -10619
rect 7763 -10899 7823 -10629
rect 8093 -10639 8163 -10629
rect 7903 -10689 7933 -10669
rect 7883 -10729 7933 -10689
rect 7993 -10689 8023 -10669
rect 7993 -10729 8043 -10689
rect 7883 -10799 8043 -10729
rect 7883 -10839 7933 -10799
rect 7903 -10859 7933 -10839
rect 7993 -10839 8043 -10799
rect 7993 -10859 8023 -10839
rect 8103 -10899 8163 -10639
rect 7763 -10909 7843 -10899
rect 7763 -10969 7773 -10909
rect 7833 -10919 7843 -10909
rect 8083 -10909 8163 -10899
rect 8083 -10919 8093 -10909
rect 7833 -10969 8093 -10919
rect 8153 -10969 8163 -10909
rect 7763 -10979 8163 -10969
rect 8237 -10559 8637 -10549
rect 8237 -10619 8247 -10559
rect 8307 -10609 8567 -10559
rect 8307 -10619 8317 -10609
rect 8237 -10629 8317 -10619
rect 8557 -10619 8567 -10609
rect 8627 -10619 8637 -10559
rect 8557 -10629 8637 -10619
rect 8237 -10899 8297 -10629
rect 8567 -10639 8637 -10629
rect 8377 -10689 8407 -10669
rect 8357 -10729 8407 -10689
rect 8467 -10689 8497 -10669
rect 8467 -10729 8517 -10689
rect 8357 -10799 8517 -10729
rect 8357 -10839 8407 -10799
rect 8377 -10859 8407 -10839
rect 8467 -10839 8517 -10799
rect 8467 -10859 8497 -10839
rect 8577 -10899 8637 -10639
rect 8237 -10909 8317 -10899
rect 8237 -10969 8247 -10909
rect 8307 -10919 8317 -10909
rect 8557 -10909 8637 -10899
rect 8557 -10919 8567 -10909
rect 8307 -10969 8567 -10919
rect 8627 -10969 8637 -10909
rect 8237 -10979 8637 -10969
rect 8693 -10559 9093 -10549
rect 8693 -10619 8703 -10559
rect 8763 -10609 9023 -10559
rect 8763 -10619 8773 -10609
rect 8693 -10629 8773 -10619
rect 9013 -10619 9023 -10609
rect 9083 -10619 9093 -10559
rect 9013 -10629 9093 -10619
rect 8693 -10899 8753 -10629
rect 9023 -10639 9093 -10629
rect 8833 -10689 8863 -10669
rect 8813 -10729 8863 -10689
rect 8923 -10689 8953 -10669
rect 8923 -10729 8973 -10689
rect 8813 -10799 8973 -10729
rect 8813 -10839 8863 -10799
rect 8833 -10859 8863 -10839
rect 8923 -10839 8973 -10799
rect 8923 -10859 8953 -10839
rect 9033 -10899 9093 -10639
rect 8693 -10909 8773 -10899
rect 8693 -10969 8703 -10909
rect 8763 -10919 8773 -10909
rect 9013 -10909 9093 -10899
rect 9013 -10919 9023 -10909
rect 8763 -10969 9023 -10919
rect 9083 -10969 9093 -10909
rect 8693 -10979 9093 -10969
rect 9151 -10559 9551 -10549
rect 9151 -10619 9161 -10559
rect 9221 -10609 9481 -10559
rect 9221 -10619 9231 -10609
rect 9151 -10629 9231 -10619
rect 9471 -10619 9481 -10609
rect 9541 -10619 9551 -10559
rect 9471 -10629 9551 -10619
rect 9151 -10899 9211 -10629
rect 9481 -10639 9551 -10629
rect 9291 -10689 9321 -10669
rect 9271 -10729 9321 -10689
rect 9381 -10689 9411 -10669
rect 9381 -10729 9431 -10689
rect 9271 -10799 9431 -10729
rect 9271 -10839 9321 -10799
rect 9291 -10859 9321 -10839
rect 9381 -10839 9431 -10799
rect 9381 -10859 9411 -10839
rect 9491 -10899 9551 -10639
rect 9151 -10909 9231 -10899
rect 9151 -10969 9161 -10909
rect 9221 -10919 9231 -10909
rect 9471 -10909 9551 -10899
rect 9471 -10919 9481 -10909
rect 9221 -10969 9481 -10919
rect 9541 -10969 9551 -10909
rect 9151 -10979 9551 -10969
rect 9607 -10559 10007 -10549
rect 9607 -10619 9617 -10559
rect 9677 -10609 9937 -10559
rect 9677 -10619 9687 -10609
rect 9607 -10629 9687 -10619
rect 9927 -10619 9937 -10609
rect 9997 -10619 10007 -10559
rect 9927 -10629 10007 -10619
rect 9607 -10899 9667 -10629
rect 9937 -10639 10007 -10629
rect 9747 -10689 9777 -10669
rect 9727 -10729 9777 -10689
rect 9837 -10689 9867 -10669
rect 9837 -10729 9887 -10689
rect 9727 -10799 9887 -10729
rect 9727 -10839 9777 -10799
rect 9747 -10859 9777 -10839
rect 9837 -10839 9887 -10799
rect 9837 -10859 9867 -10839
rect 9947 -10899 10007 -10639
rect 9607 -10909 9687 -10899
rect 9607 -10969 9617 -10909
rect 9677 -10919 9687 -10909
rect 9927 -10909 10007 -10899
rect 9927 -10919 9937 -10909
rect 9677 -10969 9937 -10919
rect 9997 -10969 10007 -10909
rect 9607 -10979 10007 -10969
rect 10063 -10559 10463 -10549
rect 10063 -10619 10073 -10559
rect 10133 -10609 10393 -10559
rect 10133 -10619 10143 -10609
rect 10063 -10629 10143 -10619
rect 10383 -10619 10393 -10609
rect 10453 -10619 10463 -10559
rect 10383 -10629 10463 -10619
rect 10063 -10899 10123 -10629
rect 10393 -10639 10463 -10629
rect 10203 -10689 10233 -10669
rect 10183 -10729 10233 -10689
rect 10293 -10689 10323 -10669
rect 10293 -10729 10343 -10689
rect 10183 -10799 10343 -10729
rect 10183 -10839 10233 -10799
rect 10203 -10859 10233 -10839
rect 10293 -10839 10343 -10799
rect 10293 -10859 10323 -10839
rect 10403 -10899 10463 -10639
rect 10063 -10909 10143 -10899
rect 10063 -10969 10073 -10909
rect 10133 -10919 10143 -10909
rect 10383 -10909 10463 -10899
rect 10383 -10919 10393 -10909
rect 10133 -10969 10393 -10919
rect 10453 -10969 10463 -10909
rect 10063 -10979 10463 -10969
rect 10521 -10559 10921 -10549
rect 10521 -10619 10531 -10559
rect 10591 -10609 10851 -10559
rect 10591 -10619 10601 -10609
rect 10521 -10629 10601 -10619
rect 10841 -10619 10851 -10609
rect 10911 -10619 10921 -10559
rect 10841 -10629 10921 -10619
rect 10521 -10899 10581 -10629
rect 10851 -10639 10921 -10629
rect 10661 -10689 10691 -10669
rect 10641 -10729 10691 -10689
rect 10751 -10689 10781 -10669
rect 10751 -10729 10801 -10689
rect 10641 -10799 10801 -10729
rect 10641 -10839 10691 -10799
rect 10661 -10859 10691 -10839
rect 10751 -10839 10801 -10799
rect 10751 -10859 10781 -10839
rect 10861 -10899 10921 -10639
rect 10521 -10909 10601 -10899
rect 10521 -10969 10531 -10909
rect 10591 -10919 10601 -10909
rect 10841 -10909 10921 -10899
rect 10841 -10919 10851 -10909
rect 10591 -10969 10851 -10919
rect 10911 -10969 10921 -10909
rect 10521 -10979 10921 -10969
rect 10977 -10559 11377 -10549
rect 10977 -10619 10987 -10559
rect 11047 -10609 11307 -10559
rect 11047 -10619 11057 -10609
rect 10977 -10629 11057 -10619
rect 11297 -10619 11307 -10609
rect 11367 -10619 11377 -10559
rect 11297 -10629 11377 -10619
rect 10977 -10899 11037 -10629
rect 11307 -10639 11377 -10629
rect 11117 -10689 11147 -10669
rect 11097 -10729 11147 -10689
rect 11207 -10689 11237 -10669
rect 11207 -10729 11257 -10689
rect 11097 -10799 11257 -10729
rect 11097 -10839 11147 -10799
rect 11117 -10859 11147 -10839
rect 11207 -10839 11257 -10799
rect 11207 -10859 11237 -10839
rect 11317 -10899 11377 -10639
rect 10977 -10909 11057 -10899
rect 10977 -10969 10987 -10909
rect 11047 -10919 11057 -10909
rect 11297 -10909 11377 -10899
rect 11297 -10919 11307 -10909
rect 11047 -10969 11307 -10919
rect 11367 -10969 11377 -10909
rect 10977 -10979 11377 -10969
rect 11433 -10559 11833 -10549
rect 11433 -10619 11443 -10559
rect 11503 -10609 11763 -10559
rect 11503 -10619 11513 -10609
rect 11433 -10629 11513 -10619
rect 11753 -10619 11763 -10609
rect 11823 -10619 11833 -10559
rect 11753 -10629 11833 -10619
rect 11433 -10899 11493 -10629
rect 11763 -10639 11833 -10629
rect 11573 -10689 11603 -10669
rect 11553 -10729 11603 -10689
rect 11663 -10689 11693 -10669
rect 11663 -10729 11713 -10689
rect 11553 -10799 11713 -10729
rect 11553 -10839 11603 -10799
rect 11573 -10859 11603 -10839
rect 11663 -10839 11713 -10799
rect 11663 -10859 11693 -10839
rect 11773 -10899 11833 -10639
rect 11433 -10909 11513 -10899
rect 11433 -10969 11443 -10909
rect 11503 -10919 11513 -10909
rect 11753 -10909 11833 -10899
rect 11753 -10919 11763 -10909
rect 11503 -10969 11763 -10919
rect 11823 -10969 11833 -10909
rect 11433 -10979 11833 -10969
rect 11891 -10559 12291 -10549
rect 11891 -10619 11901 -10559
rect 11961 -10609 12221 -10559
rect 11961 -10619 11971 -10609
rect 11891 -10629 11971 -10619
rect 12211 -10619 12221 -10609
rect 12281 -10619 12291 -10559
rect 12211 -10629 12291 -10619
rect 11891 -10899 11951 -10629
rect 12221 -10639 12291 -10629
rect 12031 -10689 12061 -10669
rect 12011 -10729 12061 -10689
rect 12121 -10689 12151 -10669
rect 12121 -10729 12171 -10689
rect 12011 -10799 12171 -10729
rect 12011 -10839 12061 -10799
rect 12031 -10859 12061 -10839
rect 12121 -10839 12171 -10799
rect 12121 -10859 12151 -10839
rect 12231 -10899 12291 -10639
rect 11891 -10909 11971 -10899
rect 11891 -10969 11901 -10909
rect 11961 -10919 11971 -10909
rect 12211 -10909 12291 -10899
rect 12211 -10919 12221 -10909
rect 11961 -10969 12221 -10919
rect 12281 -10969 12291 -10909
rect 11891 -10979 12291 -10969
rect 12347 -10559 12747 -10549
rect 12347 -10619 12357 -10559
rect 12417 -10609 12677 -10559
rect 12417 -10619 12427 -10609
rect 12347 -10629 12427 -10619
rect 12667 -10619 12677 -10609
rect 12737 -10619 12747 -10559
rect 12667 -10629 12747 -10619
rect 12347 -10899 12407 -10629
rect 12677 -10639 12747 -10629
rect 12487 -10689 12517 -10669
rect 12467 -10729 12517 -10689
rect 12577 -10689 12607 -10669
rect 12577 -10729 12627 -10689
rect 12467 -10799 12627 -10729
rect 12467 -10839 12517 -10799
rect 12487 -10859 12517 -10839
rect 12577 -10839 12627 -10799
rect 12577 -10859 12607 -10839
rect 12687 -10899 12747 -10639
rect 12347 -10909 12427 -10899
rect 12347 -10969 12357 -10909
rect 12417 -10919 12427 -10909
rect 12667 -10909 12747 -10899
rect 12667 -10919 12677 -10909
rect 12417 -10969 12677 -10919
rect 12737 -10969 12747 -10909
rect 12347 -10979 12747 -10969
rect 12803 -10559 13203 -10549
rect 12803 -10619 12813 -10559
rect 12873 -10609 13133 -10559
rect 12873 -10619 12883 -10609
rect 12803 -10629 12883 -10619
rect 13123 -10619 13133 -10609
rect 13193 -10619 13203 -10559
rect 13123 -10629 13203 -10619
rect 12803 -10899 12863 -10629
rect 13133 -10639 13203 -10629
rect 12943 -10689 12973 -10669
rect 12923 -10729 12973 -10689
rect 13033 -10689 13063 -10669
rect 13033 -10729 13083 -10689
rect 12923 -10799 13083 -10729
rect 12923 -10839 12973 -10799
rect 12943 -10859 12973 -10839
rect 13033 -10839 13083 -10799
rect 13033 -10859 13063 -10839
rect 13143 -10899 13203 -10639
rect 12803 -10909 12883 -10899
rect 12803 -10969 12813 -10909
rect 12873 -10919 12883 -10909
rect 13123 -10909 13203 -10899
rect 13123 -10919 13133 -10909
rect 12873 -10969 13133 -10919
rect 13193 -10969 13203 -10909
rect 12803 -10979 13203 -10969
rect 13261 -10559 13661 -10549
rect 13261 -10619 13271 -10559
rect 13331 -10609 13591 -10559
rect 13331 -10619 13341 -10609
rect 13261 -10629 13341 -10619
rect 13581 -10619 13591 -10609
rect 13651 -10619 13661 -10559
rect 13581 -10629 13661 -10619
rect 13261 -10899 13321 -10629
rect 13591 -10639 13661 -10629
rect 13401 -10689 13431 -10669
rect 13381 -10729 13431 -10689
rect 13491 -10689 13521 -10669
rect 13491 -10729 13541 -10689
rect 13381 -10799 13541 -10729
rect 13381 -10839 13431 -10799
rect 13401 -10859 13431 -10839
rect 13491 -10839 13541 -10799
rect 13491 -10859 13521 -10839
rect 13601 -10899 13661 -10639
rect 13261 -10909 13341 -10899
rect 13261 -10969 13271 -10909
rect 13331 -10919 13341 -10909
rect 13581 -10909 13661 -10899
rect 13581 -10919 13591 -10909
rect 13331 -10969 13591 -10919
rect 13651 -10969 13661 -10909
rect 13261 -10979 13661 -10969
rect 13717 -10559 14117 -10549
rect 13717 -10619 13727 -10559
rect 13787 -10609 14047 -10559
rect 13787 -10619 13797 -10609
rect 13717 -10629 13797 -10619
rect 14037 -10619 14047 -10609
rect 14107 -10619 14117 -10559
rect 14037 -10629 14117 -10619
rect 13717 -10899 13777 -10629
rect 14047 -10639 14117 -10629
rect 13857 -10689 13887 -10669
rect 13837 -10729 13887 -10689
rect 13947 -10689 13977 -10669
rect 13947 -10729 13997 -10689
rect 13837 -10799 13997 -10729
rect 13837 -10839 13887 -10799
rect 13857 -10859 13887 -10839
rect 13947 -10839 13997 -10799
rect 13947 -10859 13977 -10839
rect 14057 -10899 14117 -10639
rect 13717 -10909 13797 -10899
rect 13717 -10969 13727 -10909
rect 13787 -10919 13797 -10909
rect 14037 -10909 14117 -10899
rect 14037 -10919 14047 -10909
rect 13787 -10969 14047 -10919
rect 14107 -10969 14117 -10909
rect 13717 -10979 14117 -10969
rect 14173 -10559 14573 -10549
rect 14173 -10619 14183 -10559
rect 14243 -10609 14503 -10559
rect 14243 -10619 14253 -10609
rect 14173 -10629 14253 -10619
rect 14493 -10619 14503 -10609
rect 14563 -10619 14573 -10559
rect 14493 -10629 14573 -10619
rect 14173 -10899 14233 -10629
rect 14503 -10639 14573 -10629
rect 14313 -10689 14343 -10669
rect 14293 -10729 14343 -10689
rect 14403 -10689 14433 -10669
rect 14403 -10729 14453 -10689
rect 14293 -10799 14453 -10729
rect 14293 -10839 14343 -10799
rect 14313 -10859 14343 -10839
rect 14403 -10839 14453 -10799
rect 14403 -10859 14433 -10839
rect 14513 -10899 14573 -10639
rect 14173 -10909 14253 -10899
rect 14173 -10969 14183 -10909
rect 14243 -10919 14253 -10909
rect 14493 -10909 14573 -10899
rect 14493 -10919 14503 -10909
rect 14243 -10969 14503 -10919
rect 14563 -10969 14573 -10909
rect 14173 -10979 14573 -10969
rect 14631 -10559 15031 -10549
rect 14631 -10619 14641 -10559
rect 14701 -10609 14961 -10559
rect 14701 -10619 14711 -10609
rect 14631 -10629 14711 -10619
rect 14951 -10619 14961 -10609
rect 15021 -10619 15031 -10559
rect 14951 -10629 15031 -10619
rect 14631 -10899 14691 -10629
rect 14961 -10639 15031 -10629
rect 14771 -10689 14801 -10669
rect 14751 -10729 14801 -10689
rect 14861 -10689 14891 -10669
rect 14861 -10729 14911 -10689
rect 14751 -10799 14911 -10729
rect 14751 -10839 14801 -10799
rect 14771 -10859 14801 -10839
rect 14861 -10839 14911 -10799
rect 14861 -10859 14891 -10839
rect 14971 -10899 15031 -10639
rect 14631 -10909 14711 -10899
rect 14631 -10969 14641 -10909
rect 14701 -10919 14711 -10909
rect 14951 -10909 15031 -10899
rect 14951 -10919 14961 -10909
rect 14701 -10969 14961 -10919
rect 15021 -10969 15031 -10909
rect 14631 -10979 15031 -10969
rect 15087 -10559 15487 -10549
rect 15087 -10619 15097 -10559
rect 15157 -10609 15417 -10559
rect 15157 -10619 15167 -10609
rect 15087 -10629 15167 -10619
rect 15407 -10619 15417 -10609
rect 15477 -10619 15487 -10559
rect 15407 -10629 15487 -10619
rect 15087 -10899 15147 -10629
rect 15417 -10639 15487 -10629
rect 15227 -10689 15257 -10669
rect 15207 -10729 15257 -10689
rect 15317 -10689 15347 -10669
rect 15317 -10729 15367 -10689
rect 15207 -10799 15367 -10729
rect 15207 -10839 15257 -10799
rect 15227 -10859 15257 -10839
rect 15317 -10839 15367 -10799
rect 15317 -10859 15347 -10839
rect 15427 -10899 15487 -10639
rect 15087 -10909 15167 -10899
rect 15087 -10969 15097 -10909
rect 15157 -10919 15167 -10909
rect 15407 -10909 15487 -10899
rect 15407 -10919 15417 -10909
rect 15157 -10969 15417 -10919
rect 15477 -10969 15487 -10909
rect 15087 -10979 15487 -10969
rect 1 -11051 401 -11041
rect 1 -11111 11 -11051
rect 71 -11101 331 -11051
rect 71 -11111 81 -11101
rect 1 -11121 81 -11111
rect 321 -11111 331 -11101
rect 391 -11111 401 -11051
rect 321 -11121 401 -11111
rect 1 -11391 61 -11121
rect 331 -11131 401 -11121
rect 141 -11181 171 -11161
rect 121 -11221 171 -11181
rect 231 -11181 261 -11161
rect 231 -11221 281 -11181
rect 121 -11291 281 -11221
rect 121 -11331 171 -11291
rect 141 -11351 171 -11331
rect 231 -11331 281 -11291
rect 231 -11351 261 -11331
rect 341 -11391 401 -11131
rect 1 -11401 81 -11391
rect 1 -11461 11 -11401
rect 71 -11411 81 -11401
rect 321 -11401 401 -11391
rect 321 -11411 331 -11401
rect 71 -11461 331 -11411
rect 391 -11461 401 -11401
rect 1 -11471 401 -11461
rect 457 -11051 857 -11041
rect 457 -11111 467 -11051
rect 527 -11101 787 -11051
rect 527 -11111 537 -11101
rect 457 -11121 537 -11111
rect 777 -11111 787 -11101
rect 847 -11111 857 -11051
rect 777 -11121 857 -11111
rect 457 -11391 517 -11121
rect 787 -11131 857 -11121
rect 597 -11181 627 -11161
rect 577 -11221 627 -11181
rect 687 -11181 717 -11161
rect 687 -11221 737 -11181
rect 577 -11291 737 -11221
rect 577 -11331 627 -11291
rect 597 -11351 627 -11331
rect 687 -11331 737 -11291
rect 687 -11351 717 -11331
rect 797 -11391 857 -11131
rect 457 -11401 537 -11391
rect 457 -11461 467 -11401
rect 527 -11411 537 -11401
rect 777 -11401 857 -11391
rect 777 -11411 787 -11401
rect 527 -11461 787 -11411
rect 847 -11461 857 -11401
rect 457 -11471 857 -11461
rect 913 -11051 1313 -11041
rect 913 -11111 923 -11051
rect 983 -11101 1243 -11051
rect 983 -11111 993 -11101
rect 913 -11121 993 -11111
rect 1233 -11111 1243 -11101
rect 1303 -11111 1313 -11051
rect 1233 -11121 1313 -11111
rect 913 -11391 973 -11121
rect 1243 -11131 1313 -11121
rect 1053 -11181 1083 -11161
rect 1033 -11221 1083 -11181
rect 1143 -11181 1173 -11161
rect 1143 -11221 1193 -11181
rect 1033 -11291 1193 -11221
rect 1033 -11331 1083 -11291
rect 1053 -11351 1083 -11331
rect 1143 -11331 1193 -11291
rect 1143 -11351 1173 -11331
rect 1253 -11391 1313 -11131
rect 913 -11401 993 -11391
rect 913 -11461 923 -11401
rect 983 -11411 993 -11401
rect 1233 -11401 1313 -11391
rect 1233 -11411 1243 -11401
rect 983 -11461 1243 -11411
rect 1303 -11461 1313 -11401
rect 913 -11471 1313 -11461
rect 1371 -11051 1771 -11041
rect 1371 -11111 1381 -11051
rect 1441 -11101 1701 -11051
rect 1441 -11111 1451 -11101
rect 1371 -11121 1451 -11111
rect 1691 -11111 1701 -11101
rect 1761 -11111 1771 -11051
rect 1691 -11121 1771 -11111
rect 1371 -11391 1431 -11121
rect 1701 -11131 1771 -11121
rect 1511 -11181 1541 -11161
rect 1491 -11221 1541 -11181
rect 1601 -11181 1631 -11161
rect 1601 -11221 1651 -11181
rect 1491 -11291 1651 -11221
rect 1491 -11331 1541 -11291
rect 1511 -11351 1541 -11331
rect 1601 -11331 1651 -11291
rect 1601 -11351 1631 -11331
rect 1711 -11391 1771 -11131
rect 1371 -11401 1451 -11391
rect 1371 -11461 1381 -11401
rect 1441 -11411 1451 -11401
rect 1691 -11401 1771 -11391
rect 1691 -11411 1701 -11401
rect 1441 -11461 1701 -11411
rect 1761 -11461 1771 -11401
rect 1371 -11471 1771 -11461
rect 1827 -11051 2227 -11041
rect 1827 -11111 1837 -11051
rect 1897 -11101 2157 -11051
rect 1897 -11111 1907 -11101
rect 1827 -11121 1907 -11111
rect 2147 -11111 2157 -11101
rect 2217 -11111 2227 -11051
rect 2147 -11121 2227 -11111
rect 1827 -11391 1887 -11121
rect 2157 -11131 2227 -11121
rect 1967 -11181 1997 -11161
rect 1947 -11221 1997 -11181
rect 2057 -11181 2087 -11161
rect 2057 -11221 2107 -11181
rect 1947 -11291 2107 -11221
rect 1947 -11331 1997 -11291
rect 1967 -11351 1997 -11331
rect 2057 -11331 2107 -11291
rect 2057 -11351 2087 -11331
rect 2167 -11391 2227 -11131
rect 1827 -11401 1907 -11391
rect 1827 -11461 1837 -11401
rect 1897 -11411 1907 -11401
rect 2147 -11401 2227 -11391
rect 2147 -11411 2157 -11401
rect 1897 -11461 2157 -11411
rect 2217 -11461 2227 -11401
rect 1827 -11471 2227 -11461
rect 2283 -11051 2683 -11041
rect 2283 -11111 2293 -11051
rect 2353 -11101 2613 -11051
rect 2353 -11111 2363 -11101
rect 2283 -11121 2363 -11111
rect 2603 -11111 2613 -11101
rect 2673 -11111 2683 -11051
rect 2603 -11121 2683 -11111
rect 2283 -11391 2343 -11121
rect 2613 -11131 2683 -11121
rect 2423 -11181 2453 -11161
rect 2403 -11221 2453 -11181
rect 2513 -11181 2543 -11161
rect 2513 -11221 2563 -11181
rect 2403 -11291 2563 -11221
rect 2403 -11331 2453 -11291
rect 2423 -11351 2453 -11331
rect 2513 -11331 2563 -11291
rect 2513 -11351 2543 -11331
rect 2623 -11391 2683 -11131
rect 2283 -11401 2363 -11391
rect 2283 -11461 2293 -11401
rect 2353 -11411 2363 -11401
rect 2603 -11401 2683 -11391
rect 2603 -11411 2613 -11401
rect 2353 -11461 2613 -11411
rect 2673 -11461 2683 -11401
rect 2283 -11471 2683 -11461
rect 2741 -11051 3141 -11041
rect 2741 -11111 2751 -11051
rect 2811 -11101 3071 -11051
rect 2811 -11111 2821 -11101
rect 2741 -11121 2821 -11111
rect 3061 -11111 3071 -11101
rect 3131 -11111 3141 -11051
rect 3061 -11121 3141 -11111
rect 2741 -11391 2801 -11121
rect 3071 -11131 3141 -11121
rect 2881 -11181 2911 -11161
rect 2861 -11221 2911 -11181
rect 2971 -11181 3001 -11161
rect 2971 -11221 3021 -11181
rect 2861 -11291 3021 -11221
rect 2861 -11331 2911 -11291
rect 2881 -11351 2911 -11331
rect 2971 -11331 3021 -11291
rect 2971 -11351 3001 -11331
rect 3081 -11391 3141 -11131
rect 2741 -11401 2821 -11391
rect 2741 -11461 2751 -11401
rect 2811 -11411 2821 -11401
rect 3061 -11401 3141 -11391
rect 3061 -11411 3071 -11401
rect 2811 -11461 3071 -11411
rect 3131 -11461 3141 -11401
rect 2741 -11471 3141 -11461
rect 3197 -11051 3597 -11041
rect 3197 -11111 3207 -11051
rect 3267 -11101 3527 -11051
rect 3267 -11111 3277 -11101
rect 3197 -11121 3277 -11111
rect 3517 -11111 3527 -11101
rect 3587 -11111 3597 -11051
rect 3517 -11121 3597 -11111
rect 3197 -11391 3257 -11121
rect 3527 -11131 3597 -11121
rect 3337 -11181 3367 -11161
rect 3317 -11221 3367 -11181
rect 3427 -11181 3457 -11161
rect 3427 -11221 3477 -11181
rect 3317 -11291 3477 -11221
rect 3317 -11331 3367 -11291
rect 3337 -11351 3367 -11331
rect 3427 -11331 3477 -11291
rect 3427 -11351 3457 -11331
rect 3537 -11391 3597 -11131
rect 3197 -11401 3277 -11391
rect 3197 -11461 3207 -11401
rect 3267 -11411 3277 -11401
rect 3517 -11401 3597 -11391
rect 3517 -11411 3527 -11401
rect 3267 -11461 3527 -11411
rect 3587 -11461 3597 -11401
rect 3197 -11471 3597 -11461
rect 3653 -11051 4053 -11041
rect 3653 -11111 3663 -11051
rect 3723 -11101 3983 -11051
rect 3723 -11111 3733 -11101
rect 3653 -11121 3733 -11111
rect 3973 -11111 3983 -11101
rect 4043 -11111 4053 -11051
rect 3973 -11121 4053 -11111
rect 3653 -11391 3713 -11121
rect 3983 -11131 4053 -11121
rect 3793 -11181 3823 -11161
rect 3773 -11221 3823 -11181
rect 3883 -11181 3913 -11161
rect 3883 -11221 3933 -11181
rect 3773 -11291 3933 -11221
rect 3773 -11331 3823 -11291
rect 3793 -11351 3823 -11331
rect 3883 -11331 3933 -11291
rect 3883 -11351 3913 -11331
rect 3993 -11391 4053 -11131
rect 3653 -11401 3733 -11391
rect 3653 -11461 3663 -11401
rect 3723 -11411 3733 -11401
rect 3973 -11401 4053 -11391
rect 3973 -11411 3983 -11401
rect 3723 -11461 3983 -11411
rect 4043 -11461 4053 -11401
rect 3653 -11471 4053 -11461
rect 4111 -11051 4511 -11041
rect 4111 -11111 4121 -11051
rect 4181 -11101 4441 -11051
rect 4181 -11111 4191 -11101
rect 4111 -11121 4191 -11111
rect 4431 -11111 4441 -11101
rect 4501 -11111 4511 -11051
rect 4431 -11121 4511 -11111
rect 4111 -11391 4171 -11121
rect 4441 -11131 4511 -11121
rect 4251 -11181 4281 -11161
rect 4231 -11221 4281 -11181
rect 4341 -11181 4371 -11161
rect 4341 -11221 4391 -11181
rect 4231 -11291 4391 -11221
rect 4231 -11331 4281 -11291
rect 4251 -11351 4281 -11331
rect 4341 -11331 4391 -11291
rect 4341 -11351 4371 -11331
rect 4451 -11391 4511 -11131
rect 4111 -11401 4191 -11391
rect 4111 -11461 4121 -11401
rect 4181 -11411 4191 -11401
rect 4431 -11401 4511 -11391
rect 4431 -11411 4441 -11401
rect 4181 -11461 4441 -11411
rect 4501 -11461 4511 -11401
rect 4111 -11471 4511 -11461
rect 4567 -11051 4967 -11041
rect 4567 -11111 4577 -11051
rect 4637 -11101 4897 -11051
rect 4637 -11111 4647 -11101
rect 4567 -11121 4647 -11111
rect 4887 -11111 4897 -11101
rect 4957 -11111 4967 -11051
rect 4887 -11121 4967 -11111
rect 4567 -11391 4627 -11121
rect 4897 -11131 4967 -11121
rect 4707 -11181 4737 -11161
rect 4687 -11221 4737 -11181
rect 4797 -11181 4827 -11161
rect 4797 -11221 4847 -11181
rect 4687 -11291 4847 -11221
rect 4687 -11331 4737 -11291
rect 4707 -11351 4737 -11331
rect 4797 -11331 4847 -11291
rect 4797 -11351 4827 -11331
rect 4907 -11391 4967 -11131
rect 4567 -11401 4647 -11391
rect 4567 -11461 4577 -11401
rect 4637 -11411 4647 -11401
rect 4887 -11401 4967 -11391
rect 4887 -11411 4897 -11401
rect 4637 -11461 4897 -11411
rect 4957 -11461 4967 -11401
rect 4567 -11471 4967 -11461
rect 5023 -11051 5423 -11041
rect 5023 -11111 5033 -11051
rect 5093 -11101 5353 -11051
rect 5093 -11111 5103 -11101
rect 5023 -11121 5103 -11111
rect 5343 -11111 5353 -11101
rect 5413 -11111 5423 -11051
rect 5343 -11121 5423 -11111
rect 5023 -11391 5083 -11121
rect 5353 -11131 5423 -11121
rect 5163 -11181 5193 -11161
rect 5143 -11221 5193 -11181
rect 5253 -11181 5283 -11161
rect 5253 -11221 5303 -11181
rect 5143 -11291 5303 -11221
rect 5143 -11331 5193 -11291
rect 5163 -11351 5193 -11331
rect 5253 -11331 5303 -11291
rect 5253 -11351 5283 -11331
rect 5363 -11391 5423 -11131
rect 5023 -11401 5103 -11391
rect 5023 -11461 5033 -11401
rect 5093 -11411 5103 -11401
rect 5343 -11401 5423 -11391
rect 5343 -11411 5353 -11401
rect 5093 -11461 5353 -11411
rect 5413 -11461 5423 -11401
rect 5023 -11471 5423 -11461
rect 5481 -11051 5881 -11041
rect 5481 -11111 5491 -11051
rect 5551 -11101 5811 -11051
rect 5551 -11111 5561 -11101
rect 5481 -11121 5561 -11111
rect 5801 -11111 5811 -11101
rect 5871 -11111 5881 -11051
rect 5801 -11121 5881 -11111
rect 5481 -11391 5541 -11121
rect 5811 -11131 5881 -11121
rect 5621 -11181 5651 -11161
rect 5601 -11221 5651 -11181
rect 5711 -11181 5741 -11161
rect 5711 -11221 5761 -11181
rect 5601 -11291 5761 -11221
rect 5601 -11331 5651 -11291
rect 5621 -11351 5651 -11331
rect 5711 -11331 5761 -11291
rect 5711 -11351 5741 -11331
rect 5821 -11391 5881 -11131
rect 5481 -11401 5561 -11391
rect 5481 -11461 5491 -11401
rect 5551 -11411 5561 -11401
rect 5801 -11401 5881 -11391
rect 5801 -11411 5811 -11401
rect 5551 -11461 5811 -11411
rect 5871 -11461 5881 -11401
rect 5481 -11471 5881 -11461
rect 5937 -11051 6337 -11041
rect 5937 -11111 5947 -11051
rect 6007 -11101 6267 -11051
rect 6007 -11111 6017 -11101
rect 5937 -11121 6017 -11111
rect 6257 -11111 6267 -11101
rect 6327 -11111 6337 -11051
rect 6257 -11121 6337 -11111
rect 5937 -11391 5997 -11121
rect 6267 -11131 6337 -11121
rect 6077 -11181 6107 -11161
rect 6057 -11221 6107 -11181
rect 6167 -11181 6197 -11161
rect 6167 -11221 6217 -11181
rect 6057 -11291 6217 -11221
rect 6057 -11331 6107 -11291
rect 6077 -11351 6107 -11331
rect 6167 -11331 6217 -11291
rect 6167 -11351 6197 -11331
rect 6277 -11391 6337 -11131
rect 5937 -11401 6017 -11391
rect 5937 -11461 5947 -11401
rect 6007 -11411 6017 -11401
rect 6257 -11401 6337 -11391
rect 6257 -11411 6267 -11401
rect 6007 -11461 6267 -11411
rect 6327 -11461 6337 -11401
rect 5937 -11471 6337 -11461
rect 6393 -11051 6793 -11041
rect 6393 -11111 6403 -11051
rect 6463 -11101 6723 -11051
rect 6463 -11111 6473 -11101
rect 6393 -11121 6473 -11111
rect 6713 -11111 6723 -11101
rect 6783 -11111 6793 -11051
rect 6713 -11121 6793 -11111
rect 6393 -11391 6453 -11121
rect 6723 -11131 6793 -11121
rect 6533 -11181 6563 -11161
rect 6513 -11221 6563 -11181
rect 6623 -11181 6653 -11161
rect 6623 -11221 6673 -11181
rect 6513 -11291 6673 -11221
rect 6513 -11331 6563 -11291
rect 6533 -11351 6563 -11331
rect 6623 -11331 6673 -11291
rect 6623 -11351 6653 -11331
rect 6733 -11391 6793 -11131
rect 6393 -11401 6473 -11391
rect 6393 -11461 6403 -11401
rect 6463 -11411 6473 -11401
rect 6713 -11401 6793 -11391
rect 6713 -11411 6723 -11401
rect 6463 -11461 6723 -11411
rect 6783 -11461 6793 -11401
rect 6393 -11471 6793 -11461
rect 6851 -11051 7251 -11041
rect 6851 -11111 6861 -11051
rect 6921 -11101 7181 -11051
rect 6921 -11111 6931 -11101
rect 6851 -11121 6931 -11111
rect 7171 -11111 7181 -11101
rect 7241 -11111 7251 -11051
rect 7171 -11121 7251 -11111
rect 6851 -11391 6911 -11121
rect 7181 -11131 7251 -11121
rect 6991 -11181 7021 -11161
rect 6971 -11221 7021 -11181
rect 7081 -11181 7111 -11161
rect 7081 -11221 7131 -11181
rect 6971 -11291 7131 -11221
rect 6971 -11331 7021 -11291
rect 6991 -11351 7021 -11331
rect 7081 -11331 7131 -11291
rect 7081 -11351 7111 -11331
rect 7191 -11391 7251 -11131
rect 6851 -11401 6931 -11391
rect 6851 -11461 6861 -11401
rect 6921 -11411 6931 -11401
rect 7171 -11401 7251 -11391
rect 7171 -11411 7181 -11401
rect 6921 -11461 7181 -11411
rect 7241 -11461 7251 -11401
rect 6851 -11471 7251 -11461
rect 7307 -11051 7707 -11041
rect 7307 -11111 7317 -11051
rect 7377 -11101 7637 -11051
rect 7377 -11111 7387 -11101
rect 7307 -11121 7387 -11111
rect 7627 -11111 7637 -11101
rect 7697 -11111 7707 -11051
rect 7627 -11121 7707 -11111
rect 7307 -11391 7367 -11121
rect 7637 -11131 7707 -11121
rect 7447 -11181 7477 -11161
rect 7427 -11221 7477 -11181
rect 7537 -11181 7567 -11161
rect 7537 -11221 7587 -11181
rect 7427 -11291 7587 -11221
rect 7427 -11331 7477 -11291
rect 7447 -11351 7477 -11331
rect 7537 -11331 7587 -11291
rect 7537 -11351 7567 -11331
rect 7647 -11391 7707 -11131
rect 7307 -11401 7387 -11391
rect 7307 -11461 7317 -11401
rect 7377 -11411 7387 -11401
rect 7627 -11401 7707 -11391
rect 7627 -11411 7637 -11401
rect 7377 -11461 7637 -11411
rect 7697 -11461 7707 -11401
rect 7307 -11471 7707 -11461
rect 7763 -11051 8163 -11041
rect 7763 -11111 7773 -11051
rect 7833 -11101 8093 -11051
rect 7833 -11111 7843 -11101
rect 7763 -11121 7843 -11111
rect 8083 -11111 8093 -11101
rect 8153 -11111 8163 -11051
rect 8083 -11121 8163 -11111
rect 7763 -11391 7823 -11121
rect 8093 -11131 8163 -11121
rect 7903 -11181 7933 -11161
rect 7883 -11221 7933 -11181
rect 7993 -11181 8023 -11161
rect 7993 -11221 8043 -11181
rect 7883 -11291 8043 -11221
rect 7883 -11331 7933 -11291
rect 7903 -11351 7933 -11331
rect 7993 -11331 8043 -11291
rect 7993 -11351 8023 -11331
rect 8103 -11391 8163 -11131
rect 7763 -11401 7843 -11391
rect 7763 -11461 7773 -11401
rect 7833 -11411 7843 -11401
rect 8083 -11401 8163 -11391
rect 8083 -11411 8093 -11401
rect 7833 -11461 8093 -11411
rect 8153 -11461 8163 -11401
rect 7763 -11471 8163 -11461
rect 8237 -11051 8637 -11041
rect 8237 -11111 8247 -11051
rect 8307 -11101 8567 -11051
rect 8307 -11111 8317 -11101
rect 8237 -11121 8317 -11111
rect 8557 -11111 8567 -11101
rect 8627 -11111 8637 -11051
rect 8557 -11121 8637 -11111
rect 8237 -11391 8297 -11121
rect 8567 -11131 8637 -11121
rect 8377 -11181 8407 -11161
rect 8357 -11221 8407 -11181
rect 8467 -11181 8497 -11161
rect 8467 -11221 8517 -11181
rect 8357 -11291 8517 -11221
rect 8357 -11331 8407 -11291
rect 8377 -11351 8407 -11331
rect 8467 -11331 8517 -11291
rect 8467 -11351 8497 -11331
rect 8577 -11391 8637 -11131
rect 8237 -11401 8317 -11391
rect 8237 -11461 8247 -11401
rect 8307 -11411 8317 -11401
rect 8557 -11401 8637 -11391
rect 8557 -11411 8567 -11401
rect 8307 -11461 8567 -11411
rect 8627 -11461 8637 -11401
rect 8237 -11471 8637 -11461
rect 8693 -11051 9093 -11041
rect 8693 -11111 8703 -11051
rect 8763 -11101 9023 -11051
rect 8763 -11111 8773 -11101
rect 8693 -11121 8773 -11111
rect 9013 -11111 9023 -11101
rect 9083 -11111 9093 -11051
rect 9013 -11121 9093 -11111
rect 8693 -11391 8753 -11121
rect 9023 -11131 9093 -11121
rect 8833 -11181 8863 -11161
rect 8813 -11221 8863 -11181
rect 8923 -11181 8953 -11161
rect 8923 -11221 8973 -11181
rect 8813 -11291 8973 -11221
rect 8813 -11331 8863 -11291
rect 8833 -11351 8863 -11331
rect 8923 -11331 8973 -11291
rect 8923 -11351 8953 -11331
rect 9033 -11391 9093 -11131
rect 8693 -11401 8773 -11391
rect 8693 -11461 8703 -11401
rect 8763 -11411 8773 -11401
rect 9013 -11401 9093 -11391
rect 9013 -11411 9023 -11401
rect 8763 -11461 9023 -11411
rect 9083 -11461 9093 -11401
rect 8693 -11471 9093 -11461
rect 9151 -11051 9551 -11041
rect 9151 -11111 9161 -11051
rect 9221 -11101 9481 -11051
rect 9221 -11111 9231 -11101
rect 9151 -11121 9231 -11111
rect 9471 -11111 9481 -11101
rect 9541 -11111 9551 -11051
rect 9471 -11121 9551 -11111
rect 9151 -11391 9211 -11121
rect 9481 -11131 9551 -11121
rect 9291 -11181 9321 -11161
rect 9271 -11221 9321 -11181
rect 9381 -11181 9411 -11161
rect 9491 -11170 9551 -11131
rect 9607 -11051 10007 -11041
rect 9607 -11111 9617 -11051
rect 9677 -11101 9937 -11051
rect 9677 -11111 9687 -11101
rect 9607 -11121 9687 -11111
rect 9927 -11111 9937 -11101
rect 9997 -11111 10007 -11051
rect 9927 -11121 10007 -11111
rect 9381 -11221 9431 -11181
rect 9271 -11291 9431 -11221
rect 9271 -11331 9321 -11291
rect 9291 -11351 9321 -11331
rect 9381 -11331 9431 -11291
rect 9381 -11351 9411 -11331
rect 9491 -11391 9550 -11170
rect 9151 -11401 9231 -11391
rect 9151 -11461 9161 -11401
rect 9221 -11411 9231 -11401
rect 9471 -11401 9550 -11391
rect 9471 -11411 9481 -11401
rect 9221 -11461 9481 -11411
rect 9541 -11461 9550 -11401
rect 9151 -11471 9550 -11461
rect 9607 -11391 9667 -11121
rect 9937 -11131 10007 -11121
rect 9747 -11181 9777 -11161
rect 9727 -11221 9777 -11181
rect 9837 -11181 9867 -11161
rect 9837 -11221 9887 -11181
rect 9727 -11291 9887 -11221
rect 9727 -11331 9777 -11291
rect 9747 -11351 9777 -11331
rect 9837 -11331 9887 -11291
rect 9837 -11351 9867 -11331
rect 9947 -11391 10007 -11131
rect 9607 -11401 9687 -11391
rect 9607 -11461 9617 -11401
rect 9677 -11411 9687 -11401
rect 9927 -11401 10007 -11391
rect 9927 -11411 9937 -11401
rect 9677 -11461 9937 -11411
rect 9997 -11461 10007 -11401
rect 9607 -11471 10007 -11461
rect 10063 -11051 10463 -11041
rect 10063 -11111 10073 -11051
rect 10133 -11101 10393 -11051
rect 10133 -11111 10143 -11101
rect 10063 -11121 10143 -11111
rect 10383 -11111 10393 -11101
rect 10453 -11111 10463 -11051
rect 10383 -11121 10463 -11111
rect 10063 -11391 10123 -11121
rect 10393 -11131 10463 -11121
rect 10203 -11181 10233 -11161
rect 10183 -11221 10233 -11181
rect 10293 -11181 10323 -11161
rect 10293 -11221 10343 -11181
rect 10183 -11291 10343 -11221
rect 10183 -11331 10233 -11291
rect 10203 -11351 10233 -11331
rect 10293 -11331 10343 -11291
rect 10293 -11351 10323 -11331
rect 10403 -11391 10463 -11131
rect 10063 -11401 10143 -11391
rect 10063 -11461 10073 -11401
rect 10133 -11411 10143 -11401
rect 10383 -11401 10463 -11391
rect 10383 -11411 10393 -11401
rect 10133 -11461 10393 -11411
rect 10453 -11461 10463 -11401
rect 10063 -11471 10463 -11461
rect 10521 -11051 10921 -11041
rect 10521 -11111 10531 -11051
rect 10591 -11101 10851 -11051
rect 10591 -11111 10601 -11101
rect 10521 -11121 10601 -11111
rect 10841 -11111 10851 -11101
rect 10911 -11111 10921 -11051
rect 10841 -11121 10921 -11111
rect 10521 -11391 10581 -11121
rect 10851 -11131 10921 -11121
rect 10661 -11181 10691 -11161
rect 10641 -11221 10691 -11181
rect 10751 -11181 10781 -11161
rect 10751 -11221 10801 -11181
rect 10641 -11291 10801 -11221
rect 10641 -11331 10691 -11291
rect 10661 -11351 10691 -11331
rect 10751 -11331 10801 -11291
rect 10751 -11351 10781 -11331
rect 10861 -11391 10921 -11131
rect 10521 -11401 10601 -11391
rect 10521 -11461 10531 -11401
rect 10591 -11411 10601 -11401
rect 10841 -11401 10921 -11391
rect 10841 -11411 10851 -11401
rect 10591 -11461 10851 -11411
rect 10911 -11461 10921 -11401
rect 10521 -11471 10921 -11461
rect 10977 -11051 11377 -11041
rect 10977 -11111 10987 -11051
rect 11047 -11101 11307 -11051
rect 11047 -11111 11057 -11101
rect 10977 -11121 11057 -11111
rect 11297 -11111 11307 -11101
rect 11367 -11111 11377 -11051
rect 11297 -11121 11377 -11111
rect 10977 -11391 11037 -11121
rect 11307 -11131 11377 -11121
rect 11117 -11181 11147 -11161
rect 11097 -11221 11147 -11181
rect 11207 -11181 11237 -11161
rect 11207 -11221 11257 -11181
rect 11097 -11291 11257 -11221
rect 11097 -11331 11147 -11291
rect 11117 -11351 11147 -11331
rect 11207 -11331 11257 -11291
rect 11207 -11351 11237 -11331
rect 11317 -11391 11377 -11131
rect 10977 -11401 11057 -11391
rect 10977 -11461 10987 -11401
rect 11047 -11411 11057 -11401
rect 11297 -11401 11377 -11391
rect 11297 -11411 11307 -11401
rect 11047 -11461 11307 -11411
rect 11367 -11461 11377 -11401
rect 10977 -11471 11377 -11461
rect 11433 -11051 11833 -11041
rect 11433 -11111 11443 -11051
rect 11503 -11101 11763 -11051
rect 11503 -11111 11513 -11101
rect 11433 -11121 11513 -11111
rect 11753 -11111 11763 -11101
rect 11823 -11111 11833 -11051
rect 11753 -11121 11833 -11111
rect 11433 -11391 11493 -11121
rect 11763 -11131 11833 -11121
rect 11573 -11181 11603 -11161
rect 11553 -11221 11603 -11181
rect 11663 -11181 11693 -11161
rect 11663 -11221 11713 -11181
rect 11553 -11291 11713 -11221
rect 11553 -11331 11603 -11291
rect 11573 -11351 11603 -11331
rect 11663 -11331 11713 -11291
rect 11663 -11351 11693 -11331
rect 11773 -11391 11833 -11131
rect 11433 -11401 11513 -11391
rect 11433 -11461 11443 -11401
rect 11503 -11411 11513 -11401
rect 11753 -11401 11833 -11391
rect 11753 -11411 11763 -11401
rect 11503 -11461 11763 -11411
rect 11823 -11461 11833 -11401
rect 11433 -11471 11833 -11461
rect 11891 -11051 12291 -11041
rect 11891 -11111 11901 -11051
rect 11961 -11101 12221 -11051
rect 11961 -11111 11971 -11101
rect 11891 -11121 11971 -11111
rect 12211 -11111 12221 -11101
rect 12281 -11111 12291 -11051
rect 12211 -11121 12291 -11111
rect 11891 -11391 11951 -11121
rect 12221 -11131 12291 -11121
rect 12031 -11181 12061 -11161
rect 12011 -11221 12061 -11181
rect 12121 -11181 12151 -11161
rect 12121 -11221 12171 -11181
rect 12011 -11291 12171 -11221
rect 12011 -11331 12061 -11291
rect 12031 -11351 12061 -11331
rect 12121 -11331 12171 -11291
rect 12121 -11351 12151 -11331
rect 12231 -11391 12291 -11131
rect 11891 -11401 11971 -11391
rect 11891 -11461 11901 -11401
rect 11961 -11411 11971 -11401
rect 12211 -11401 12291 -11391
rect 12211 -11411 12221 -11401
rect 11961 -11461 12221 -11411
rect 12281 -11461 12291 -11401
rect 11891 -11471 12291 -11461
rect 12347 -11051 12747 -11041
rect 12347 -11111 12357 -11051
rect 12417 -11101 12677 -11051
rect 12417 -11111 12427 -11101
rect 12347 -11121 12427 -11111
rect 12667 -11111 12677 -11101
rect 12737 -11111 12747 -11051
rect 12667 -11121 12747 -11111
rect 12347 -11391 12407 -11121
rect 12677 -11131 12747 -11121
rect 12487 -11181 12517 -11161
rect 12467 -11221 12517 -11181
rect 12577 -11181 12607 -11161
rect 12577 -11221 12627 -11181
rect 12467 -11291 12627 -11221
rect 12467 -11331 12517 -11291
rect 12487 -11351 12517 -11331
rect 12577 -11331 12627 -11291
rect 12577 -11351 12607 -11331
rect 12687 -11391 12747 -11131
rect 12347 -11401 12427 -11391
rect 12347 -11461 12357 -11401
rect 12417 -11411 12427 -11401
rect 12667 -11401 12747 -11391
rect 12667 -11411 12677 -11401
rect 12417 -11461 12677 -11411
rect 12737 -11461 12747 -11401
rect 12347 -11471 12747 -11461
rect 12803 -11051 13203 -11041
rect 12803 -11111 12813 -11051
rect 12873 -11101 13133 -11051
rect 12873 -11111 12883 -11101
rect 12803 -11121 12883 -11111
rect 13123 -11111 13133 -11101
rect 13193 -11111 13203 -11051
rect 13123 -11121 13203 -11111
rect 12803 -11391 12863 -11121
rect 13133 -11131 13203 -11121
rect 12943 -11181 12973 -11161
rect 12923 -11221 12973 -11181
rect 13033 -11181 13063 -11161
rect 13033 -11221 13083 -11181
rect 12923 -11291 13083 -11221
rect 12923 -11331 12973 -11291
rect 12943 -11351 12973 -11331
rect 13033 -11331 13083 -11291
rect 13033 -11351 13063 -11331
rect 13143 -11391 13203 -11131
rect 12803 -11401 12883 -11391
rect 12803 -11461 12813 -11401
rect 12873 -11411 12883 -11401
rect 13123 -11401 13203 -11391
rect 13123 -11411 13133 -11401
rect 12873 -11461 13133 -11411
rect 13193 -11461 13203 -11401
rect 12803 -11471 13203 -11461
rect 13261 -11051 13661 -11041
rect 13261 -11111 13271 -11051
rect 13331 -11101 13591 -11051
rect 13331 -11111 13341 -11101
rect 13261 -11121 13341 -11111
rect 13581 -11111 13591 -11101
rect 13651 -11111 13661 -11051
rect 13581 -11121 13661 -11111
rect 13261 -11391 13321 -11121
rect 13591 -11131 13661 -11121
rect 13401 -11181 13431 -11161
rect 13381 -11221 13431 -11181
rect 13491 -11181 13521 -11161
rect 13491 -11221 13541 -11181
rect 13381 -11291 13541 -11221
rect 13381 -11331 13431 -11291
rect 13401 -11351 13431 -11331
rect 13491 -11331 13541 -11291
rect 13491 -11351 13521 -11331
rect 13601 -11391 13661 -11131
rect 13261 -11401 13341 -11391
rect 13261 -11461 13271 -11401
rect 13331 -11411 13341 -11401
rect 13581 -11401 13661 -11391
rect 13581 -11411 13591 -11401
rect 13331 -11461 13591 -11411
rect 13651 -11461 13661 -11401
rect 13261 -11471 13661 -11461
rect 13717 -11051 14117 -11041
rect 13717 -11111 13727 -11051
rect 13787 -11101 14047 -11051
rect 13787 -11111 13797 -11101
rect 13717 -11121 13797 -11111
rect 14037 -11111 14047 -11101
rect 14107 -11111 14117 -11051
rect 14037 -11121 14117 -11111
rect 13717 -11391 13777 -11121
rect 14047 -11131 14117 -11121
rect 13857 -11181 13887 -11161
rect 13837 -11221 13887 -11181
rect 13947 -11181 13977 -11161
rect 13947 -11221 13997 -11181
rect 13837 -11291 13997 -11221
rect 13837 -11331 13887 -11291
rect 13857 -11351 13887 -11331
rect 13947 -11331 13997 -11291
rect 13947 -11351 13977 -11331
rect 14057 -11391 14117 -11131
rect 13717 -11401 13797 -11391
rect 13717 -11461 13727 -11401
rect 13787 -11411 13797 -11401
rect 14037 -11401 14117 -11391
rect 14037 -11411 14047 -11401
rect 13787 -11461 14047 -11411
rect 14107 -11461 14117 -11401
rect 13717 -11471 14117 -11461
rect 14173 -11051 14573 -11041
rect 14173 -11111 14183 -11051
rect 14243 -11101 14503 -11051
rect 14243 -11111 14253 -11101
rect 14173 -11121 14253 -11111
rect 14493 -11111 14503 -11101
rect 14563 -11111 14573 -11051
rect 14493 -11121 14573 -11111
rect 14173 -11391 14233 -11121
rect 14503 -11131 14573 -11121
rect 14313 -11181 14343 -11161
rect 14293 -11221 14343 -11181
rect 14403 -11181 14433 -11161
rect 14403 -11221 14453 -11181
rect 14293 -11291 14453 -11221
rect 14293 -11331 14343 -11291
rect 14313 -11351 14343 -11331
rect 14403 -11331 14453 -11291
rect 14403 -11351 14433 -11331
rect 14513 -11391 14573 -11131
rect 14173 -11401 14253 -11391
rect 14173 -11461 14183 -11401
rect 14243 -11411 14253 -11401
rect 14493 -11401 14573 -11391
rect 14493 -11411 14503 -11401
rect 14243 -11461 14503 -11411
rect 14563 -11461 14573 -11401
rect 14173 -11471 14573 -11461
rect 14631 -11051 15031 -11041
rect 14631 -11111 14641 -11051
rect 14701 -11101 14961 -11051
rect 14701 -11111 14711 -11101
rect 14631 -11121 14711 -11111
rect 14951 -11111 14961 -11101
rect 15021 -11111 15031 -11051
rect 14951 -11121 15031 -11111
rect 14631 -11391 14691 -11121
rect 14961 -11131 15031 -11121
rect 14771 -11181 14801 -11161
rect 14751 -11221 14801 -11181
rect 14861 -11181 14891 -11161
rect 14861 -11221 14911 -11181
rect 14751 -11291 14911 -11221
rect 14751 -11331 14801 -11291
rect 14771 -11351 14801 -11331
rect 14861 -11331 14911 -11291
rect 14861 -11351 14891 -11331
rect 14971 -11391 15031 -11131
rect 14631 -11401 14711 -11391
rect 14631 -11461 14641 -11401
rect 14701 -11411 14711 -11401
rect 14951 -11401 15031 -11391
rect 14951 -11411 14961 -11401
rect 14701 -11461 14961 -11411
rect 15021 -11461 15031 -11401
rect 14631 -11471 15031 -11461
rect 15087 -11051 15487 -11041
rect 15087 -11111 15097 -11051
rect 15157 -11101 15417 -11051
rect 15157 -11111 15167 -11101
rect 15087 -11121 15167 -11111
rect 15407 -11111 15417 -11101
rect 15477 -11111 15487 -11051
rect 15407 -11121 15487 -11111
rect 15087 -11391 15147 -11121
rect 15417 -11131 15487 -11121
rect 15227 -11181 15257 -11161
rect 15207 -11221 15257 -11181
rect 15317 -11181 15347 -11161
rect 15317 -11221 15367 -11181
rect 15207 -11291 15367 -11221
rect 15207 -11331 15257 -11291
rect 15227 -11351 15257 -11331
rect 15317 -11331 15367 -11291
rect 15317 -11351 15347 -11331
rect 15427 -11391 15487 -11131
rect 15087 -11401 15167 -11391
rect 15087 -11461 15097 -11401
rect 15157 -11411 15167 -11401
rect 15407 -11401 15487 -11391
rect 15407 -11411 15417 -11401
rect 15157 -11461 15417 -11411
rect 15477 -11461 15487 -11401
rect 15087 -11471 15487 -11461
rect 0 -11544 400 -11534
rect 0 -11604 10 -11544
rect 70 -11594 330 -11544
rect 70 -11604 80 -11594
rect 0 -11614 80 -11604
rect 320 -11604 330 -11594
rect 390 -11604 400 -11544
rect 320 -11614 400 -11604
rect 0 -11884 60 -11614
rect 330 -11624 400 -11614
rect 140 -11674 170 -11654
rect 120 -11714 170 -11674
rect 230 -11674 260 -11654
rect 230 -11714 280 -11674
rect 120 -11784 280 -11714
rect 120 -11824 170 -11784
rect 140 -11844 170 -11824
rect 230 -11824 280 -11784
rect 230 -11844 260 -11824
rect 340 -11884 400 -11624
rect 0 -11894 80 -11884
rect 0 -11954 10 -11894
rect 70 -11904 80 -11894
rect 320 -11894 400 -11884
rect 320 -11904 330 -11894
rect 70 -11954 330 -11904
rect 390 -11954 400 -11894
rect 0 -11964 400 -11954
rect 456 -11544 856 -11534
rect 456 -11604 466 -11544
rect 526 -11594 786 -11544
rect 526 -11604 536 -11594
rect 456 -11614 536 -11604
rect 776 -11604 786 -11594
rect 846 -11604 856 -11544
rect 776 -11614 856 -11604
rect 456 -11884 516 -11614
rect 786 -11624 856 -11614
rect 596 -11674 626 -11654
rect 576 -11714 626 -11674
rect 686 -11674 716 -11654
rect 686 -11714 736 -11674
rect 576 -11784 736 -11714
rect 576 -11824 626 -11784
rect 596 -11844 626 -11824
rect 686 -11824 736 -11784
rect 686 -11844 716 -11824
rect 796 -11884 856 -11624
rect 456 -11894 536 -11884
rect 456 -11954 466 -11894
rect 526 -11904 536 -11894
rect 776 -11894 856 -11884
rect 776 -11904 786 -11894
rect 526 -11954 786 -11904
rect 846 -11954 856 -11894
rect 456 -11964 856 -11954
rect 912 -11544 1312 -11534
rect 912 -11604 922 -11544
rect 982 -11594 1242 -11544
rect 982 -11604 992 -11594
rect 912 -11614 992 -11604
rect 1232 -11604 1242 -11594
rect 1302 -11604 1312 -11544
rect 1232 -11614 1312 -11604
rect 912 -11884 972 -11614
rect 1242 -11624 1312 -11614
rect 1052 -11674 1082 -11654
rect 1032 -11714 1082 -11674
rect 1142 -11674 1172 -11654
rect 1142 -11714 1192 -11674
rect 1032 -11784 1192 -11714
rect 1032 -11824 1082 -11784
rect 1052 -11844 1082 -11824
rect 1142 -11824 1192 -11784
rect 1142 -11844 1172 -11824
rect 1252 -11884 1312 -11624
rect 912 -11894 992 -11884
rect 912 -11954 922 -11894
rect 982 -11904 992 -11894
rect 1232 -11894 1312 -11884
rect 1232 -11904 1242 -11894
rect 982 -11954 1242 -11904
rect 1302 -11954 1312 -11894
rect 912 -11964 1312 -11954
rect 1370 -11544 1770 -11534
rect 1370 -11604 1380 -11544
rect 1440 -11594 1700 -11544
rect 1440 -11604 1450 -11594
rect 1370 -11614 1450 -11604
rect 1690 -11604 1700 -11594
rect 1760 -11604 1770 -11544
rect 1690 -11614 1770 -11604
rect 1370 -11884 1430 -11614
rect 1700 -11624 1770 -11614
rect 1510 -11674 1540 -11654
rect 1490 -11714 1540 -11674
rect 1600 -11674 1630 -11654
rect 1600 -11714 1650 -11674
rect 1490 -11784 1650 -11714
rect 1490 -11824 1540 -11784
rect 1510 -11844 1540 -11824
rect 1600 -11824 1650 -11784
rect 1600 -11844 1630 -11824
rect 1710 -11884 1770 -11624
rect 1370 -11894 1450 -11884
rect 1370 -11954 1380 -11894
rect 1440 -11904 1450 -11894
rect 1690 -11894 1770 -11884
rect 1690 -11904 1700 -11894
rect 1440 -11954 1700 -11904
rect 1760 -11954 1770 -11894
rect 1370 -11964 1770 -11954
rect 1826 -11544 2226 -11534
rect 1826 -11604 1836 -11544
rect 1896 -11594 2156 -11544
rect 1896 -11604 1906 -11594
rect 1826 -11614 1906 -11604
rect 2146 -11604 2156 -11594
rect 2216 -11604 2226 -11544
rect 2146 -11614 2226 -11604
rect 1826 -11884 1886 -11614
rect 2156 -11624 2226 -11614
rect 1966 -11674 1996 -11654
rect 1946 -11714 1996 -11674
rect 2056 -11674 2086 -11654
rect 2056 -11714 2106 -11674
rect 1946 -11784 2106 -11714
rect 1946 -11824 1996 -11784
rect 1966 -11844 1996 -11824
rect 2056 -11824 2106 -11784
rect 2056 -11844 2086 -11824
rect 2166 -11884 2226 -11624
rect 1826 -11894 1906 -11884
rect 1826 -11954 1836 -11894
rect 1896 -11904 1906 -11894
rect 2146 -11894 2226 -11884
rect 2146 -11904 2156 -11894
rect 1896 -11954 2156 -11904
rect 2216 -11954 2226 -11894
rect 1826 -11964 2226 -11954
rect 2282 -11544 2682 -11534
rect 2282 -11604 2292 -11544
rect 2352 -11594 2612 -11544
rect 2352 -11604 2362 -11594
rect 2282 -11614 2362 -11604
rect 2602 -11604 2612 -11594
rect 2672 -11604 2682 -11544
rect 2602 -11614 2682 -11604
rect 2282 -11884 2342 -11614
rect 2612 -11624 2682 -11614
rect 2422 -11674 2452 -11654
rect 2402 -11714 2452 -11674
rect 2512 -11674 2542 -11654
rect 2512 -11714 2562 -11674
rect 2402 -11784 2562 -11714
rect 2402 -11824 2452 -11784
rect 2422 -11844 2452 -11824
rect 2512 -11824 2562 -11784
rect 2512 -11844 2542 -11824
rect 2622 -11884 2682 -11624
rect 2282 -11894 2362 -11884
rect 2282 -11954 2292 -11894
rect 2352 -11904 2362 -11894
rect 2602 -11894 2682 -11884
rect 2602 -11904 2612 -11894
rect 2352 -11954 2612 -11904
rect 2672 -11954 2682 -11894
rect 2282 -11964 2682 -11954
rect 2740 -11544 3140 -11534
rect 2740 -11604 2750 -11544
rect 2810 -11594 3070 -11544
rect 2810 -11604 2820 -11594
rect 2740 -11614 2820 -11604
rect 3060 -11604 3070 -11594
rect 3130 -11604 3140 -11544
rect 3060 -11614 3140 -11604
rect 2740 -11884 2800 -11614
rect 3070 -11624 3140 -11614
rect 2880 -11674 2910 -11654
rect 2860 -11714 2910 -11674
rect 2970 -11674 3000 -11654
rect 2970 -11714 3020 -11674
rect 2860 -11784 3020 -11714
rect 2860 -11824 2910 -11784
rect 2880 -11844 2910 -11824
rect 2970 -11824 3020 -11784
rect 2970 -11844 3000 -11824
rect 3080 -11884 3140 -11624
rect 2740 -11894 2820 -11884
rect 2740 -11954 2750 -11894
rect 2810 -11904 2820 -11894
rect 3060 -11894 3140 -11884
rect 3060 -11904 3070 -11894
rect 2810 -11954 3070 -11904
rect 3130 -11954 3140 -11894
rect 2740 -11964 3140 -11954
rect 3196 -11544 3596 -11534
rect 3196 -11604 3206 -11544
rect 3266 -11594 3526 -11544
rect 3266 -11604 3276 -11594
rect 3196 -11614 3276 -11604
rect 3516 -11604 3526 -11594
rect 3586 -11604 3596 -11544
rect 3516 -11614 3596 -11604
rect 3196 -11884 3256 -11614
rect 3526 -11624 3596 -11614
rect 3336 -11674 3366 -11654
rect 3316 -11714 3366 -11674
rect 3426 -11674 3456 -11654
rect 3426 -11714 3476 -11674
rect 3316 -11784 3476 -11714
rect 3316 -11824 3366 -11784
rect 3336 -11844 3366 -11824
rect 3426 -11824 3476 -11784
rect 3426 -11844 3456 -11824
rect 3536 -11884 3596 -11624
rect 3196 -11894 3276 -11884
rect 3196 -11954 3206 -11894
rect 3266 -11904 3276 -11894
rect 3516 -11894 3596 -11884
rect 3516 -11904 3526 -11894
rect 3266 -11954 3526 -11904
rect 3586 -11954 3596 -11894
rect 3196 -11964 3596 -11954
rect 3652 -11544 4052 -11534
rect 3652 -11604 3662 -11544
rect 3722 -11594 3982 -11544
rect 3722 -11604 3732 -11594
rect 3652 -11614 3732 -11604
rect 3972 -11604 3982 -11594
rect 4042 -11604 4052 -11544
rect 3972 -11614 4052 -11604
rect 3652 -11884 3712 -11614
rect 3982 -11624 4052 -11614
rect 3792 -11674 3822 -11654
rect 3772 -11714 3822 -11674
rect 3882 -11674 3912 -11654
rect 3882 -11714 3932 -11674
rect 3772 -11784 3932 -11714
rect 3772 -11824 3822 -11784
rect 3792 -11844 3822 -11824
rect 3882 -11824 3932 -11784
rect 3882 -11844 3912 -11824
rect 3992 -11884 4052 -11624
rect 3652 -11894 3732 -11884
rect 3652 -11954 3662 -11894
rect 3722 -11904 3732 -11894
rect 3972 -11894 4052 -11884
rect 3972 -11904 3982 -11894
rect 3722 -11954 3982 -11904
rect 4042 -11954 4052 -11894
rect 3652 -11964 4052 -11954
rect 4110 -11544 4510 -11534
rect 4110 -11604 4120 -11544
rect 4180 -11594 4440 -11544
rect 4180 -11604 4190 -11594
rect 4110 -11614 4190 -11604
rect 4430 -11604 4440 -11594
rect 4500 -11604 4510 -11544
rect 4430 -11614 4510 -11604
rect 4110 -11884 4170 -11614
rect 4440 -11624 4510 -11614
rect 4250 -11674 4280 -11654
rect 4230 -11714 4280 -11674
rect 4340 -11674 4370 -11654
rect 4340 -11714 4390 -11674
rect 4230 -11784 4390 -11714
rect 4230 -11824 4280 -11784
rect 4250 -11844 4280 -11824
rect 4340 -11824 4390 -11784
rect 4340 -11844 4370 -11824
rect 4450 -11884 4510 -11624
rect 4110 -11894 4190 -11884
rect 4110 -11954 4120 -11894
rect 4180 -11904 4190 -11894
rect 4430 -11894 4510 -11884
rect 4430 -11904 4440 -11894
rect 4180 -11954 4440 -11904
rect 4500 -11954 4510 -11894
rect 4110 -11964 4510 -11954
rect 4566 -11544 4966 -11534
rect 4566 -11604 4576 -11544
rect 4636 -11594 4896 -11544
rect 4636 -11604 4646 -11594
rect 4566 -11614 4646 -11604
rect 4886 -11604 4896 -11594
rect 4956 -11604 4966 -11544
rect 4886 -11614 4966 -11604
rect 4566 -11884 4626 -11614
rect 4896 -11624 4966 -11614
rect 4706 -11674 4736 -11654
rect 4686 -11714 4736 -11674
rect 4796 -11674 4826 -11654
rect 4796 -11714 4846 -11674
rect 4686 -11784 4846 -11714
rect 4686 -11824 4736 -11784
rect 4706 -11844 4736 -11824
rect 4796 -11824 4846 -11784
rect 4796 -11844 4826 -11824
rect 4906 -11884 4966 -11624
rect 4566 -11894 4646 -11884
rect 4566 -11954 4576 -11894
rect 4636 -11904 4646 -11894
rect 4886 -11894 4966 -11884
rect 4886 -11904 4896 -11894
rect 4636 -11954 4896 -11904
rect 4956 -11954 4966 -11894
rect 4566 -11964 4966 -11954
rect 5022 -11544 5422 -11534
rect 5022 -11604 5032 -11544
rect 5092 -11594 5352 -11544
rect 5092 -11604 5102 -11594
rect 5022 -11614 5102 -11604
rect 5342 -11604 5352 -11594
rect 5412 -11604 5422 -11544
rect 5342 -11614 5422 -11604
rect 5022 -11884 5082 -11614
rect 5352 -11624 5422 -11614
rect 5162 -11674 5192 -11654
rect 5142 -11714 5192 -11674
rect 5252 -11674 5282 -11654
rect 5252 -11714 5302 -11674
rect 5142 -11784 5302 -11714
rect 5142 -11824 5192 -11784
rect 5162 -11844 5192 -11824
rect 5252 -11824 5302 -11784
rect 5252 -11844 5282 -11824
rect 5362 -11884 5422 -11624
rect 5022 -11894 5102 -11884
rect 5022 -11954 5032 -11894
rect 5092 -11904 5102 -11894
rect 5342 -11894 5422 -11884
rect 5342 -11904 5352 -11894
rect 5092 -11954 5352 -11904
rect 5412 -11954 5422 -11894
rect 5022 -11964 5422 -11954
rect 5480 -11544 5880 -11534
rect 5480 -11604 5490 -11544
rect 5550 -11594 5810 -11544
rect 5550 -11604 5560 -11594
rect 5480 -11614 5560 -11604
rect 5800 -11604 5810 -11594
rect 5870 -11604 5880 -11544
rect 5800 -11614 5880 -11604
rect 5480 -11884 5540 -11614
rect 5810 -11624 5880 -11614
rect 5620 -11674 5650 -11654
rect 5600 -11714 5650 -11674
rect 5710 -11674 5740 -11654
rect 5710 -11714 5760 -11674
rect 5600 -11784 5760 -11714
rect 5600 -11824 5650 -11784
rect 5620 -11844 5650 -11824
rect 5710 -11824 5760 -11784
rect 5710 -11844 5740 -11824
rect 5820 -11884 5880 -11624
rect 5480 -11894 5560 -11884
rect 5480 -11954 5490 -11894
rect 5550 -11904 5560 -11894
rect 5800 -11894 5880 -11884
rect 5800 -11904 5810 -11894
rect 5550 -11954 5810 -11904
rect 5870 -11954 5880 -11894
rect 5480 -11964 5880 -11954
rect 5936 -11544 6336 -11534
rect 5936 -11604 5946 -11544
rect 6006 -11594 6266 -11544
rect 6006 -11604 6016 -11594
rect 5936 -11614 6016 -11604
rect 6256 -11604 6266 -11594
rect 6326 -11604 6336 -11544
rect 6256 -11614 6336 -11604
rect 5936 -11884 5996 -11614
rect 6266 -11624 6336 -11614
rect 6076 -11674 6106 -11654
rect 6056 -11714 6106 -11674
rect 6166 -11674 6196 -11654
rect 6166 -11714 6216 -11674
rect 6056 -11784 6216 -11714
rect 6056 -11824 6106 -11784
rect 6076 -11844 6106 -11824
rect 6166 -11824 6216 -11784
rect 6166 -11844 6196 -11824
rect 6276 -11884 6336 -11624
rect 5936 -11894 6016 -11884
rect 5936 -11954 5946 -11894
rect 6006 -11904 6016 -11894
rect 6256 -11894 6336 -11884
rect 6256 -11904 6266 -11894
rect 6006 -11954 6266 -11904
rect 6326 -11954 6336 -11894
rect 5936 -11964 6336 -11954
rect 6392 -11544 6792 -11534
rect 6392 -11604 6402 -11544
rect 6462 -11594 6722 -11544
rect 6462 -11604 6472 -11594
rect 6392 -11614 6472 -11604
rect 6712 -11604 6722 -11594
rect 6782 -11604 6792 -11544
rect 6712 -11614 6792 -11604
rect 6392 -11884 6452 -11614
rect 6722 -11624 6792 -11614
rect 6532 -11674 6562 -11654
rect 6512 -11714 6562 -11674
rect 6622 -11674 6652 -11654
rect 6622 -11714 6672 -11674
rect 6512 -11784 6672 -11714
rect 6512 -11824 6562 -11784
rect 6532 -11844 6562 -11824
rect 6622 -11824 6672 -11784
rect 6622 -11844 6652 -11824
rect 6732 -11884 6792 -11624
rect 6392 -11894 6472 -11884
rect 6392 -11954 6402 -11894
rect 6462 -11904 6472 -11894
rect 6712 -11894 6792 -11884
rect 6712 -11904 6722 -11894
rect 6462 -11954 6722 -11904
rect 6782 -11954 6792 -11894
rect 6392 -11964 6792 -11954
rect 6850 -11544 7250 -11534
rect 6850 -11604 6860 -11544
rect 6920 -11594 7180 -11544
rect 6920 -11604 6930 -11594
rect 6850 -11614 6930 -11604
rect 7170 -11604 7180 -11594
rect 7240 -11604 7250 -11544
rect 7170 -11614 7250 -11604
rect 6850 -11884 6910 -11614
rect 7180 -11624 7250 -11614
rect 6990 -11674 7020 -11654
rect 6970 -11714 7020 -11674
rect 7080 -11674 7110 -11654
rect 7080 -11714 7130 -11674
rect 6970 -11784 7130 -11714
rect 6970 -11824 7020 -11784
rect 6990 -11844 7020 -11824
rect 7080 -11824 7130 -11784
rect 7080 -11844 7110 -11824
rect 7190 -11884 7250 -11624
rect 6850 -11894 6930 -11884
rect 6850 -11954 6860 -11894
rect 6920 -11904 6930 -11894
rect 7170 -11894 7250 -11884
rect 7170 -11904 7180 -11894
rect 6920 -11954 7180 -11904
rect 7240 -11954 7250 -11894
rect 6850 -11964 7250 -11954
rect 7306 -11544 7706 -11534
rect 7306 -11604 7316 -11544
rect 7376 -11594 7636 -11544
rect 7376 -11604 7386 -11594
rect 7306 -11614 7386 -11604
rect 7626 -11604 7636 -11594
rect 7696 -11604 7706 -11544
rect 7626 -11614 7706 -11604
rect 7306 -11884 7366 -11614
rect 7636 -11624 7706 -11614
rect 7446 -11674 7476 -11654
rect 7426 -11714 7476 -11674
rect 7536 -11674 7566 -11654
rect 7536 -11714 7586 -11674
rect 7426 -11784 7586 -11714
rect 7426 -11824 7476 -11784
rect 7446 -11844 7476 -11824
rect 7536 -11824 7586 -11784
rect 7536 -11844 7566 -11824
rect 7646 -11884 7706 -11624
rect 7306 -11894 7386 -11884
rect 7306 -11954 7316 -11894
rect 7376 -11904 7386 -11894
rect 7626 -11894 7706 -11884
rect 7626 -11904 7636 -11894
rect 7376 -11954 7636 -11904
rect 7696 -11954 7706 -11894
rect 7306 -11964 7706 -11954
rect 7762 -11544 8162 -11534
rect 7762 -11604 7772 -11544
rect 7832 -11594 8092 -11544
rect 7832 -11604 7842 -11594
rect 7762 -11614 7842 -11604
rect 8082 -11604 8092 -11594
rect 8152 -11604 8162 -11544
rect 8082 -11614 8162 -11604
rect 7762 -11884 7822 -11614
rect 8092 -11624 8162 -11614
rect 7902 -11674 7932 -11654
rect 7882 -11714 7932 -11674
rect 7992 -11674 8022 -11654
rect 7992 -11714 8042 -11674
rect 7882 -11784 8042 -11714
rect 7882 -11824 7932 -11784
rect 7902 -11844 7932 -11824
rect 7992 -11824 8042 -11784
rect 7992 -11844 8022 -11824
rect 8102 -11884 8162 -11624
rect 7762 -11894 7842 -11884
rect 7762 -11954 7772 -11894
rect 7832 -11904 7842 -11894
rect 8082 -11894 8162 -11884
rect 8082 -11904 8092 -11894
rect 7832 -11954 8092 -11904
rect 8152 -11954 8162 -11894
rect 7762 -11964 8162 -11954
rect 8236 -11544 8636 -11534
rect 8236 -11604 8246 -11544
rect 8306 -11594 8566 -11544
rect 8306 -11604 8316 -11594
rect 8236 -11614 8316 -11604
rect 8556 -11604 8566 -11594
rect 8626 -11604 8636 -11544
rect 8556 -11614 8636 -11604
rect 8236 -11884 8296 -11614
rect 8566 -11624 8636 -11614
rect 8376 -11674 8406 -11654
rect 8356 -11714 8406 -11674
rect 8466 -11674 8496 -11654
rect 8466 -11714 8516 -11674
rect 8356 -11784 8516 -11714
rect 8356 -11824 8406 -11784
rect 8376 -11844 8406 -11824
rect 8466 -11824 8516 -11784
rect 8466 -11844 8496 -11824
rect 8576 -11884 8636 -11624
rect 8236 -11894 8316 -11884
rect 8236 -11954 8246 -11894
rect 8306 -11904 8316 -11894
rect 8556 -11894 8636 -11884
rect 8556 -11904 8566 -11894
rect 8306 -11954 8566 -11904
rect 8626 -11954 8636 -11894
rect 8236 -11964 8636 -11954
rect 8692 -11544 9092 -11534
rect 8692 -11604 8702 -11544
rect 8762 -11594 9022 -11544
rect 8762 -11604 8772 -11594
rect 8692 -11614 8772 -11604
rect 9012 -11604 9022 -11594
rect 9082 -11604 9092 -11544
rect 9012 -11614 9092 -11604
rect 8692 -11884 8752 -11614
rect 9022 -11624 9092 -11614
rect 8832 -11674 8862 -11654
rect 8812 -11714 8862 -11674
rect 8922 -11674 8952 -11654
rect 8922 -11714 8972 -11674
rect 8812 -11784 8972 -11714
rect 8812 -11824 8862 -11784
rect 8832 -11844 8862 -11824
rect 8922 -11824 8972 -11784
rect 8922 -11844 8952 -11824
rect 9032 -11884 9092 -11624
rect 8692 -11894 8772 -11884
rect 8692 -11954 8702 -11894
rect 8762 -11904 8772 -11894
rect 9012 -11894 9092 -11884
rect 9012 -11904 9022 -11894
rect 8762 -11954 9022 -11904
rect 9082 -11954 9092 -11894
rect 8692 -11964 9092 -11954
rect 9150 -11544 9550 -11534
rect 9150 -11604 9160 -11544
rect 9220 -11594 9480 -11544
rect 9220 -11604 9230 -11594
rect 9150 -11614 9230 -11604
rect 9470 -11604 9480 -11594
rect 9540 -11604 9550 -11544
rect 9470 -11614 9550 -11604
rect 9150 -11884 9210 -11614
rect 9480 -11624 9550 -11614
rect 9290 -11674 9320 -11654
rect 9270 -11714 9320 -11674
rect 9380 -11674 9410 -11654
rect 9380 -11714 9430 -11674
rect 9270 -11784 9430 -11714
rect 9270 -11824 9320 -11784
rect 9290 -11844 9320 -11824
rect 9380 -11824 9430 -11784
rect 9380 -11844 9410 -11824
rect 9490 -11884 9550 -11624
rect 9607 -11544 10006 -11534
rect 9607 -11604 9616 -11544
rect 9676 -11594 9936 -11544
rect 9676 -11604 9686 -11594
rect 9607 -11614 9686 -11604
rect 9926 -11604 9936 -11594
rect 9996 -11604 10006 -11544
rect 9926 -11614 10006 -11604
rect 9607 -11787 9666 -11614
rect 9936 -11624 10006 -11614
rect 9746 -11674 9776 -11654
rect 9150 -11894 9230 -11884
rect 9150 -11954 9160 -11894
rect 9220 -11904 9230 -11894
rect 9470 -11894 9550 -11884
rect 9470 -11904 9480 -11894
rect 9220 -11954 9480 -11904
rect 9540 -11954 9550 -11894
rect 9150 -11964 9550 -11954
rect 9606 -11884 9666 -11787
rect 9726 -11714 9776 -11674
rect 9836 -11674 9866 -11654
rect 9836 -11714 9886 -11674
rect 9726 -11784 9886 -11714
rect 9726 -11824 9776 -11784
rect 9746 -11844 9776 -11824
rect 9836 -11824 9886 -11784
rect 9836 -11844 9866 -11824
rect 9946 -11884 10006 -11624
rect 9606 -11894 9686 -11884
rect 9606 -11954 9616 -11894
rect 9676 -11904 9686 -11894
rect 9926 -11894 10006 -11884
rect 9926 -11904 9936 -11894
rect 9676 -11954 9936 -11904
rect 9996 -11954 10006 -11894
rect 9606 -11964 10006 -11954
rect 10062 -11544 10462 -11534
rect 10062 -11604 10072 -11544
rect 10132 -11594 10392 -11544
rect 10132 -11604 10142 -11594
rect 10062 -11614 10142 -11604
rect 10382 -11604 10392 -11594
rect 10452 -11604 10462 -11544
rect 10382 -11614 10462 -11604
rect 10062 -11884 10122 -11614
rect 10392 -11624 10462 -11614
rect 10202 -11674 10232 -11654
rect 10182 -11714 10232 -11674
rect 10292 -11674 10322 -11654
rect 10292 -11714 10342 -11674
rect 10182 -11784 10342 -11714
rect 10182 -11824 10232 -11784
rect 10202 -11844 10232 -11824
rect 10292 -11824 10342 -11784
rect 10292 -11844 10322 -11824
rect 10402 -11884 10462 -11624
rect 10062 -11894 10142 -11884
rect 10062 -11954 10072 -11894
rect 10132 -11904 10142 -11894
rect 10382 -11894 10462 -11884
rect 10382 -11904 10392 -11894
rect 10132 -11954 10392 -11904
rect 10452 -11954 10462 -11894
rect 10062 -11964 10462 -11954
rect 10520 -11544 10920 -11534
rect 10520 -11604 10530 -11544
rect 10590 -11594 10850 -11544
rect 10590 -11604 10600 -11594
rect 10520 -11614 10600 -11604
rect 10840 -11604 10850 -11594
rect 10910 -11604 10920 -11544
rect 10840 -11614 10920 -11604
rect 10520 -11884 10580 -11614
rect 10850 -11624 10920 -11614
rect 10660 -11674 10690 -11654
rect 10640 -11714 10690 -11674
rect 10750 -11674 10780 -11654
rect 10750 -11714 10800 -11674
rect 10640 -11784 10800 -11714
rect 10640 -11824 10690 -11784
rect 10660 -11844 10690 -11824
rect 10750 -11824 10800 -11784
rect 10750 -11844 10780 -11824
rect 10860 -11884 10920 -11624
rect 10520 -11894 10600 -11884
rect 10520 -11954 10530 -11894
rect 10590 -11904 10600 -11894
rect 10840 -11894 10920 -11884
rect 10840 -11904 10850 -11894
rect 10590 -11954 10850 -11904
rect 10910 -11954 10920 -11894
rect 10520 -11964 10920 -11954
rect 10976 -11544 11376 -11534
rect 10976 -11604 10986 -11544
rect 11046 -11594 11306 -11544
rect 11046 -11604 11056 -11594
rect 10976 -11614 11056 -11604
rect 11296 -11604 11306 -11594
rect 11366 -11604 11376 -11544
rect 11296 -11614 11376 -11604
rect 10976 -11884 11036 -11614
rect 11306 -11624 11376 -11614
rect 11116 -11674 11146 -11654
rect 11096 -11714 11146 -11674
rect 11206 -11674 11236 -11654
rect 11206 -11714 11256 -11674
rect 11096 -11784 11256 -11714
rect 11096 -11824 11146 -11784
rect 11116 -11844 11146 -11824
rect 11206 -11824 11256 -11784
rect 11206 -11844 11236 -11824
rect 11316 -11884 11376 -11624
rect 10976 -11894 11056 -11884
rect 10976 -11954 10986 -11894
rect 11046 -11904 11056 -11894
rect 11296 -11894 11376 -11884
rect 11296 -11904 11306 -11894
rect 11046 -11954 11306 -11904
rect 11366 -11954 11376 -11894
rect 10976 -11964 11376 -11954
rect 11432 -11544 11832 -11534
rect 11432 -11604 11442 -11544
rect 11502 -11594 11762 -11544
rect 11502 -11604 11512 -11594
rect 11432 -11614 11512 -11604
rect 11752 -11604 11762 -11594
rect 11822 -11604 11832 -11544
rect 11752 -11614 11832 -11604
rect 11432 -11884 11492 -11614
rect 11762 -11624 11832 -11614
rect 11572 -11674 11602 -11654
rect 11552 -11714 11602 -11674
rect 11662 -11674 11692 -11654
rect 11662 -11714 11712 -11674
rect 11552 -11784 11712 -11714
rect 11552 -11824 11602 -11784
rect 11572 -11844 11602 -11824
rect 11662 -11824 11712 -11784
rect 11662 -11844 11692 -11824
rect 11772 -11884 11832 -11624
rect 11432 -11894 11512 -11884
rect 11432 -11954 11442 -11894
rect 11502 -11904 11512 -11894
rect 11752 -11894 11832 -11884
rect 11752 -11904 11762 -11894
rect 11502 -11954 11762 -11904
rect 11822 -11954 11832 -11894
rect 11432 -11964 11832 -11954
rect 11890 -11544 12290 -11534
rect 11890 -11604 11900 -11544
rect 11960 -11594 12220 -11544
rect 11960 -11604 11970 -11594
rect 11890 -11614 11970 -11604
rect 12210 -11604 12220 -11594
rect 12280 -11604 12290 -11544
rect 12210 -11614 12290 -11604
rect 11890 -11884 11950 -11614
rect 12220 -11624 12290 -11614
rect 12030 -11674 12060 -11654
rect 12010 -11714 12060 -11674
rect 12120 -11674 12150 -11654
rect 12120 -11714 12170 -11674
rect 12010 -11784 12170 -11714
rect 12010 -11824 12060 -11784
rect 12030 -11844 12060 -11824
rect 12120 -11824 12170 -11784
rect 12120 -11844 12150 -11824
rect 12230 -11884 12290 -11624
rect 11890 -11894 11970 -11884
rect 11890 -11954 11900 -11894
rect 11960 -11904 11970 -11894
rect 12210 -11894 12290 -11884
rect 12210 -11904 12220 -11894
rect 11960 -11954 12220 -11904
rect 12280 -11954 12290 -11894
rect 11890 -11964 12290 -11954
rect 12346 -11544 12746 -11534
rect 12346 -11604 12356 -11544
rect 12416 -11594 12676 -11544
rect 12416 -11604 12426 -11594
rect 12346 -11614 12426 -11604
rect 12666 -11604 12676 -11594
rect 12736 -11604 12746 -11544
rect 12666 -11614 12746 -11604
rect 12346 -11884 12406 -11614
rect 12676 -11624 12746 -11614
rect 12486 -11674 12516 -11654
rect 12466 -11714 12516 -11674
rect 12576 -11674 12606 -11654
rect 12576 -11714 12626 -11674
rect 12466 -11784 12626 -11714
rect 12466 -11824 12516 -11784
rect 12486 -11844 12516 -11824
rect 12576 -11824 12626 -11784
rect 12576 -11844 12606 -11824
rect 12686 -11884 12746 -11624
rect 12346 -11894 12426 -11884
rect 12346 -11954 12356 -11894
rect 12416 -11904 12426 -11894
rect 12666 -11894 12746 -11884
rect 12666 -11904 12676 -11894
rect 12416 -11954 12676 -11904
rect 12736 -11954 12746 -11894
rect 12346 -11964 12746 -11954
rect 12802 -11544 13202 -11534
rect 12802 -11604 12812 -11544
rect 12872 -11594 13132 -11544
rect 12872 -11604 12882 -11594
rect 12802 -11614 12882 -11604
rect 13122 -11604 13132 -11594
rect 13192 -11604 13202 -11544
rect 13122 -11614 13202 -11604
rect 12802 -11884 12862 -11614
rect 13132 -11624 13202 -11614
rect 12942 -11674 12972 -11654
rect 12922 -11714 12972 -11674
rect 13032 -11674 13062 -11654
rect 13032 -11714 13082 -11674
rect 12922 -11784 13082 -11714
rect 12922 -11824 12972 -11784
rect 12942 -11844 12972 -11824
rect 13032 -11824 13082 -11784
rect 13032 -11844 13062 -11824
rect 13142 -11884 13202 -11624
rect 12802 -11894 12882 -11884
rect 12802 -11954 12812 -11894
rect 12872 -11904 12882 -11894
rect 13122 -11894 13202 -11884
rect 13122 -11904 13132 -11894
rect 12872 -11954 13132 -11904
rect 13192 -11954 13202 -11894
rect 12802 -11964 13202 -11954
rect 13260 -11544 13660 -11534
rect 13260 -11604 13270 -11544
rect 13330 -11594 13590 -11544
rect 13330 -11604 13340 -11594
rect 13260 -11614 13340 -11604
rect 13580 -11604 13590 -11594
rect 13650 -11604 13660 -11544
rect 13580 -11614 13660 -11604
rect 13260 -11884 13320 -11614
rect 13590 -11624 13660 -11614
rect 13400 -11674 13430 -11654
rect 13380 -11714 13430 -11674
rect 13490 -11674 13520 -11654
rect 13490 -11714 13540 -11674
rect 13380 -11784 13540 -11714
rect 13380 -11824 13430 -11784
rect 13400 -11844 13430 -11824
rect 13490 -11824 13540 -11784
rect 13490 -11844 13520 -11824
rect 13600 -11884 13660 -11624
rect 13260 -11894 13340 -11884
rect 13260 -11954 13270 -11894
rect 13330 -11904 13340 -11894
rect 13580 -11894 13660 -11884
rect 13580 -11904 13590 -11894
rect 13330 -11954 13590 -11904
rect 13650 -11954 13660 -11894
rect 13260 -11964 13660 -11954
rect 13716 -11544 14116 -11534
rect 13716 -11604 13726 -11544
rect 13786 -11594 14046 -11544
rect 13786 -11604 13796 -11594
rect 13716 -11614 13796 -11604
rect 14036 -11604 14046 -11594
rect 14106 -11604 14116 -11544
rect 14036 -11614 14116 -11604
rect 13716 -11884 13776 -11614
rect 14046 -11624 14116 -11614
rect 13856 -11674 13886 -11654
rect 13836 -11714 13886 -11674
rect 13946 -11674 13976 -11654
rect 13946 -11714 13996 -11674
rect 13836 -11784 13996 -11714
rect 13836 -11824 13886 -11784
rect 13856 -11844 13886 -11824
rect 13946 -11824 13996 -11784
rect 13946 -11844 13976 -11824
rect 14056 -11884 14116 -11624
rect 13716 -11894 13796 -11884
rect 13716 -11954 13726 -11894
rect 13786 -11904 13796 -11894
rect 14036 -11894 14116 -11884
rect 14036 -11904 14046 -11894
rect 13786 -11954 14046 -11904
rect 14106 -11954 14116 -11894
rect 13716 -11964 14116 -11954
rect 14172 -11544 14572 -11534
rect 14172 -11604 14182 -11544
rect 14242 -11594 14502 -11544
rect 14242 -11604 14252 -11594
rect 14172 -11614 14252 -11604
rect 14492 -11604 14502 -11594
rect 14562 -11604 14572 -11544
rect 14492 -11614 14572 -11604
rect 14172 -11884 14232 -11614
rect 14502 -11624 14572 -11614
rect 14312 -11674 14342 -11654
rect 14292 -11714 14342 -11674
rect 14402 -11674 14432 -11654
rect 14402 -11714 14452 -11674
rect 14292 -11784 14452 -11714
rect 14292 -11824 14342 -11784
rect 14312 -11844 14342 -11824
rect 14402 -11824 14452 -11784
rect 14402 -11844 14432 -11824
rect 14512 -11884 14572 -11624
rect 14172 -11894 14252 -11884
rect 14172 -11954 14182 -11894
rect 14242 -11904 14252 -11894
rect 14492 -11894 14572 -11884
rect 14492 -11904 14502 -11894
rect 14242 -11954 14502 -11904
rect 14562 -11954 14572 -11894
rect 14172 -11964 14572 -11954
rect 14630 -11544 15030 -11534
rect 14630 -11604 14640 -11544
rect 14700 -11594 14960 -11544
rect 14700 -11604 14710 -11594
rect 14630 -11614 14710 -11604
rect 14950 -11604 14960 -11594
rect 15020 -11604 15030 -11544
rect 14950 -11614 15030 -11604
rect 14630 -11884 14690 -11614
rect 14960 -11624 15030 -11614
rect 14770 -11674 14800 -11654
rect 14750 -11714 14800 -11674
rect 14860 -11674 14890 -11654
rect 14860 -11714 14910 -11674
rect 14750 -11784 14910 -11714
rect 14750 -11824 14800 -11784
rect 14770 -11844 14800 -11824
rect 14860 -11824 14910 -11784
rect 14860 -11844 14890 -11824
rect 14970 -11884 15030 -11624
rect 14630 -11894 14710 -11884
rect 14630 -11954 14640 -11894
rect 14700 -11904 14710 -11894
rect 14950 -11894 15030 -11884
rect 14950 -11904 14960 -11894
rect 14700 -11954 14960 -11904
rect 15020 -11954 15030 -11894
rect 14630 -11964 15030 -11954
rect 15086 -11544 15486 -11534
rect 15086 -11604 15096 -11544
rect 15156 -11594 15416 -11544
rect 15156 -11604 15166 -11594
rect 15086 -11614 15166 -11604
rect 15406 -11604 15416 -11594
rect 15476 -11604 15486 -11544
rect 15406 -11614 15486 -11604
rect 15086 -11884 15146 -11614
rect 15416 -11624 15486 -11614
rect 15226 -11674 15256 -11654
rect 15206 -11714 15256 -11674
rect 15316 -11674 15346 -11654
rect 15316 -11714 15366 -11674
rect 15206 -11784 15366 -11714
rect 15206 -11824 15256 -11784
rect 15226 -11844 15256 -11824
rect 15316 -11824 15366 -11784
rect 15316 -11844 15346 -11824
rect 15426 -11884 15486 -11624
rect 15086 -11894 15166 -11884
rect 15086 -11954 15096 -11894
rect 15156 -11904 15166 -11894
rect 15406 -11894 15486 -11884
rect 15406 -11904 15416 -11894
rect 15156 -11954 15416 -11904
rect 15476 -11954 15486 -11894
rect 15086 -11964 15486 -11954
rect 0 -12036 400 -12026
rect 0 -12096 10 -12036
rect 70 -12086 330 -12036
rect 70 -12096 80 -12086
rect 0 -12106 80 -12096
rect 320 -12096 330 -12086
rect 390 -12096 400 -12036
rect 320 -12106 400 -12096
rect 0 -12376 60 -12106
rect 330 -12116 400 -12106
rect 140 -12166 170 -12146
rect 120 -12206 170 -12166
rect 230 -12166 260 -12146
rect 230 -12206 280 -12166
rect 120 -12276 280 -12206
rect 120 -12316 170 -12276
rect 140 -12336 170 -12316
rect 230 -12316 280 -12276
rect 230 -12336 260 -12316
rect 340 -12376 400 -12116
rect 0 -12386 80 -12376
rect 0 -12446 10 -12386
rect 70 -12396 80 -12386
rect 320 -12386 400 -12376
rect 320 -12396 330 -12386
rect 70 -12446 330 -12396
rect 390 -12446 400 -12386
rect 0 -12456 400 -12446
rect 456 -12036 856 -12026
rect 456 -12096 466 -12036
rect 526 -12086 786 -12036
rect 526 -12096 536 -12086
rect 456 -12106 536 -12096
rect 776 -12096 786 -12086
rect 846 -12096 856 -12036
rect 776 -12106 856 -12096
rect 456 -12376 516 -12106
rect 786 -12116 856 -12106
rect 596 -12166 626 -12146
rect 576 -12206 626 -12166
rect 686 -12166 716 -12146
rect 686 -12206 736 -12166
rect 576 -12276 736 -12206
rect 576 -12316 626 -12276
rect 596 -12336 626 -12316
rect 686 -12316 736 -12276
rect 686 -12336 716 -12316
rect 796 -12376 856 -12116
rect 456 -12386 536 -12376
rect 456 -12446 466 -12386
rect 526 -12396 536 -12386
rect 776 -12386 856 -12376
rect 776 -12396 786 -12386
rect 526 -12446 786 -12396
rect 846 -12446 856 -12386
rect 456 -12456 856 -12446
rect 912 -12036 1312 -12026
rect 912 -12096 922 -12036
rect 982 -12086 1242 -12036
rect 982 -12096 992 -12086
rect 912 -12106 992 -12096
rect 1232 -12096 1242 -12086
rect 1302 -12096 1312 -12036
rect 1232 -12106 1312 -12096
rect 912 -12376 972 -12106
rect 1242 -12116 1312 -12106
rect 1052 -12166 1082 -12146
rect 1032 -12206 1082 -12166
rect 1142 -12166 1172 -12146
rect 1142 -12206 1192 -12166
rect 1032 -12276 1192 -12206
rect 1032 -12316 1082 -12276
rect 1052 -12336 1082 -12316
rect 1142 -12316 1192 -12276
rect 1142 -12336 1172 -12316
rect 1252 -12376 1312 -12116
rect 912 -12386 992 -12376
rect 912 -12446 922 -12386
rect 982 -12396 992 -12386
rect 1232 -12386 1312 -12376
rect 1232 -12396 1242 -12386
rect 982 -12446 1242 -12396
rect 1302 -12446 1312 -12386
rect 912 -12456 1312 -12446
rect 1370 -12036 1770 -12026
rect 1370 -12096 1380 -12036
rect 1440 -12086 1700 -12036
rect 1440 -12096 1450 -12086
rect 1370 -12106 1450 -12096
rect 1690 -12096 1700 -12086
rect 1760 -12096 1770 -12036
rect 1690 -12106 1770 -12096
rect 1370 -12376 1430 -12106
rect 1700 -12116 1770 -12106
rect 1510 -12166 1540 -12146
rect 1490 -12206 1540 -12166
rect 1600 -12166 1630 -12146
rect 1600 -12206 1650 -12166
rect 1490 -12276 1650 -12206
rect 1490 -12316 1540 -12276
rect 1510 -12336 1540 -12316
rect 1600 -12316 1650 -12276
rect 1600 -12336 1630 -12316
rect 1710 -12376 1770 -12116
rect 1370 -12386 1450 -12376
rect 1370 -12446 1380 -12386
rect 1440 -12396 1450 -12386
rect 1690 -12386 1770 -12376
rect 1690 -12396 1700 -12386
rect 1440 -12446 1700 -12396
rect 1760 -12446 1770 -12386
rect 1370 -12456 1770 -12446
rect 1826 -12036 2226 -12026
rect 1826 -12096 1836 -12036
rect 1896 -12086 2156 -12036
rect 1896 -12096 1906 -12086
rect 1826 -12106 1906 -12096
rect 2146 -12096 2156 -12086
rect 2216 -12096 2226 -12036
rect 2146 -12106 2226 -12096
rect 1826 -12376 1886 -12106
rect 2156 -12116 2226 -12106
rect 1966 -12166 1996 -12146
rect 1946 -12206 1996 -12166
rect 2056 -12166 2086 -12146
rect 2056 -12206 2106 -12166
rect 1946 -12276 2106 -12206
rect 1946 -12316 1996 -12276
rect 1966 -12336 1996 -12316
rect 2056 -12316 2106 -12276
rect 2056 -12336 2086 -12316
rect 2166 -12376 2226 -12116
rect 1826 -12386 1906 -12376
rect 1826 -12446 1836 -12386
rect 1896 -12396 1906 -12386
rect 2146 -12386 2226 -12376
rect 2146 -12396 2156 -12386
rect 1896 -12446 2156 -12396
rect 2216 -12446 2226 -12386
rect 1826 -12456 2226 -12446
rect 2282 -12036 2682 -12026
rect 2282 -12096 2292 -12036
rect 2352 -12086 2612 -12036
rect 2352 -12096 2362 -12086
rect 2282 -12106 2362 -12096
rect 2602 -12096 2612 -12086
rect 2672 -12096 2682 -12036
rect 2602 -12106 2682 -12096
rect 2282 -12376 2342 -12106
rect 2612 -12116 2682 -12106
rect 2422 -12166 2452 -12146
rect 2402 -12206 2452 -12166
rect 2512 -12166 2542 -12146
rect 2512 -12206 2562 -12166
rect 2402 -12276 2562 -12206
rect 2402 -12316 2452 -12276
rect 2422 -12336 2452 -12316
rect 2512 -12316 2562 -12276
rect 2512 -12336 2542 -12316
rect 2622 -12376 2682 -12116
rect 2282 -12386 2362 -12376
rect 2282 -12446 2292 -12386
rect 2352 -12396 2362 -12386
rect 2602 -12386 2682 -12376
rect 2602 -12396 2612 -12386
rect 2352 -12446 2612 -12396
rect 2672 -12446 2682 -12386
rect 2282 -12456 2682 -12446
rect 2740 -12036 3140 -12026
rect 2740 -12096 2750 -12036
rect 2810 -12086 3070 -12036
rect 2810 -12096 2820 -12086
rect 2740 -12106 2820 -12096
rect 3060 -12096 3070 -12086
rect 3130 -12096 3140 -12036
rect 3060 -12106 3140 -12096
rect 2740 -12376 2800 -12106
rect 3070 -12116 3140 -12106
rect 2880 -12166 2910 -12146
rect 2860 -12206 2910 -12166
rect 2970 -12166 3000 -12146
rect 2970 -12206 3020 -12166
rect 2860 -12276 3020 -12206
rect 2860 -12316 2910 -12276
rect 2880 -12336 2910 -12316
rect 2970 -12316 3020 -12276
rect 2970 -12336 3000 -12316
rect 3080 -12376 3140 -12116
rect 2740 -12386 2820 -12376
rect 2740 -12446 2750 -12386
rect 2810 -12396 2820 -12386
rect 3060 -12386 3140 -12376
rect 3060 -12396 3070 -12386
rect 2810 -12446 3070 -12396
rect 3130 -12446 3140 -12386
rect 2740 -12456 3140 -12446
rect 3196 -12036 3596 -12026
rect 3196 -12096 3206 -12036
rect 3266 -12086 3526 -12036
rect 3266 -12096 3276 -12086
rect 3196 -12106 3276 -12096
rect 3516 -12096 3526 -12086
rect 3586 -12096 3596 -12036
rect 3516 -12106 3596 -12096
rect 3196 -12376 3256 -12106
rect 3526 -12116 3596 -12106
rect 3336 -12166 3366 -12146
rect 3316 -12206 3366 -12166
rect 3426 -12166 3456 -12146
rect 3426 -12206 3476 -12166
rect 3316 -12276 3476 -12206
rect 3316 -12316 3366 -12276
rect 3336 -12336 3366 -12316
rect 3426 -12316 3476 -12276
rect 3426 -12336 3456 -12316
rect 3536 -12376 3596 -12116
rect 3196 -12386 3276 -12376
rect 3196 -12446 3206 -12386
rect 3266 -12396 3276 -12386
rect 3516 -12386 3596 -12376
rect 3516 -12396 3526 -12386
rect 3266 -12446 3526 -12396
rect 3586 -12446 3596 -12386
rect 3196 -12456 3596 -12446
rect 3652 -12036 4052 -12026
rect 3652 -12096 3662 -12036
rect 3722 -12086 3982 -12036
rect 3722 -12096 3732 -12086
rect 3652 -12106 3732 -12096
rect 3972 -12096 3982 -12086
rect 4042 -12096 4052 -12036
rect 3972 -12106 4052 -12096
rect 3652 -12376 3712 -12106
rect 3982 -12116 4052 -12106
rect 3792 -12166 3822 -12146
rect 3772 -12206 3822 -12166
rect 3882 -12166 3912 -12146
rect 3882 -12206 3932 -12166
rect 3772 -12276 3932 -12206
rect 3772 -12316 3822 -12276
rect 3792 -12336 3822 -12316
rect 3882 -12316 3932 -12276
rect 3882 -12336 3912 -12316
rect 3992 -12376 4052 -12116
rect 3652 -12386 3732 -12376
rect 3652 -12446 3662 -12386
rect 3722 -12396 3732 -12386
rect 3972 -12386 4052 -12376
rect 3972 -12396 3982 -12386
rect 3722 -12446 3982 -12396
rect 4042 -12446 4052 -12386
rect 3652 -12456 4052 -12446
rect 4110 -12036 4510 -12026
rect 4110 -12096 4120 -12036
rect 4180 -12086 4440 -12036
rect 4180 -12096 4190 -12086
rect 4110 -12106 4190 -12096
rect 4430 -12096 4440 -12086
rect 4500 -12096 4510 -12036
rect 4430 -12106 4510 -12096
rect 4110 -12376 4170 -12106
rect 4440 -12116 4510 -12106
rect 4250 -12166 4280 -12146
rect 4230 -12206 4280 -12166
rect 4340 -12166 4370 -12146
rect 4340 -12206 4390 -12166
rect 4230 -12276 4390 -12206
rect 4230 -12316 4280 -12276
rect 4250 -12336 4280 -12316
rect 4340 -12316 4390 -12276
rect 4340 -12336 4370 -12316
rect 4450 -12376 4510 -12116
rect 4110 -12386 4190 -12376
rect 4110 -12446 4120 -12386
rect 4180 -12396 4190 -12386
rect 4430 -12386 4510 -12376
rect 4430 -12396 4440 -12386
rect 4180 -12446 4440 -12396
rect 4500 -12446 4510 -12386
rect 4110 -12456 4510 -12446
rect 4566 -12036 4966 -12026
rect 4566 -12096 4576 -12036
rect 4636 -12086 4896 -12036
rect 4636 -12096 4646 -12086
rect 4566 -12106 4646 -12096
rect 4886 -12096 4896 -12086
rect 4956 -12096 4966 -12036
rect 4886 -12106 4966 -12096
rect 4566 -12376 4626 -12106
rect 4896 -12116 4966 -12106
rect 4706 -12166 4736 -12146
rect 4686 -12206 4736 -12166
rect 4796 -12166 4826 -12146
rect 4796 -12206 4846 -12166
rect 4686 -12276 4846 -12206
rect 4686 -12316 4736 -12276
rect 4706 -12336 4736 -12316
rect 4796 -12316 4846 -12276
rect 4796 -12336 4826 -12316
rect 4906 -12376 4966 -12116
rect 4566 -12386 4646 -12376
rect 4566 -12446 4576 -12386
rect 4636 -12396 4646 -12386
rect 4886 -12386 4966 -12376
rect 4886 -12396 4896 -12386
rect 4636 -12446 4896 -12396
rect 4956 -12446 4966 -12386
rect 4566 -12456 4966 -12446
rect 5022 -12036 5422 -12026
rect 5022 -12096 5032 -12036
rect 5092 -12086 5352 -12036
rect 5092 -12096 5102 -12086
rect 5022 -12106 5102 -12096
rect 5342 -12096 5352 -12086
rect 5412 -12096 5422 -12036
rect 5342 -12106 5422 -12096
rect 5022 -12376 5082 -12106
rect 5352 -12116 5422 -12106
rect 5162 -12166 5192 -12146
rect 5142 -12206 5192 -12166
rect 5252 -12166 5282 -12146
rect 5252 -12206 5302 -12166
rect 5142 -12276 5302 -12206
rect 5142 -12316 5192 -12276
rect 5162 -12336 5192 -12316
rect 5252 -12316 5302 -12276
rect 5252 -12336 5282 -12316
rect 5362 -12376 5422 -12116
rect 5022 -12386 5102 -12376
rect 5022 -12446 5032 -12386
rect 5092 -12396 5102 -12386
rect 5342 -12386 5422 -12376
rect 5342 -12396 5352 -12386
rect 5092 -12446 5352 -12396
rect 5412 -12446 5422 -12386
rect 5022 -12456 5422 -12446
rect 5480 -12036 5880 -12026
rect 5480 -12096 5490 -12036
rect 5550 -12086 5810 -12036
rect 5550 -12096 5560 -12086
rect 5480 -12106 5560 -12096
rect 5800 -12096 5810 -12086
rect 5870 -12096 5880 -12036
rect 5800 -12106 5880 -12096
rect 5480 -12376 5540 -12106
rect 5810 -12116 5880 -12106
rect 5620 -12166 5650 -12146
rect 5600 -12206 5650 -12166
rect 5710 -12166 5740 -12146
rect 5710 -12206 5760 -12166
rect 5600 -12276 5760 -12206
rect 5600 -12316 5650 -12276
rect 5620 -12336 5650 -12316
rect 5710 -12316 5760 -12276
rect 5710 -12336 5740 -12316
rect 5820 -12376 5880 -12116
rect 5480 -12386 5560 -12376
rect 5480 -12446 5490 -12386
rect 5550 -12396 5560 -12386
rect 5800 -12386 5880 -12376
rect 5800 -12396 5810 -12386
rect 5550 -12446 5810 -12396
rect 5870 -12446 5880 -12386
rect 5480 -12456 5880 -12446
rect 5936 -12036 6336 -12026
rect 5936 -12096 5946 -12036
rect 6006 -12086 6266 -12036
rect 6006 -12096 6016 -12086
rect 5936 -12106 6016 -12096
rect 6256 -12096 6266 -12086
rect 6326 -12096 6336 -12036
rect 6256 -12106 6336 -12096
rect 5936 -12376 5996 -12106
rect 6266 -12116 6336 -12106
rect 6076 -12166 6106 -12146
rect 6056 -12206 6106 -12166
rect 6166 -12166 6196 -12146
rect 6166 -12206 6216 -12166
rect 6056 -12276 6216 -12206
rect 6056 -12316 6106 -12276
rect 6076 -12336 6106 -12316
rect 6166 -12316 6216 -12276
rect 6166 -12336 6196 -12316
rect 6276 -12376 6336 -12116
rect 5936 -12386 6016 -12376
rect 5936 -12446 5946 -12386
rect 6006 -12396 6016 -12386
rect 6256 -12386 6336 -12376
rect 6256 -12396 6266 -12386
rect 6006 -12446 6266 -12396
rect 6326 -12446 6336 -12386
rect 5936 -12456 6336 -12446
rect 6392 -12036 6792 -12026
rect 6392 -12096 6402 -12036
rect 6462 -12086 6722 -12036
rect 6462 -12096 6472 -12086
rect 6392 -12106 6472 -12096
rect 6712 -12096 6722 -12086
rect 6782 -12096 6792 -12036
rect 6712 -12106 6792 -12096
rect 6392 -12376 6452 -12106
rect 6722 -12116 6792 -12106
rect 6532 -12166 6562 -12146
rect 6512 -12206 6562 -12166
rect 6622 -12166 6652 -12146
rect 6622 -12206 6672 -12166
rect 6512 -12276 6672 -12206
rect 6512 -12316 6562 -12276
rect 6532 -12336 6562 -12316
rect 6622 -12316 6672 -12276
rect 6622 -12336 6652 -12316
rect 6732 -12376 6792 -12116
rect 6392 -12386 6472 -12376
rect 6392 -12446 6402 -12386
rect 6462 -12396 6472 -12386
rect 6712 -12386 6792 -12376
rect 6712 -12396 6722 -12386
rect 6462 -12446 6722 -12396
rect 6782 -12446 6792 -12386
rect 6392 -12456 6792 -12446
rect 6850 -12036 7250 -12026
rect 6850 -12096 6860 -12036
rect 6920 -12086 7180 -12036
rect 6920 -12096 6930 -12086
rect 6850 -12106 6930 -12096
rect 7170 -12096 7180 -12086
rect 7240 -12096 7250 -12036
rect 7170 -12106 7250 -12096
rect 6850 -12376 6910 -12106
rect 7180 -12116 7250 -12106
rect 6990 -12166 7020 -12146
rect 6970 -12206 7020 -12166
rect 7080 -12166 7110 -12146
rect 7080 -12206 7130 -12166
rect 6970 -12276 7130 -12206
rect 6970 -12316 7020 -12276
rect 6990 -12336 7020 -12316
rect 7080 -12316 7130 -12276
rect 7080 -12336 7110 -12316
rect 7190 -12376 7250 -12116
rect 6850 -12386 6930 -12376
rect 6850 -12446 6860 -12386
rect 6920 -12396 6930 -12386
rect 7170 -12386 7250 -12376
rect 7170 -12396 7180 -12386
rect 6920 -12446 7180 -12396
rect 7240 -12446 7250 -12386
rect 6850 -12456 7250 -12446
rect 7306 -12036 7706 -12026
rect 7306 -12096 7316 -12036
rect 7376 -12086 7636 -12036
rect 7376 -12096 7386 -12086
rect 7306 -12106 7386 -12096
rect 7626 -12096 7636 -12086
rect 7696 -12096 7706 -12036
rect 7626 -12106 7706 -12096
rect 7306 -12376 7366 -12106
rect 7636 -12116 7706 -12106
rect 7446 -12166 7476 -12146
rect 7426 -12206 7476 -12166
rect 7536 -12166 7566 -12146
rect 7536 -12206 7586 -12166
rect 7426 -12276 7586 -12206
rect 7426 -12316 7476 -12276
rect 7446 -12336 7476 -12316
rect 7536 -12316 7586 -12276
rect 7536 -12336 7566 -12316
rect 7646 -12376 7706 -12116
rect 7306 -12386 7386 -12376
rect 7306 -12446 7316 -12386
rect 7376 -12396 7386 -12386
rect 7626 -12386 7706 -12376
rect 7626 -12396 7636 -12386
rect 7376 -12446 7636 -12396
rect 7696 -12446 7706 -12386
rect 7306 -12456 7706 -12446
rect 7762 -12036 8162 -12026
rect 7762 -12096 7772 -12036
rect 7832 -12086 8092 -12036
rect 7832 -12096 7842 -12086
rect 7762 -12106 7842 -12096
rect 8082 -12096 8092 -12086
rect 8152 -12096 8162 -12036
rect 8082 -12106 8162 -12096
rect 7762 -12376 7822 -12106
rect 8092 -12116 8162 -12106
rect 7902 -12166 7932 -12146
rect 7882 -12206 7932 -12166
rect 7992 -12166 8022 -12146
rect 7992 -12206 8042 -12166
rect 7882 -12276 8042 -12206
rect 7882 -12316 7932 -12276
rect 7902 -12336 7932 -12316
rect 7992 -12316 8042 -12276
rect 7992 -12336 8022 -12316
rect 8102 -12376 8162 -12116
rect 7762 -12386 7842 -12376
rect 7762 -12446 7772 -12386
rect 7832 -12396 7842 -12386
rect 8082 -12386 8162 -12376
rect 8082 -12396 8092 -12386
rect 7832 -12446 8092 -12396
rect 8152 -12446 8162 -12386
rect 7762 -12456 8162 -12446
rect 8236 -12036 8636 -12026
rect 8236 -12096 8246 -12036
rect 8306 -12086 8566 -12036
rect 8306 -12096 8316 -12086
rect 8236 -12106 8316 -12096
rect 8556 -12096 8566 -12086
rect 8626 -12096 8636 -12036
rect 8556 -12106 8636 -12096
rect 8236 -12376 8296 -12106
rect 8566 -12116 8636 -12106
rect 8376 -12166 8406 -12146
rect 8356 -12206 8406 -12166
rect 8466 -12166 8496 -12146
rect 8466 -12206 8516 -12166
rect 8356 -12276 8516 -12206
rect 8356 -12316 8406 -12276
rect 8376 -12336 8406 -12316
rect 8466 -12316 8516 -12276
rect 8466 -12336 8496 -12316
rect 8576 -12376 8636 -12116
rect 8236 -12386 8316 -12376
rect 8236 -12446 8246 -12386
rect 8306 -12396 8316 -12386
rect 8556 -12386 8636 -12376
rect 8556 -12396 8566 -12386
rect 8306 -12446 8566 -12396
rect 8626 -12446 8636 -12386
rect 8236 -12456 8636 -12446
rect 8692 -12036 9092 -12026
rect 8692 -12096 8702 -12036
rect 8762 -12086 9022 -12036
rect 8762 -12096 8772 -12086
rect 8692 -12106 8772 -12096
rect 9012 -12096 9022 -12086
rect 9082 -12096 9092 -12036
rect 9012 -12106 9092 -12096
rect 8692 -12376 8752 -12106
rect 9022 -12116 9092 -12106
rect 8832 -12166 8862 -12146
rect 8812 -12206 8862 -12166
rect 8922 -12166 8952 -12146
rect 8922 -12206 8972 -12166
rect 8812 -12276 8972 -12206
rect 8812 -12316 8862 -12276
rect 8832 -12336 8862 -12316
rect 8922 -12316 8972 -12276
rect 8922 -12336 8952 -12316
rect 9032 -12376 9092 -12116
rect 8692 -12386 8772 -12376
rect 8692 -12446 8702 -12386
rect 8762 -12396 8772 -12386
rect 9012 -12386 9092 -12376
rect 9012 -12396 9022 -12386
rect 8762 -12446 9022 -12396
rect 9082 -12446 9092 -12386
rect 8692 -12456 9092 -12446
rect 9150 -12036 9550 -12026
rect 9150 -12096 9160 -12036
rect 9220 -12086 9480 -12036
rect 9220 -12096 9230 -12086
rect 9150 -12106 9230 -12096
rect 9470 -12096 9480 -12086
rect 9540 -12096 9550 -12036
rect 9470 -12106 9550 -12096
rect 9150 -12376 9210 -12106
rect 9480 -12116 9550 -12106
rect 9290 -12166 9320 -12146
rect 9270 -12206 9320 -12166
rect 9380 -12166 9410 -12146
rect 9380 -12206 9430 -12166
rect 9270 -12276 9430 -12206
rect 9270 -12316 9320 -12276
rect 9290 -12336 9320 -12316
rect 9380 -12316 9430 -12276
rect 9380 -12336 9410 -12316
rect 9490 -12376 9550 -12116
rect 9150 -12386 9230 -12376
rect 9150 -12446 9160 -12386
rect 9220 -12396 9230 -12386
rect 9470 -12386 9550 -12376
rect 9470 -12396 9480 -12386
rect 9220 -12446 9480 -12396
rect 9540 -12446 9550 -12386
rect 9150 -12456 9550 -12446
rect 9606 -12036 10006 -12026
rect 9606 -12096 9616 -12036
rect 9676 -12086 9936 -12036
rect 9676 -12096 9686 -12086
rect 9606 -12106 9686 -12096
rect 9926 -12096 9936 -12086
rect 9996 -12096 10006 -12036
rect 9926 -12106 10006 -12096
rect 9606 -12376 9666 -12106
rect 9936 -12116 10006 -12106
rect 9746 -12166 9776 -12146
rect 9726 -12206 9776 -12166
rect 9836 -12166 9866 -12146
rect 9836 -12206 9886 -12166
rect 9726 -12276 9886 -12206
rect 9726 -12316 9776 -12276
rect 9746 -12336 9776 -12316
rect 9836 -12316 9886 -12276
rect 9836 -12336 9866 -12316
rect 9946 -12376 10006 -12116
rect 9606 -12386 9686 -12376
rect 9606 -12446 9616 -12386
rect 9676 -12396 9686 -12386
rect 9926 -12386 10006 -12376
rect 9926 -12396 9936 -12386
rect 9676 -12446 9936 -12396
rect 9996 -12446 10006 -12386
rect 9606 -12456 10006 -12446
rect 10062 -12036 10462 -12026
rect 10062 -12096 10072 -12036
rect 10132 -12086 10392 -12036
rect 10132 -12096 10142 -12086
rect 10062 -12106 10142 -12096
rect 10382 -12096 10392 -12086
rect 10452 -12096 10462 -12036
rect 10382 -12106 10462 -12096
rect 10062 -12376 10122 -12106
rect 10392 -12116 10462 -12106
rect 10202 -12166 10232 -12146
rect 10182 -12206 10232 -12166
rect 10292 -12166 10322 -12146
rect 10292 -12206 10342 -12166
rect 10182 -12276 10342 -12206
rect 10182 -12316 10232 -12276
rect 10202 -12336 10232 -12316
rect 10292 -12316 10342 -12276
rect 10292 -12336 10322 -12316
rect 10402 -12376 10462 -12116
rect 10062 -12386 10142 -12376
rect 10062 -12446 10072 -12386
rect 10132 -12396 10142 -12386
rect 10382 -12386 10462 -12376
rect 10382 -12396 10392 -12386
rect 10132 -12446 10392 -12396
rect 10452 -12446 10462 -12386
rect 10062 -12456 10462 -12446
rect 10520 -12036 10920 -12026
rect 10520 -12096 10530 -12036
rect 10590 -12086 10850 -12036
rect 10590 -12096 10600 -12086
rect 10520 -12106 10600 -12096
rect 10840 -12096 10850 -12086
rect 10910 -12096 10920 -12036
rect 10840 -12106 10920 -12096
rect 10520 -12376 10580 -12106
rect 10850 -12116 10920 -12106
rect 10660 -12166 10690 -12146
rect 10640 -12206 10690 -12166
rect 10750 -12166 10780 -12146
rect 10750 -12206 10800 -12166
rect 10640 -12276 10800 -12206
rect 10640 -12316 10690 -12276
rect 10660 -12336 10690 -12316
rect 10750 -12316 10800 -12276
rect 10750 -12336 10780 -12316
rect 10860 -12376 10920 -12116
rect 10520 -12386 10600 -12376
rect 10520 -12446 10530 -12386
rect 10590 -12396 10600 -12386
rect 10840 -12386 10920 -12376
rect 10840 -12396 10850 -12386
rect 10590 -12446 10850 -12396
rect 10910 -12446 10920 -12386
rect 10520 -12456 10920 -12446
rect 10976 -12036 11376 -12026
rect 10976 -12096 10986 -12036
rect 11046 -12086 11306 -12036
rect 11046 -12096 11056 -12086
rect 10976 -12106 11056 -12096
rect 11296 -12096 11306 -12086
rect 11366 -12096 11376 -12036
rect 11296 -12106 11376 -12096
rect 10976 -12376 11036 -12106
rect 11306 -12116 11376 -12106
rect 11116 -12166 11146 -12146
rect 11096 -12206 11146 -12166
rect 11206 -12166 11236 -12146
rect 11206 -12206 11256 -12166
rect 11096 -12276 11256 -12206
rect 11096 -12316 11146 -12276
rect 11116 -12336 11146 -12316
rect 11206 -12316 11256 -12276
rect 11206 -12336 11236 -12316
rect 11316 -12376 11376 -12116
rect 10976 -12386 11056 -12376
rect 10976 -12446 10986 -12386
rect 11046 -12396 11056 -12386
rect 11296 -12386 11376 -12376
rect 11296 -12396 11306 -12386
rect 11046 -12446 11306 -12396
rect 11366 -12446 11376 -12386
rect 10976 -12456 11376 -12446
rect 11432 -12036 11832 -12026
rect 11432 -12096 11442 -12036
rect 11502 -12086 11762 -12036
rect 11502 -12096 11512 -12086
rect 11432 -12106 11512 -12096
rect 11752 -12096 11762 -12086
rect 11822 -12096 11832 -12036
rect 11752 -12106 11832 -12096
rect 11432 -12376 11492 -12106
rect 11762 -12116 11832 -12106
rect 11572 -12166 11602 -12146
rect 11552 -12206 11602 -12166
rect 11662 -12166 11692 -12146
rect 11662 -12206 11712 -12166
rect 11552 -12276 11712 -12206
rect 11552 -12316 11602 -12276
rect 11572 -12336 11602 -12316
rect 11662 -12316 11712 -12276
rect 11662 -12336 11692 -12316
rect 11772 -12376 11832 -12116
rect 11432 -12386 11512 -12376
rect 11432 -12446 11442 -12386
rect 11502 -12396 11512 -12386
rect 11752 -12386 11832 -12376
rect 11752 -12396 11762 -12386
rect 11502 -12446 11762 -12396
rect 11822 -12446 11832 -12386
rect 11432 -12456 11832 -12446
rect 11890 -12036 12290 -12026
rect 11890 -12096 11900 -12036
rect 11960 -12086 12220 -12036
rect 11960 -12096 11970 -12086
rect 11890 -12106 11970 -12096
rect 12210 -12096 12220 -12086
rect 12280 -12096 12290 -12036
rect 12210 -12106 12290 -12096
rect 11890 -12376 11950 -12106
rect 12220 -12116 12290 -12106
rect 12030 -12166 12060 -12146
rect 12010 -12206 12060 -12166
rect 12120 -12166 12150 -12146
rect 12120 -12206 12170 -12166
rect 12010 -12276 12170 -12206
rect 12010 -12316 12060 -12276
rect 12030 -12336 12060 -12316
rect 12120 -12316 12170 -12276
rect 12120 -12336 12150 -12316
rect 12230 -12376 12290 -12116
rect 11890 -12386 11970 -12376
rect 11890 -12446 11900 -12386
rect 11960 -12396 11970 -12386
rect 12210 -12386 12290 -12376
rect 12210 -12396 12220 -12386
rect 11960 -12446 12220 -12396
rect 12280 -12446 12290 -12386
rect 11890 -12456 12290 -12446
rect 12346 -12036 12746 -12026
rect 12346 -12096 12356 -12036
rect 12416 -12086 12676 -12036
rect 12416 -12096 12426 -12086
rect 12346 -12106 12426 -12096
rect 12666 -12096 12676 -12086
rect 12736 -12096 12746 -12036
rect 12666 -12106 12746 -12096
rect 12346 -12376 12406 -12106
rect 12676 -12116 12746 -12106
rect 12486 -12166 12516 -12146
rect 12466 -12206 12516 -12166
rect 12576 -12166 12606 -12146
rect 12576 -12206 12626 -12166
rect 12466 -12276 12626 -12206
rect 12466 -12316 12516 -12276
rect 12486 -12336 12516 -12316
rect 12576 -12316 12626 -12276
rect 12576 -12336 12606 -12316
rect 12686 -12376 12746 -12116
rect 12346 -12386 12426 -12376
rect 12346 -12446 12356 -12386
rect 12416 -12396 12426 -12386
rect 12666 -12386 12746 -12376
rect 12666 -12396 12676 -12386
rect 12416 -12446 12676 -12396
rect 12736 -12446 12746 -12386
rect 12346 -12456 12746 -12446
rect 12802 -12036 13202 -12026
rect 12802 -12096 12812 -12036
rect 12872 -12086 13132 -12036
rect 12872 -12096 12882 -12086
rect 12802 -12106 12882 -12096
rect 13122 -12096 13132 -12086
rect 13192 -12096 13202 -12036
rect 13122 -12106 13202 -12096
rect 12802 -12376 12862 -12106
rect 13132 -12116 13202 -12106
rect 12942 -12166 12972 -12146
rect 12922 -12206 12972 -12166
rect 13032 -12166 13062 -12146
rect 13032 -12206 13082 -12166
rect 12922 -12276 13082 -12206
rect 12922 -12316 12972 -12276
rect 12942 -12336 12972 -12316
rect 13032 -12316 13082 -12276
rect 13032 -12336 13062 -12316
rect 13142 -12376 13202 -12116
rect 12802 -12386 12882 -12376
rect 12802 -12446 12812 -12386
rect 12872 -12396 12882 -12386
rect 13122 -12386 13202 -12376
rect 13122 -12396 13132 -12386
rect 12872 -12446 13132 -12396
rect 13192 -12446 13202 -12386
rect 12802 -12456 13202 -12446
rect 13260 -12036 13660 -12026
rect 13260 -12096 13270 -12036
rect 13330 -12086 13590 -12036
rect 13330 -12096 13340 -12086
rect 13260 -12106 13340 -12096
rect 13580 -12096 13590 -12086
rect 13650 -12096 13660 -12036
rect 13580 -12106 13660 -12096
rect 13260 -12376 13320 -12106
rect 13590 -12116 13660 -12106
rect 13400 -12166 13430 -12146
rect 13380 -12206 13430 -12166
rect 13490 -12166 13520 -12146
rect 13490 -12206 13540 -12166
rect 13380 -12276 13540 -12206
rect 13380 -12316 13430 -12276
rect 13400 -12336 13430 -12316
rect 13490 -12316 13540 -12276
rect 13490 -12336 13520 -12316
rect 13600 -12376 13660 -12116
rect 13260 -12386 13340 -12376
rect 13260 -12446 13270 -12386
rect 13330 -12396 13340 -12386
rect 13580 -12386 13660 -12376
rect 13580 -12396 13590 -12386
rect 13330 -12446 13590 -12396
rect 13650 -12446 13660 -12386
rect 13260 -12456 13660 -12446
rect 13716 -12036 14116 -12026
rect 13716 -12096 13726 -12036
rect 13786 -12086 14046 -12036
rect 13786 -12096 13796 -12086
rect 13716 -12106 13796 -12096
rect 14036 -12096 14046 -12086
rect 14106 -12096 14116 -12036
rect 14036 -12106 14116 -12096
rect 13716 -12376 13776 -12106
rect 14046 -12116 14116 -12106
rect 13856 -12166 13886 -12146
rect 13836 -12206 13886 -12166
rect 13946 -12166 13976 -12146
rect 13946 -12206 13996 -12166
rect 13836 -12276 13996 -12206
rect 13836 -12316 13886 -12276
rect 13856 -12336 13886 -12316
rect 13946 -12316 13996 -12276
rect 13946 -12336 13976 -12316
rect 14056 -12376 14116 -12116
rect 13716 -12386 13796 -12376
rect 13716 -12446 13726 -12386
rect 13786 -12396 13796 -12386
rect 14036 -12386 14116 -12376
rect 14036 -12396 14046 -12386
rect 13786 -12446 14046 -12396
rect 14106 -12446 14116 -12386
rect 13716 -12456 14116 -12446
rect 14172 -12036 14572 -12026
rect 14172 -12096 14182 -12036
rect 14242 -12086 14502 -12036
rect 14242 -12096 14252 -12086
rect 14172 -12106 14252 -12096
rect 14492 -12096 14502 -12086
rect 14562 -12096 14572 -12036
rect 14492 -12106 14572 -12096
rect 14172 -12376 14232 -12106
rect 14502 -12116 14572 -12106
rect 14312 -12166 14342 -12146
rect 14292 -12206 14342 -12166
rect 14402 -12166 14432 -12146
rect 14402 -12206 14452 -12166
rect 14292 -12276 14452 -12206
rect 14292 -12316 14342 -12276
rect 14312 -12336 14342 -12316
rect 14402 -12316 14452 -12276
rect 14402 -12336 14432 -12316
rect 14512 -12376 14572 -12116
rect 14172 -12386 14252 -12376
rect 14172 -12446 14182 -12386
rect 14242 -12396 14252 -12386
rect 14492 -12386 14572 -12376
rect 14492 -12396 14502 -12386
rect 14242 -12446 14502 -12396
rect 14562 -12446 14572 -12386
rect 14172 -12456 14572 -12446
rect 14630 -12036 15030 -12026
rect 14630 -12096 14640 -12036
rect 14700 -12086 14960 -12036
rect 14700 -12096 14710 -12086
rect 14630 -12106 14710 -12096
rect 14950 -12096 14960 -12086
rect 15020 -12096 15030 -12036
rect 14950 -12106 15030 -12096
rect 14630 -12376 14690 -12106
rect 14960 -12116 15030 -12106
rect 14770 -12166 14800 -12146
rect 14750 -12206 14800 -12166
rect 14860 -12166 14890 -12146
rect 14860 -12206 14910 -12166
rect 14750 -12276 14910 -12206
rect 14750 -12316 14800 -12276
rect 14770 -12336 14800 -12316
rect 14860 -12316 14910 -12276
rect 14860 -12336 14890 -12316
rect 14970 -12376 15030 -12116
rect 14630 -12386 14710 -12376
rect 14630 -12446 14640 -12386
rect 14700 -12396 14710 -12386
rect 14950 -12386 15030 -12376
rect 14950 -12396 14960 -12386
rect 14700 -12446 14960 -12396
rect 15020 -12446 15030 -12386
rect 14630 -12456 15030 -12446
rect 15086 -12036 15486 -12026
rect 15086 -12096 15096 -12036
rect 15156 -12086 15416 -12036
rect 15156 -12096 15166 -12086
rect 15086 -12106 15166 -12096
rect 15406 -12096 15416 -12086
rect 15476 -12096 15486 -12036
rect 15406 -12106 15486 -12096
rect 15086 -12376 15146 -12106
rect 15416 -12116 15486 -12106
rect 15226 -12166 15256 -12146
rect 15206 -12206 15256 -12166
rect 15316 -12166 15346 -12146
rect 15316 -12206 15366 -12166
rect 15206 -12276 15366 -12206
rect 15206 -12316 15256 -12276
rect 15226 -12336 15256 -12316
rect 15316 -12316 15366 -12276
rect 15316 -12336 15346 -12316
rect 15426 -12376 15486 -12116
rect 15086 -12386 15166 -12376
rect 15086 -12446 15096 -12386
rect 15156 -12396 15166 -12386
rect 15406 -12386 15486 -12376
rect 15406 -12396 15416 -12386
rect 15156 -12446 15416 -12396
rect 15476 -12446 15486 -12386
rect 15086 -12456 15486 -12446
rect 0 -12552 400 -12542
rect 0 -12612 10 -12552
rect 70 -12602 330 -12552
rect 70 -12612 80 -12602
rect 0 -12622 80 -12612
rect 320 -12612 330 -12602
rect 390 -12612 400 -12552
rect 320 -12622 400 -12612
rect 0 -12892 60 -12622
rect 330 -12632 400 -12622
rect 140 -12682 170 -12662
rect 120 -12722 170 -12682
rect 230 -12682 260 -12662
rect 230 -12722 280 -12682
rect 120 -12792 280 -12722
rect 120 -12832 170 -12792
rect 140 -12852 170 -12832
rect 230 -12832 280 -12792
rect 230 -12852 260 -12832
rect 340 -12892 400 -12632
rect 0 -12902 80 -12892
rect 0 -12962 10 -12902
rect 70 -12912 80 -12902
rect 320 -12902 400 -12892
rect 320 -12912 330 -12902
rect 70 -12962 330 -12912
rect 390 -12962 400 -12902
rect 0 -12972 400 -12962
rect 456 -12552 856 -12542
rect 456 -12612 466 -12552
rect 526 -12602 786 -12552
rect 526 -12612 536 -12602
rect 456 -12622 536 -12612
rect 776 -12612 786 -12602
rect 846 -12612 856 -12552
rect 776 -12622 856 -12612
rect 456 -12892 516 -12622
rect 786 -12632 856 -12622
rect 596 -12682 626 -12662
rect 576 -12722 626 -12682
rect 686 -12682 716 -12662
rect 686 -12722 736 -12682
rect 576 -12792 736 -12722
rect 576 -12832 626 -12792
rect 596 -12852 626 -12832
rect 686 -12832 736 -12792
rect 686 -12852 716 -12832
rect 796 -12892 856 -12632
rect 456 -12902 536 -12892
rect 456 -12962 466 -12902
rect 526 -12912 536 -12902
rect 776 -12902 856 -12892
rect 776 -12912 786 -12902
rect 526 -12962 786 -12912
rect 846 -12962 856 -12902
rect 456 -12972 856 -12962
rect 912 -12552 1312 -12542
rect 912 -12612 922 -12552
rect 982 -12602 1242 -12552
rect 982 -12612 992 -12602
rect 912 -12622 992 -12612
rect 1232 -12612 1242 -12602
rect 1302 -12612 1312 -12552
rect 1232 -12622 1312 -12612
rect 912 -12892 972 -12622
rect 1242 -12632 1312 -12622
rect 1052 -12682 1082 -12662
rect 1032 -12722 1082 -12682
rect 1142 -12682 1172 -12662
rect 1142 -12722 1192 -12682
rect 1032 -12792 1192 -12722
rect 1032 -12832 1082 -12792
rect 1052 -12852 1082 -12832
rect 1142 -12832 1192 -12792
rect 1142 -12852 1172 -12832
rect 1252 -12892 1312 -12632
rect 912 -12902 992 -12892
rect 912 -12962 922 -12902
rect 982 -12912 992 -12902
rect 1232 -12902 1312 -12892
rect 1232 -12912 1242 -12902
rect 982 -12962 1242 -12912
rect 1302 -12962 1312 -12902
rect 912 -12972 1312 -12962
rect 1370 -12552 1770 -12542
rect 1370 -12612 1380 -12552
rect 1440 -12602 1700 -12552
rect 1440 -12612 1450 -12602
rect 1370 -12622 1450 -12612
rect 1690 -12612 1700 -12602
rect 1760 -12612 1770 -12552
rect 1690 -12622 1770 -12612
rect 1370 -12892 1430 -12622
rect 1700 -12632 1770 -12622
rect 1510 -12682 1540 -12662
rect 1490 -12722 1540 -12682
rect 1600 -12682 1630 -12662
rect 1600 -12722 1650 -12682
rect 1490 -12792 1650 -12722
rect 1490 -12832 1540 -12792
rect 1510 -12852 1540 -12832
rect 1600 -12832 1650 -12792
rect 1600 -12852 1630 -12832
rect 1710 -12892 1770 -12632
rect 1370 -12902 1450 -12892
rect 1370 -12962 1380 -12902
rect 1440 -12912 1450 -12902
rect 1690 -12902 1770 -12892
rect 1690 -12912 1700 -12902
rect 1440 -12962 1700 -12912
rect 1760 -12962 1770 -12902
rect 1370 -12972 1770 -12962
rect 1826 -12552 2226 -12542
rect 1826 -12612 1836 -12552
rect 1896 -12602 2156 -12552
rect 1896 -12612 1906 -12602
rect 1826 -12622 1906 -12612
rect 2146 -12612 2156 -12602
rect 2216 -12612 2226 -12552
rect 2146 -12622 2226 -12612
rect 1826 -12892 1886 -12622
rect 2156 -12632 2226 -12622
rect 1966 -12682 1996 -12662
rect 1946 -12722 1996 -12682
rect 2056 -12682 2086 -12662
rect 2056 -12722 2106 -12682
rect 1946 -12792 2106 -12722
rect 1946 -12832 1996 -12792
rect 1966 -12852 1996 -12832
rect 2056 -12832 2106 -12792
rect 2056 -12852 2086 -12832
rect 2166 -12892 2226 -12632
rect 1826 -12902 1906 -12892
rect 1826 -12962 1836 -12902
rect 1896 -12912 1906 -12902
rect 2146 -12902 2226 -12892
rect 2146 -12912 2156 -12902
rect 1896 -12962 2156 -12912
rect 2216 -12962 2226 -12902
rect 1826 -12972 2226 -12962
rect 2282 -12552 2682 -12542
rect 2282 -12612 2292 -12552
rect 2352 -12602 2612 -12552
rect 2352 -12612 2362 -12602
rect 2282 -12622 2362 -12612
rect 2602 -12612 2612 -12602
rect 2672 -12612 2682 -12552
rect 2602 -12622 2682 -12612
rect 2282 -12892 2342 -12622
rect 2612 -12632 2682 -12622
rect 2422 -12682 2452 -12662
rect 2402 -12722 2452 -12682
rect 2512 -12682 2542 -12662
rect 2512 -12722 2562 -12682
rect 2402 -12792 2562 -12722
rect 2402 -12832 2452 -12792
rect 2422 -12852 2452 -12832
rect 2512 -12832 2562 -12792
rect 2512 -12852 2542 -12832
rect 2622 -12892 2682 -12632
rect 2282 -12902 2362 -12892
rect 2282 -12962 2292 -12902
rect 2352 -12912 2362 -12902
rect 2602 -12902 2682 -12892
rect 2602 -12912 2612 -12902
rect 2352 -12962 2612 -12912
rect 2672 -12962 2682 -12902
rect 2282 -12972 2682 -12962
rect 2740 -12552 3140 -12542
rect 2740 -12612 2750 -12552
rect 2810 -12602 3070 -12552
rect 2810 -12612 2820 -12602
rect 2740 -12622 2820 -12612
rect 3060 -12612 3070 -12602
rect 3130 -12612 3140 -12552
rect 3060 -12622 3140 -12612
rect 2740 -12892 2800 -12622
rect 3070 -12632 3140 -12622
rect 2880 -12682 2910 -12662
rect 2860 -12722 2910 -12682
rect 2970 -12682 3000 -12662
rect 2970 -12722 3020 -12682
rect 2860 -12792 3020 -12722
rect 2860 -12832 2910 -12792
rect 2880 -12852 2910 -12832
rect 2970 -12832 3020 -12792
rect 2970 -12852 3000 -12832
rect 3080 -12892 3140 -12632
rect 2740 -12902 2820 -12892
rect 2740 -12962 2750 -12902
rect 2810 -12912 2820 -12902
rect 3060 -12902 3140 -12892
rect 3060 -12912 3070 -12902
rect 2810 -12962 3070 -12912
rect 3130 -12962 3140 -12902
rect 2740 -12972 3140 -12962
rect 3196 -12552 3596 -12542
rect 3196 -12612 3206 -12552
rect 3266 -12602 3526 -12552
rect 3266 -12612 3276 -12602
rect 3196 -12622 3276 -12612
rect 3516 -12612 3526 -12602
rect 3586 -12612 3596 -12552
rect 3516 -12622 3596 -12612
rect 3196 -12892 3256 -12622
rect 3526 -12632 3596 -12622
rect 3336 -12682 3366 -12662
rect 3316 -12722 3366 -12682
rect 3426 -12682 3456 -12662
rect 3426 -12722 3476 -12682
rect 3316 -12792 3476 -12722
rect 3316 -12832 3366 -12792
rect 3336 -12852 3366 -12832
rect 3426 -12832 3476 -12792
rect 3426 -12852 3456 -12832
rect 3536 -12892 3596 -12632
rect 3196 -12902 3276 -12892
rect 3196 -12962 3206 -12902
rect 3266 -12912 3276 -12902
rect 3516 -12902 3596 -12892
rect 3516 -12912 3526 -12902
rect 3266 -12962 3526 -12912
rect 3586 -12962 3596 -12902
rect 3196 -12972 3596 -12962
rect 3652 -12552 4052 -12542
rect 3652 -12612 3662 -12552
rect 3722 -12602 3982 -12552
rect 3722 -12612 3732 -12602
rect 3652 -12622 3732 -12612
rect 3972 -12612 3982 -12602
rect 4042 -12612 4052 -12552
rect 3972 -12622 4052 -12612
rect 3652 -12892 3712 -12622
rect 3982 -12632 4052 -12622
rect 3792 -12682 3822 -12662
rect 3772 -12722 3822 -12682
rect 3882 -12682 3912 -12662
rect 3882 -12722 3932 -12682
rect 3772 -12792 3932 -12722
rect 3772 -12832 3822 -12792
rect 3792 -12852 3822 -12832
rect 3882 -12832 3932 -12792
rect 3882 -12852 3912 -12832
rect 3992 -12892 4052 -12632
rect 3652 -12902 3732 -12892
rect 3652 -12962 3662 -12902
rect 3722 -12912 3732 -12902
rect 3972 -12902 4052 -12892
rect 3972 -12912 3982 -12902
rect 3722 -12962 3982 -12912
rect 4042 -12962 4052 -12902
rect 3652 -12972 4052 -12962
rect 4110 -12552 4510 -12542
rect 4110 -12612 4120 -12552
rect 4180 -12602 4440 -12552
rect 4180 -12612 4190 -12602
rect 4110 -12622 4190 -12612
rect 4430 -12612 4440 -12602
rect 4500 -12612 4510 -12552
rect 4430 -12622 4510 -12612
rect 4110 -12892 4170 -12622
rect 4440 -12632 4510 -12622
rect 4250 -12682 4280 -12662
rect 4230 -12722 4280 -12682
rect 4340 -12682 4370 -12662
rect 4340 -12722 4390 -12682
rect 4230 -12792 4390 -12722
rect 4230 -12832 4280 -12792
rect 4250 -12852 4280 -12832
rect 4340 -12832 4390 -12792
rect 4340 -12852 4370 -12832
rect 4450 -12892 4510 -12632
rect 4110 -12902 4190 -12892
rect 4110 -12962 4120 -12902
rect 4180 -12912 4190 -12902
rect 4430 -12902 4510 -12892
rect 4430 -12912 4440 -12902
rect 4180 -12962 4440 -12912
rect 4500 -12962 4510 -12902
rect 4110 -12972 4510 -12962
rect 4566 -12552 4966 -12542
rect 4566 -12612 4576 -12552
rect 4636 -12602 4896 -12552
rect 4636 -12612 4646 -12602
rect 4566 -12622 4646 -12612
rect 4886 -12612 4896 -12602
rect 4956 -12612 4966 -12552
rect 4886 -12622 4966 -12612
rect 4566 -12892 4626 -12622
rect 4896 -12632 4966 -12622
rect 4706 -12682 4736 -12662
rect 4686 -12722 4736 -12682
rect 4796 -12682 4826 -12662
rect 4796 -12722 4846 -12682
rect 4686 -12792 4846 -12722
rect 4686 -12832 4736 -12792
rect 4706 -12852 4736 -12832
rect 4796 -12832 4846 -12792
rect 4796 -12852 4826 -12832
rect 4906 -12892 4966 -12632
rect 4566 -12902 4646 -12892
rect 4566 -12962 4576 -12902
rect 4636 -12912 4646 -12902
rect 4886 -12902 4966 -12892
rect 4886 -12912 4896 -12902
rect 4636 -12962 4896 -12912
rect 4956 -12962 4966 -12902
rect 4566 -12972 4966 -12962
rect 5022 -12552 5422 -12542
rect 5022 -12612 5032 -12552
rect 5092 -12602 5352 -12552
rect 5092 -12612 5102 -12602
rect 5022 -12622 5102 -12612
rect 5342 -12612 5352 -12602
rect 5412 -12612 5422 -12552
rect 5342 -12622 5422 -12612
rect 5022 -12892 5082 -12622
rect 5352 -12632 5422 -12622
rect 5162 -12682 5192 -12662
rect 5142 -12722 5192 -12682
rect 5252 -12682 5282 -12662
rect 5252 -12722 5302 -12682
rect 5142 -12792 5302 -12722
rect 5142 -12832 5192 -12792
rect 5162 -12852 5192 -12832
rect 5252 -12832 5302 -12792
rect 5252 -12852 5282 -12832
rect 5362 -12892 5422 -12632
rect 5022 -12902 5102 -12892
rect 5022 -12962 5032 -12902
rect 5092 -12912 5102 -12902
rect 5342 -12902 5422 -12892
rect 5342 -12912 5352 -12902
rect 5092 -12962 5352 -12912
rect 5412 -12962 5422 -12902
rect 5022 -12972 5422 -12962
rect 5480 -12552 5880 -12542
rect 5480 -12612 5490 -12552
rect 5550 -12602 5810 -12552
rect 5550 -12612 5560 -12602
rect 5480 -12622 5560 -12612
rect 5800 -12612 5810 -12602
rect 5870 -12612 5880 -12552
rect 5800 -12622 5880 -12612
rect 5480 -12892 5540 -12622
rect 5810 -12632 5880 -12622
rect 5620 -12682 5650 -12662
rect 5600 -12722 5650 -12682
rect 5710 -12682 5740 -12662
rect 5710 -12722 5760 -12682
rect 5600 -12792 5760 -12722
rect 5600 -12832 5650 -12792
rect 5620 -12852 5650 -12832
rect 5710 -12832 5760 -12792
rect 5710 -12852 5740 -12832
rect 5820 -12892 5880 -12632
rect 5480 -12902 5560 -12892
rect 5480 -12962 5490 -12902
rect 5550 -12912 5560 -12902
rect 5800 -12902 5880 -12892
rect 5800 -12912 5810 -12902
rect 5550 -12962 5810 -12912
rect 5870 -12962 5880 -12902
rect 5480 -12972 5880 -12962
rect 5936 -12552 6336 -12542
rect 5936 -12612 5946 -12552
rect 6006 -12602 6266 -12552
rect 6006 -12612 6016 -12602
rect 5936 -12622 6016 -12612
rect 6256 -12612 6266 -12602
rect 6326 -12612 6336 -12552
rect 6256 -12622 6336 -12612
rect 5936 -12892 5996 -12622
rect 6266 -12632 6336 -12622
rect 6076 -12682 6106 -12662
rect 6056 -12722 6106 -12682
rect 6166 -12682 6196 -12662
rect 6166 -12722 6216 -12682
rect 6056 -12792 6216 -12722
rect 6056 -12832 6106 -12792
rect 6076 -12852 6106 -12832
rect 6166 -12832 6216 -12792
rect 6166 -12852 6196 -12832
rect 6276 -12892 6336 -12632
rect 5936 -12902 6016 -12892
rect 5936 -12962 5946 -12902
rect 6006 -12912 6016 -12902
rect 6256 -12902 6336 -12892
rect 6256 -12912 6266 -12902
rect 6006 -12962 6266 -12912
rect 6326 -12962 6336 -12902
rect 5936 -12972 6336 -12962
rect 6392 -12552 6792 -12542
rect 6392 -12612 6402 -12552
rect 6462 -12602 6722 -12552
rect 6462 -12612 6472 -12602
rect 6392 -12622 6472 -12612
rect 6712 -12612 6722 -12602
rect 6782 -12612 6792 -12552
rect 6712 -12622 6792 -12612
rect 6392 -12892 6452 -12622
rect 6722 -12632 6792 -12622
rect 6532 -12682 6562 -12662
rect 6512 -12722 6562 -12682
rect 6622 -12682 6652 -12662
rect 6622 -12722 6672 -12682
rect 6512 -12792 6672 -12722
rect 6512 -12832 6562 -12792
rect 6532 -12852 6562 -12832
rect 6622 -12832 6672 -12792
rect 6622 -12852 6652 -12832
rect 6732 -12892 6792 -12632
rect 6392 -12902 6472 -12892
rect 6392 -12962 6402 -12902
rect 6462 -12912 6472 -12902
rect 6712 -12902 6792 -12892
rect 6712 -12912 6722 -12902
rect 6462 -12962 6722 -12912
rect 6782 -12962 6792 -12902
rect 6392 -12972 6792 -12962
rect 6850 -12552 7250 -12542
rect 6850 -12612 6860 -12552
rect 6920 -12602 7180 -12552
rect 6920 -12612 6930 -12602
rect 6850 -12622 6930 -12612
rect 7170 -12612 7180 -12602
rect 7240 -12612 7250 -12552
rect 7170 -12622 7250 -12612
rect 6850 -12892 6910 -12622
rect 7180 -12632 7250 -12622
rect 6990 -12682 7020 -12662
rect 6970 -12722 7020 -12682
rect 7080 -12682 7110 -12662
rect 7080 -12722 7130 -12682
rect 6970 -12792 7130 -12722
rect 6970 -12832 7020 -12792
rect 6990 -12852 7020 -12832
rect 7080 -12832 7130 -12792
rect 7080 -12852 7110 -12832
rect 7190 -12892 7250 -12632
rect 6850 -12902 6930 -12892
rect 6850 -12962 6860 -12902
rect 6920 -12912 6930 -12902
rect 7170 -12902 7250 -12892
rect 7170 -12912 7180 -12902
rect 6920 -12962 7180 -12912
rect 7240 -12962 7250 -12902
rect 6850 -12972 7250 -12962
rect 7306 -12552 7706 -12542
rect 7306 -12612 7316 -12552
rect 7376 -12602 7636 -12552
rect 7376 -12612 7386 -12602
rect 7306 -12622 7386 -12612
rect 7626 -12612 7636 -12602
rect 7696 -12612 7706 -12552
rect 7626 -12622 7706 -12612
rect 7306 -12892 7366 -12622
rect 7636 -12632 7706 -12622
rect 7446 -12682 7476 -12662
rect 7426 -12722 7476 -12682
rect 7536 -12682 7566 -12662
rect 7536 -12722 7586 -12682
rect 7426 -12792 7586 -12722
rect 7426 -12832 7476 -12792
rect 7446 -12852 7476 -12832
rect 7536 -12832 7586 -12792
rect 7536 -12852 7566 -12832
rect 7646 -12892 7706 -12632
rect 7306 -12902 7386 -12892
rect 7306 -12962 7316 -12902
rect 7376 -12912 7386 -12902
rect 7626 -12902 7706 -12892
rect 7626 -12912 7636 -12902
rect 7376 -12962 7636 -12912
rect 7696 -12962 7706 -12902
rect 7306 -12972 7706 -12962
rect 7762 -12552 8162 -12542
rect 7762 -12612 7772 -12552
rect 7832 -12602 8092 -12552
rect 7832 -12612 7842 -12602
rect 7762 -12622 7842 -12612
rect 8082 -12612 8092 -12602
rect 8152 -12612 8162 -12552
rect 8082 -12622 8162 -12612
rect 7762 -12892 7822 -12622
rect 8092 -12632 8162 -12622
rect 7902 -12682 7932 -12662
rect 7882 -12722 7932 -12682
rect 7992 -12682 8022 -12662
rect 7992 -12722 8042 -12682
rect 7882 -12792 8042 -12722
rect 7882 -12832 7932 -12792
rect 7902 -12852 7932 -12832
rect 7992 -12832 8042 -12792
rect 7992 -12852 8022 -12832
rect 8102 -12892 8162 -12632
rect 7762 -12902 7842 -12892
rect 7762 -12962 7772 -12902
rect 7832 -12912 7842 -12902
rect 8082 -12902 8162 -12892
rect 8082 -12912 8092 -12902
rect 7832 -12962 8092 -12912
rect 8152 -12962 8162 -12902
rect 7762 -12972 8162 -12962
rect 8236 -12552 8636 -12542
rect 8236 -12612 8246 -12552
rect 8306 -12602 8566 -12552
rect 8306 -12612 8316 -12602
rect 8236 -12622 8316 -12612
rect 8556 -12612 8566 -12602
rect 8626 -12612 8636 -12552
rect 8556 -12622 8636 -12612
rect 8236 -12892 8296 -12622
rect 8566 -12632 8636 -12622
rect 8376 -12682 8406 -12662
rect 8356 -12722 8406 -12682
rect 8466 -12682 8496 -12662
rect 8466 -12722 8516 -12682
rect 8356 -12792 8516 -12722
rect 8356 -12832 8406 -12792
rect 8376 -12852 8406 -12832
rect 8466 -12832 8516 -12792
rect 8466 -12852 8496 -12832
rect 8576 -12892 8636 -12632
rect 8236 -12902 8316 -12892
rect 8236 -12962 8246 -12902
rect 8306 -12912 8316 -12902
rect 8556 -12902 8636 -12892
rect 8556 -12912 8566 -12902
rect 8306 -12962 8566 -12912
rect 8626 -12962 8636 -12902
rect 8236 -12972 8636 -12962
rect 8692 -12552 9092 -12542
rect 8692 -12612 8702 -12552
rect 8762 -12602 9022 -12552
rect 8762 -12612 8772 -12602
rect 8692 -12622 8772 -12612
rect 9012 -12612 9022 -12602
rect 9082 -12612 9092 -12552
rect 9012 -12622 9092 -12612
rect 8692 -12892 8752 -12622
rect 9022 -12632 9092 -12622
rect 8832 -12682 8862 -12662
rect 8812 -12722 8862 -12682
rect 8922 -12682 8952 -12662
rect 8922 -12722 8972 -12682
rect 8812 -12792 8972 -12722
rect 8812 -12832 8862 -12792
rect 8832 -12852 8862 -12832
rect 8922 -12832 8972 -12792
rect 8922 -12852 8952 -12832
rect 9032 -12892 9092 -12632
rect 8692 -12902 8772 -12892
rect 8692 -12962 8702 -12902
rect 8762 -12912 8772 -12902
rect 9012 -12902 9092 -12892
rect 9012 -12912 9022 -12902
rect 8762 -12962 9022 -12912
rect 9082 -12962 9092 -12902
rect 8692 -12972 9092 -12962
rect 9150 -12552 9550 -12542
rect 9150 -12612 9160 -12552
rect 9220 -12602 9480 -12552
rect 9220 -12612 9230 -12602
rect 9150 -12622 9230 -12612
rect 9470 -12612 9480 -12602
rect 9540 -12612 9550 -12552
rect 9470 -12622 9550 -12612
rect 9150 -12892 9210 -12622
rect 9480 -12632 9550 -12622
rect 9290 -12682 9320 -12662
rect 9270 -12722 9320 -12682
rect 9380 -12682 9410 -12662
rect 9380 -12722 9430 -12682
rect 9270 -12792 9430 -12722
rect 9270 -12832 9320 -12792
rect 9290 -12852 9320 -12832
rect 9380 -12832 9430 -12792
rect 9380 -12852 9410 -12832
rect 9490 -12892 9550 -12632
rect 9150 -12902 9230 -12892
rect 9150 -12962 9160 -12902
rect 9220 -12912 9230 -12902
rect 9470 -12902 9550 -12892
rect 9470 -12912 9480 -12902
rect 9220 -12962 9480 -12912
rect 9540 -12962 9550 -12902
rect 9150 -12972 9550 -12962
rect 9606 -12552 10006 -12542
rect 9606 -12612 9616 -12552
rect 9676 -12602 9936 -12552
rect 9676 -12612 9686 -12602
rect 9606 -12622 9686 -12612
rect 9926 -12612 9936 -12602
rect 9996 -12612 10006 -12552
rect 9926 -12622 10006 -12612
rect 9606 -12892 9666 -12622
rect 9936 -12632 10006 -12622
rect 9746 -12682 9776 -12662
rect 9726 -12722 9776 -12682
rect 9836 -12682 9866 -12662
rect 9836 -12722 9886 -12682
rect 9726 -12792 9886 -12722
rect 9726 -12832 9776 -12792
rect 9746 -12852 9776 -12832
rect 9836 -12832 9886 -12792
rect 9836 -12852 9866 -12832
rect 9946 -12892 10006 -12632
rect 9606 -12902 9686 -12892
rect 9606 -12962 9616 -12902
rect 9676 -12912 9686 -12902
rect 9926 -12902 10006 -12892
rect 9926 -12912 9936 -12902
rect 9676 -12962 9936 -12912
rect 9996 -12962 10006 -12902
rect 9606 -12972 10006 -12962
rect 10062 -12552 10462 -12542
rect 10062 -12612 10072 -12552
rect 10132 -12602 10392 -12552
rect 10132 -12612 10142 -12602
rect 10062 -12622 10142 -12612
rect 10382 -12612 10392 -12602
rect 10452 -12612 10462 -12552
rect 10382 -12622 10462 -12612
rect 10062 -12892 10122 -12622
rect 10392 -12632 10462 -12622
rect 10202 -12682 10232 -12662
rect 10182 -12722 10232 -12682
rect 10292 -12682 10322 -12662
rect 10292 -12722 10342 -12682
rect 10182 -12792 10342 -12722
rect 10182 -12832 10232 -12792
rect 10202 -12852 10232 -12832
rect 10292 -12832 10342 -12792
rect 10292 -12852 10322 -12832
rect 10402 -12892 10462 -12632
rect 10062 -12902 10142 -12892
rect 10062 -12962 10072 -12902
rect 10132 -12912 10142 -12902
rect 10382 -12902 10462 -12892
rect 10382 -12912 10392 -12902
rect 10132 -12962 10392 -12912
rect 10452 -12962 10462 -12902
rect 10062 -12972 10462 -12962
rect 10520 -12552 10920 -12542
rect 10520 -12612 10530 -12552
rect 10590 -12602 10850 -12552
rect 10590 -12612 10600 -12602
rect 10520 -12622 10600 -12612
rect 10840 -12612 10850 -12602
rect 10910 -12612 10920 -12552
rect 10840 -12622 10920 -12612
rect 10520 -12892 10580 -12622
rect 10850 -12632 10920 -12622
rect 10660 -12682 10690 -12662
rect 10640 -12722 10690 -12682
rect 10750 -12682 10780 -12662
rect 10750 -12722 10800 -12682
rect 10640 -12792 10800 -12722
rect 10640 -12832 10690 -12792
rect 10660 -12852 10690 -12832
rect 10750 -12832 10800 -12792
rect 10750 -12852 10780 -12832
rect 10860 -12892 10920 -12632
rect 10520 -12902 10600 -12892
rect 10520 -12962 10530 -12902
rect 10590 -12912 10600 -12902
rect 10840 -12902 10920 -12892
rect 10840 -12912 10850 -12902
rect 10590 -12962 10850 -12912
rect 10910 -12962 10920 -12902
rect 10520 -12972 10920 -12962
rect 10976 -12552 11376 -12542
rect 10976 -12612 10986 -12552
rect 11046 -12602 11306 -12552
rect 11046 -12612 11056 -12602
rect 10976 -12622 11056 -12612
rect 11296 -12612 11306 -12602
rect 11366 -12612 11376 -12552
rect 11296 -12622 11376 -12612
rect 10976 -12892 11036 -12622
rect 11306 -12632 11376 -12622
rect 11116 -12682 11146 -12662
rect 11096 -12722 11146 -12682
rect 11206 -12682 11236 -12662
rect 11206 -12722 11256 -12682
rect 11096 -12792 11256 -12722
rect 11096 -12832 11146 -12792
rect 11116 -12852 11146 -12832
rect 11206 -12832 11256 -12792
rect 11206 -12852 11236 -12832
rect 11316 -12892 11376 -12632
rect 10976 -12902 11056 -12892
rect 10976 -12962 10986 -12902
rect 11046 -12912 11056 -12902
rect 11296 -12902 11376 -12892
rect 11296 -12912 11306 -12902
rect 11046 -12962 11306 -12912
rect 11366 -12962 11376 -12902
rect 10976 -12972 11376 -12962
rect 11432 -12552 11832 -12542
rect 11432 -12612 11442 -12552
rect 11502 -12602 11762 -12552
rect 11502 -12612 11512 -12602
rect 11432 -12622 11512 -12612
rect 11752 -12612 11762 -12602
rect 11822 -12612 11832 -12552
rect 11752 -12622 11832 -12612
rect 11432 -12892 11492 -12622
rect 11762 -12632 11832 -12622
rect 11572 -12682 11602 -12662
rect 11552 -12722 11602 -12682
rect 11662 -12682 11692 -12662
rect 11662 -12722 11712 -12682
rect 11552 -12792 11712 -12722
rect 11552 -12832 11602 -12792
rect 11572 -12852 11602 -12832
rect 11662 -12832 11712 -12792
rect 11662 -12852 11692 -12832
rect 11772 -12892 11832 -12632
rect 11432 -12902 11512 -12892
rect 11432 -12962 11442 -12902
rect 11502 -12912 11512 -12902
rect 11752 -12902 11832 -12892
rect 11752 -12912 11762 -12902
rect 11502 -12962 11762 -12912
rect 11822 -12962 11832 -12902
rect 11432 -12972 11832 -12962
rect 11890 -12552 12290 -12542
rect 11890 -12612 11900 -12552
rect 11960 -12602 12220 -12552
rect 11960 -12612 11970 -12602
rect 11890 -12622 11970 -12612
rect 12210 -12612 12220 -12602
rect 12280 -12612 12290 -12552
rect 12210 -12622 12290 -12612
rect 11890 -12892 11950 -12622
rect 12220 -12632 12290 -12622
rect 12030 -12682 12060 -12662
rect 12010 -12722 12060 -12682
rect 12120 -12682 12150 -12662
rect 12120 -12722 12170 -12682
rect 12010 -12792 12170 -12722
rect 12010 -12832 12060 -12792
rect 12030 -12852 12060 -12832
rect 12120 -12832 12170 -12792
rect 12120 -12852 12150 -12832
rect 12230 -12892 12290 -12632
rect 11890 -12902 11970 -12892
rect 11890 -12962 11900 -12902
rect 11960 -12912 11970 -12902
rect 12210 -12902 12290 -12892
rect 12210 -12912 12220 -12902
rect 11960 -12962 12220 -12912
rect 12280 -12962 12290 -12902
rect 11890 -12972 12290 -12962
rect 12346 -12552 12746 -12542
rect 12346 -12612 12356 -12552
rect 12416 -12602 12676 -12552
rect 12416 -12612 12426 -12602
rect 12346 -12622 12426 -12612
rect 12666 -12612 12676 -12602
rect 12736 -12612 12746 -12552
rect 12666 -12622 12746 -12612
rect 12346 -12892 12406 -12622
rect 12676 -12632 12746 -12622
rect 12486 -12682 12516 -12662
rect 12466 -12722 12516 -12682
rect 12576 -12682 12606 -12662
rect 12576 -12722 12626 -12682
rect 12466 -12792 12626 -12722
rect 12466 -12832 12516 -12792
rect 12486 -12852 12516 -12832
rect 12576 -12832 12626 -12792
rect 12576 -12852 12606 -12832
rect 12686 -12892 12746 -12632
rect 12346 -12902 12426 -12892
rect 12346 -12962 12356 -12902
rect 12416 -12912 12426 -12902
rect 12666 -12902 12746 -12892
rect 12666 -12912 12676 -12902
rect 12416 -12962 12676 -12912
rect 12736 -12962 12746 -12902
rect 12346 -12972 12746 -12962
rect 12802 -12552 13202 -12542
rect 12802 -12612 12812 -12552
rect 12872 -12602 13132 -12552
rect 12872 -12612 12882 -12602
rect 12802 -12622 12882 -12612
rect 13122 -12612 13132 -12602
rect 13192 -12612 13202 -12552
rect 13122 -12622 13202 -12612
rect 12802 -12892 12862 -12622
rect 13132 -12632 13202 -12622
rect 12942 -12682 12972 -12662
rect 12922 -12722 12972 -12682
rect 13032 -12682 13062 -12662
rect 13032 -12722 13082 -12682
rect 12922 -12792 13082 -12722
rect 12922 -12832 12972 -12792
rect 12942 -12852 12972 -12832
rect 13032 -12832 13082 -12792
rect 13032 -12852 13062 -12832
rect 13142 -12892 13202 -12632
rect 12802 -12902 12882 -12892
rect 12802 -12962 12812 -12902
rect 12872 -12912 12882 -12902
rect 13122 -12902 13202 -12892
rect 13122 -12912 13132 -12902
rect 12872 -12962 13132 -12912
rect 13192 -12962 13202 -12902
rect 12802 -12972 13202 -12962
rect 13260 -12552 13660 -12542
rect 13260 -12612 13270 -12552
rect 13330 -12602 13590 -12552
rect 13330 -12612 13340 -12602
rect 13260 -12622 13340 -12612
rect 13580 -12612 13590 -12602
rect 13650 -12612 13660 -12552
rect 13580 -12622 13660 -12612
rect 13260 -12892 13320 -12622
rect 13590 -12632 13660 -12622
rect 13400 -12682 13430 -12662
rect 13380 -12722 13430 -12682
rect 13490 -12682 13520 -12662
rect 13490 -12722 13540 -12682
rect 13380 -12792 13540 -12722
rect 13380 -12832 13430 -12792
rect 13400 -12852 13430 -12832
rect 13490 -12832 13540 -12792
rect 13490 -12852 13520 -12832
rect 13600 -12892 13660 -12632
rect 13260 -12902 13340 -12892
rect 13260 -12962 13270 -12902
rect 13330 -12912 13340 -12902
rect 13580 -12902 13660 -12892
rect 13580 -12912 13590 -12902
rect 13330 -12962 13590 -12912
rect 13650 -12962 13660 -12902
rect 13260 -12972 13660 -12962
rect 13716 -12552 14116 -12542
rect 13716 -12612 13726 -12552
rect 13786 -12602 14046 -12552
rect 13786 -12612 13796 -12602
rect 13716 -12622 13796 -12612
rect 14036 -12612 14046 -12602
rect 14106 -12612 14116 -12552
rect 14036 -12622 14116 -12612
rect 13716 -12892 13776 -12622
rect 14046 -12632 14116 -12622
rect 13856 -12682 13886 -12662
rect 13836 -12722 13886 -12682
rect 13946 -12682 13976 -12662
rect 13946 -12722 13996 -12682
rect 13836 -12792 13996 -12722
rect 13836 -12832 13886 -12792
rect 13856 -12852 13886 -12832
rect 13946 -12832 13996 -12792
rect 13946 -12852 13976 -12832
rect 14056 -12892 14116 -12632
rect 13716 -12902 13796 -12892
rect 13716 -12962 13726 -12902
rect 13786 -12912 13796 -12902
rect 14036 -12902 14116 -12892
rect 14036 -12912 14046 -12902
rect 13786 -12962 14046 -12912
rect 14106 -12962 14116 -12902
rect 13716 -12972 14116 -12962
rect 14172 -12552 14572 -12542
rect 14172 -12612 14182 -12552
rect 14242 -12602 14502 -12552
rect 14242 -12612 14252 -12602
rect 14172 -12622 14252 -12612
rect 14492 -12612 14502 -12602
rect 14562 -12612 14572 -12552
rect 14492 -12622 14572 -12612
rect 14172 -12892 14232 -12622
rect 14502 -12632 14572 -12622
rect 14312 -12682 14342 -12662
rect 14292 -12722 14342 -12682
rect 14402 -12682 14432 -12662
rect 14402 -12722 14452 -12682
rect 14292 -12792 14452 -12722
rect 14292 -12832 14342 -12792
rect 14312 -12852 14342 -12832
rect 14402 -12832 14452 -12792
rect 14402 -12852 14432 -12832
rect 14512 -12892 14572 -12632
rect 14172 -12902 14252 -12892
rect 14172 -12962 14182 -12902
rect 14242 -12912 14252 -12902
rect 14492 -12902 14572 -12892
rect 14492 -12912 14502 -12902
rect 14242 -12962 14502 -12912
rect 14562 -12962 14572 -12902
rect 14172 -12972 14572 -12962
rect 14630 -12552 15030 -12542
rect 14630 -12612 14640 -12552
rect 14700 -12602 14960 -12552
rect 14700 -12612 14710 -12602
rect 14630 -12622 14710 -12612
rect 14950 -12612 14960 -12602
rect 15020 -12612 15030 -12552
rect 14950 -12622 15030 -12612
rect 14630 -12892 14690 -12622
rect 14960 -12632 15030 -12622
rect 14770 -12682 14800 -12662
rect 14750 -12722 14800 -12682
rect 14860 -12682 14890 -12662
rect 14860 -12722 14910 -12682
rect 14750 -12792 14910 -12722
rect 14750 -12832 14800 -12792
rect 14770 -12852 14800 -12832
rect 14860 -12832 14910 -12792
rect 14860 -12852 14890 -12832
rect 14970 -12892 15030 -12632
rect 14630 -12902 14710 -12892
rect 14630 -12962 14640 -12902
rect 14700 -12912 14710 -12902
rect 14950 -12902 15030 -12892
rect 14950 -12912 14960 -12902
rect 14700 -12962 14960 -12912
rect 15020 -12962 15030 -12902
rect 14630 -12972 15030 -12962
rect 15086 -12552 15486 -12542
rect 15086 -12612 15096 -12552
rect 15156 -12602 15416 -12552
rect 15156 -12612 15166 -12602
rect 15086 -12622 15166 -12612
rect 15406 -12612 15416 -12602
rect 15476 -12612 15486 -12552
rect 15406 -12622 15486 -12612
rect 15086 -12892 15146 -12622
rect 15416 -12632 15486 -12622
rect 15226 -12682 15256 -12662
rect 15206 -12722 15256 -12682
rect 15316 -12682 15346 -12662
rect 15316 -12722 15366 -12682
rect 15206 -12792 15366 -12722
rect 15206 -12832 15256 -12792
rect 15226 -12852 15256 -12832
rect 15316 -12832 15366 -12792
rect 15316 -12852 15346 -12832
rect 15426 -12892 15486 -12632
rect 15086 -12902 15166 -12892
rect 15086 -12962 15096 -12902
rect 15156 -12912 15166 -12902
rect 15406 -12902 15486 -12892
rect 15406 -12912 15416 -12902
rect 15156 -12962 15416 -12912
rect 15476 -12962 15486 -12902
rect 15086 -12972 15486 -12962
rect 0 -13054 400 -13044
rect 0 -13114 10 -13054
rect 70 -13104 330 -13054
rect 70 -13114 80 -13104
rect 0 -13124 80 -13114
rect 320 -13114 330 -13104
rect 390 -13114 400 -13054
rect 320 -13124 400 -13114
rect 0 -13394 60 -13124
rect 330 -13134 400 -13124
rect 140 -13184 170 -13164
rect 120 -13224 170 -13184
rect 230 -13184 260 -13164
rect 230 -13224 280 -13184
rect 120 -13294 280 -13224
rect 120 -13334 170 -13294
rect 140 -13354 170 -13334
rect 230 -13334 280 -13294
rect 230 -13354 260 -13334
rect 340 -13394 400 -13134
rect 0 -13404 80 -13394
rect 0 -13464 10 -13404
rect 70 -13414 80 -13404
rect 320 -13404 400 -13394
rect 320 -13414 330 -13404
rect 70 -13464 330 -13414
rect 390 -13464 400 -13404
rect 0 -13474 400 -13464
rect 456 -13054 856 -13044
rect 456 -13114 466 -13054
rect 526 -13104 786 -13054
rect 526 -13114 536 -13104
rect 456 -13124 536 -13114
rect 776 -13114 786 -13104
rect 846 -13114 856 -13054
rect 776 -13124 856 -13114
rect 456 -13394 516 -13124
rect 786 -13134 856 -13124
rect 596 -13184 626 -13164
rect 576 -13224 626 -13184
rect 686 -13184 716 -13164
rect 686 -13224 736 -13184
rect 576 -13294 736 -13224
rect 576 -13334 626 -13294
rect 596 -13354 626 -13334
rect 686 -13334 736 -13294
rect 686 -13354 716 -13334
rect 796 -13394 856 -13134
rect 456 -13404 536 -13394
rect 456 -13464 466 -13404
rect 526 -13414 536 -13404
rect 776 -13404 856 -13394
rect 776 -13414 786 -13404
rect 526 -13464 786 -13414
rect 846 -13464 856 -13404
rect 456 -13474 856 -13464
rect 912 -13054 1312 -13044
rect 912 -13114 922 -13054
rect 982 -13104 1242 -13054
rect 982 -13114 992 -13104
rect 912 -13124 992 -13114
rect 1232 -13114 1242 -13104
rect 1302 -13114 1312 -13054
rect 1232 -13124 1312 -13114
rect 912 -13394 972 -13124
rect 1242 -13134 1312 -13124
rect 1052 -13184 1082 -13164
rect 1032 -13224 1082 -13184
rect 1142 -13184 1172 -13164
rect 1142 -13224 1192 -13184
rect 1032 -13294 1192 -13224
rect 1032 -13334 1082 -13294
rect 1052 -13354 1082 -13334
rect 1142 -13334 1192 -13294
rect 1142 -13354 1172 -13334
rect 1252 -13394 1312 -13134
rect 912 -13404 992 -13394
rect 912 -13464 922 -13404
rect 982 -13414 992 -13404
rect 1232 -13404 1312 -13394
rect 1232 -13414 1242 -13404
rect 982 -13464 1242 -13414
rect 1302 -13464 1312 -13404
rect 912 -13474 1312 -13464
rect 1370 -13054 1770 -13044
rect 1370 -13114 1380 -13054
rect 1440 -13104 1700 -13054
rect 1440 -13114 1450 -13104
rect 1370 -13124 1450 -13114
rect 1690 -13114 1700 -13104
rect 1760 -13114 1770 -13054
rect 1690 -13124 1770 -13114
rect 1370 -13394 1430 -13124
rect 1700 -13134 1770 -13124
rect 1510 -13184 1540 -13164
rect 1490 -13224 1540 -13184
rect 1600 -13184 1630 -13164
rect 1600 -13224 1650 -13184
rect 1490 -13294 1650 -13224
rect 1490 -13334 1540 -13294
rect 1510 -13354 1540 -13334
rect 1600 -13334 1650 -13294
rect 1600 -13354 1630 -13334
rect 1710 -13394 1770 -13134
rect 1370 -13404 1450 -13394
rect 1370 -13464 1380 -13404
rect 1440 -13414 1450 -13404
rect 1690 -13404 1770 -13394
rect 1690 -13414 1700 -13404
rect 1440 -13464 1700 -13414
rect 1760 -13464 1770 -13404
rect 1370 -13474 1770 -13464
rect 1826 -13054 2226 -13044
rect 1826 -13114 1836 -13054
rect 1896 -13104 2156 -13054
rect 1896 -13114 1906 -13104
rect 1826 -13124 1906 -13114
rect 2146 -13114 2156 -13104
rect 2216 -13114 2226 -13054
rect 2146 -13124 2226 -13114
rect 1826 -13394 1886 -13124
rect 2156 -13134 2226 -13124
rect 1966 -13184 1996 -13164
rect 1946 -13224 1996 -13184
rect 2056 -13184 2086 -13164
rect 2056 -13224 2106 -13184
rect 1946 -13294 2106 -13224
rect 1946 -13334 1996 -13294
rect 1966 -13354 1996 -13334
rect 2056 -13334 2106 -13294
rect 2056 -13354 2086 -13334
rect 2166 -13394 2226 -13134
rect 1826 -13404 1906 -13394
rect 1826 -13464 1836 -13404
rect 1896 -13414 1906 -13404
rect 2146 -13404 2226 -13394
rect 2146 -13414 2156 -13404
rect 1896 -13464 2156 -13414
rect 2216 -13464 2226 -13404
rect 1826 -13474 2226 -13464
rect 2282 -13054 2682 -13044
rect 2282 -13114 2292 -13054
rect 2352 -13104 2612 -13054
rect 2352 -13114 2362 -13104
rect 2282 -13124 2362 -13114
rect 2602 -13114 2612 -13104
rect 2672 -13114 2682 -13054
rect 2602 -13124 2682 -13114
rect 2282 -13394 2342 -13124
rect 2612 -13134 2682 -13124
rect 2422 -13184 2452 -13164
rect 2402 -13224 2452 -13184
rect 2512 -13184 2542 -13164
rect 2512 -13224 2562 -13184
rect 2402 -13294 2562 -13224
rect 2402 -13334 2452 -13294
rect 2422 -13354 2452 -13334
rect 2512 -13334 2562 -13294
rect 2512 -13354 2542 -13334
rect 2622 -13394 2682 -13134
rect 2282 -13404 2362 -13394
rect 2282 -13464 2292 -13404
rect 2352 -13414 2362 -13404
rect 2602 -13404 2682 -13394
rect 2602 -13414 2612 -13404
rect 2352 -13464 2612 -13414
rect 2672 -13464 2682 -13404
rect 2282 -13474 2682 -13464
rect 2740 -13054 3140 -13044
rect 2740 -13114 2750 -13054
rect 2810 -13104 3070 -13054
rect 2810 -13114 2820 -13104
rect 2740 -13124 2820 -13114
rect 3060 -13114 3070 -13104
rect 3130 -13114 3140 -13054
rect 3060 -13124 3140 -13114
rect 2740 -13394 2800 -13124
rect 3070 -13134 3140 -13124
rect 2880 -13184 2910 -13164
rect 2860 -13224 2910 -13184
rect 2970 -13184 3000 -13164
rect 2970 -13224 3020 -13184
rect 2860 -13294 3020 -13224
rect 2860 -13334 2910 -13294
rect 2880 -13354 2910 -13334
rect 2970 -13334 3020 -13294
rect 2970 -13354 3000 -13334
rect 3080 -13394 3140 -13134
rect 2740 -13404 2820 -13394
rect 2740 -13464 2750 -13404
rect 2810 -13414 2820 -13404
rect 3060 -13404 3140 -13394
rect 3060 -13414 3070 -13404
rect 2810 -13464 3070 -13414
rect 3130 -13464 3140 -13404
rect 2740 -13474 3140 -13464
rect 3196 -13054 3596 -13044
rect 3196 -13114 3206 -13054
rect 3266 -13104 3526 -13054
rect 3266 -13114 3276 -13104
rect 3196 -13124 3276 -13114
rect 3516 -13114 3526 -13104
rect 3586 -13114 3596 -13054
rect 3516 -13124 3596 -13114
rect 3196 -13394 3256 -13124
rect 3526 -13134 3596 -13124
rect 3336 -13184 3366 -13164
rect 3316 -13224 3366 -13184
rect 3426 -13184 3456 -13164
rect 3426 -13224 3476 -13184
rect 3316 -13294 3476 -13224
rect 3316 -13334 3366 -13294
rect 3336 -13354 3366 -13334
rect 3426 -13334 3476 -13294
rect 3426 -13354 3456 -13334
rect 3536 -13394 3596 -13134
rect 3196 -13404 3276 -13394
rect 3196 -13464 3206 -13404
rect 3266 -13414 3276 -13404
rect 3516 -13404 3596 -13394
rect 3516 -13414 3526 -13404
rect 3266 -13464 3526 -13414
rect 3586 -13464 3596 -13404
rect 3196 -13474 3596 -13464
rect 3652 -13054 4052 -13044
rect 3652 -13114 3662 -13054
rect 3722 -13104 3982 -13054
rect 3722 -13114 3732 -13104
rect 3652 -13124 3732 -13114
rect 3972 -13114 3982 -13104
rect 4042 -13114 4052 -13054
rect 3972 -13124 4052 -13114
rect 3652 -13394 3712 -13124
rect 3982 -13134 4052 -13124
rect 3792 -13184 3822 -13164
rect 3772 -13224 3822 -13184
rect 3882 -13184 3912 -13164
rect 3882 -13224 3932 -13184
rect 3772 -13294 3932 -13224
rect 3772 -13334 3822 -13294
rect 3792 -13354 3822 -13334
rect 3882 -13334 3932 -13294
rect 3882 -13354 3912 -13334
rect 3992 -13394 4052 -13134
rect 3652 -13404 3732 -13394
rect 3652 -13464 3662 -13404
rect 3722 -13414 3732 -13404
rect 3972 -13404 4052 -13394
rect 3972 -13414 3982 -13404
rect 3722 -13464 3982 -13414
rect 4042 -13464 4052 -13404
rect 3652 -13474 4052 -13464
rect 4110 -13054 4510 -13044
rect 4110 -13114 4120 -13054
rect 4180 -13104 4440 -13054
rect 4180 -13114 4190 -13104
rect 4110 -13124 4190 -13114
rect 4430 -13114 4440 -13104
rect 4500 -13114 4510 -13054
rect 4430 -13124 4510 -13114
rect 4110 -13394 4170 -13124
rect 4440 -13134 4510 -13124
rect 4250 -13184 4280 -13164
rect 4230 -13224 4280 -13184
rect 4340 -13184 4370 -13164
rect 4340 -13224 4390 -13184
rect 4230 -13294 4390 -13224
rect 4230 -13334 4280 -13294
rect 4250 -13354 4280 -13334
rect 4340 -13334 4390 -13294
rect 4340 -13354 4370 -13334
rect 4450 -13394 4510 -13134
rect 4110 -13404 4190 -13394
rect 4110 -13464 4120 -13404
rect 4180 -13414 4190 -13404
rect 4430 -13404 4510 -13394
rect 4430 -13414 4440 -13404
rect 4180 -13464 4440 -13414
rect 4500 -13464 4510 -13404
rect 4110 -13474 4510 -13464
rect 4566 -13054 4966 -13044
rect 4566 -13114 4576 -13054
rect 4636 -13104 4896 -13054
rect 4636 -13114 4646 -13104
rect 4566 -13124 4646 -13114
rect 4886 -13114 4896 -13104
rect 4956 -13114 4966 -13054
rect 4886 -13124 4966 -13114
rect 4566 -13394 4626 -13124
rect 4896 -13134 4966 -13124
rect 4706 -13184 4736 -13164
rect 4686 -13224 4736 -13184
rect 4796 -13184 4826 -13164
rect 4796 -13224 4846 -13184
rect 4686 -13294 4846 -13224
rect 4686 -13334 4736 -13294
rect 4706 -13354 4736 -13334
rect 4796 -13334 4846 -13294
rect 4796 -13354 4826 -13334
rect 4906 -13394 4966 -13134
rect 4566 -13404 4646 -13394
rect 4566 -13464 4576 -13404
rect 4636 -13414 4646 -13404
rect 4886 -13404 4966 -13394
rect 4886 -13414 4896 -13404
rect 4636 -13464 4896 -13414
rect 4956 -13464 4966 -13404
rect 4566 -13474 4966 -13464
rect 5022 -13054 5422 -13044
rect 5022 -13114 5032 -13054
rect 5092 -13104 5352 -13054
rect 5092 -13114 5102 -13104
rect 5022 -13124 5102 -13114
rect 5342 -13114 5352 -13104
rect 5412 -13114 5422 -13054
rect 5342 -13124 5422 -13114
rect 5022 -13394 5082 -13124
rect 5352 -13134 5422 -13124
rect 5162 -13184 5192 -13164
rect 5142 -13224 5192 -13184
rect 5252 -13184 5282 -13164
rect 5252 -13224 5302 -13184
rect 5142 -13294 5302 -13224
rect 5142 -13334 5192 -13294
rect 5162 -13354 5192 -13334
rect 5252 -13334 5302 -13294
rect 5252 -13354 5282 -13334
rect 5362 -13394 5422 -13134
rect 5022 -13404 5102 -13394
rect 5022 -13464 5032 -13404
rect 5092 -13414 5102 -13404
rect 5342 -13404 5422 -13394
rect 5342 -13414 5352 -13404
rect 5092 -13464 5352 -13414
rect 5412 -13464 5422 -13404
rect 5022 -13474 5422 -13464
rect 5480 -13054 5880 -13044
rect 5480 -13114 5490 -13054
rect 5550 -13104 5810 -13054
rect 5550 -13114 5560 -13104
rect 5480 -13124 5560 -13114
rect 5800 -13114 5810 -13104
rect 5870 -13114 5880 -13054
rect 5800 -13124 5880 -13114
rect 5480 -13394 5540 -13124
rect 5810 -13134 5880 -13124
rect 5620 -13184 5650 -13164
rect 5600 -13224 5650 -13184
rect 5710 -13184 5740 -13164
rect 5710 -13224 5760 -13184
rect 5600 -13294 5760 -13224
rect 5600 -13334 5650 -13294
rect 5620 -13354 5650 -13334
rect 5710 -13334 5760 -13294
rect 5710 -13354 5740 -13334
rect 5820 -13394 5880 -13134
rect 5480 -13404 5560 -13394
rect 5480 -13464 5490 -13404
rect 5550 -13414 5560 -13404
rect 5800 -13404 5880 -13394
rect 5800 -13414 5810 -13404
rect 5550 -13464 5810 -13414
rect 5870 -13464 5880 -13404
rect 5480 -13474 5880 -13464
rect 5936 -13054 6336 -13044
rect 5936 -13114 5946 -13054
rect 6006 -13104 6266 -13054
rect 6006 -13114 6016 -13104
rect 5936 -13124 6016 -13114
rect 6256 -13114 6266 -13104
rect 6326 -13114 6336 -13054
rect 6256 -13124 6336 -13114
rect 5936 -13394 5996 -13124
rect 6266 -13134 6336 -13124
rect 6076 -13184 6106 -13164
rect 6056 -13224 6106 -13184
rect 6166 -13184 6196 -13164
rect 6166 -13224 6216 -13184
rect 6056 -13294 6216 -13224
rect 6056 -13334 6106 -13294
rect 6076 -13354 6106 -13334
rect 6166 -13334 6216 -13294
rect 6166 -13354 6196 -13334
rect 6276 -13394 6336 -13134
rect 5936 -13404 6016 -13394
rect 5936 -13464 5946 -13404
rect 6006 -13414 6016 -13404
rect 6256 -13404 6336 -13394
rect 6256 -13414 6266 -13404
rect 6006 -13464 6266 -13414
rect 6326 -13464 6336 -13404
rect 5936 -13474 6336 -13464
rect 6392 -13054 6792 -13044
rect 6392 -13114 6402 -13054
rect 6462 -13104 6722 -13054
rect 6462 -13114 6472 -13104
rect 6392 -13124 6472 -13114
rect 6712 -13114 6722 -13104
rect 6782 -13114 6792 -13054
rect 6712 -13124 6792 -13114
rect 6392 -13394 6452 -13124
rect 6722 -13134 6792 -13124
rect 6532 -13184 6562 -13164
rect 6512 -13224 6562 -13184
rect 6622 -13184 6652 -13164
rect 6622 -13224 6672 -13184
rect 6512 -13294 6672 -13224
rect 6512 -13334 6562 -13294
rect 6532 -13354 6562 -13334
rect 6622 -13334 6672 -13294
rect 6622 -13354 6652 -13334
rect 6732 -13394 6792 -13134
rect 6392 -13404 6472 -13394
rect 6392 -13464 6402 -13404
rect 6462 -13414 6472 -13404
rect 6712 -13404 6792 -13394
rect 6712 -13414 6722 -13404
rect 6462 -13464 6722 -13414
rect 6782 -13464 6792 -13404
rect 6392 -13474 6792 -13464
rect 6850 -13054 7250 -13044
rect 6850 -13114 6860 -13054
rect 6920 -13104 7180 -13054
rect 6920 -13114 6930 -13104
rect 6850 -13124 6930 -13114
rect 7170 -13114 7180 -13104
rect 7240 -13114 7250 -13054
rect 7170 -13124 7250 -13114
rect 6850 -13394 6910 -13124
rect 7180 -13134 7250 -13124
rect 6990 -13184 7020 -13164
rect 6970 -13224 7020 -13184
rect 7080 -13184 7110 -13164
rect 7080 -13224 7130 -13184
rect 6970 -13294 7130 -13224
rect 6970 -13334 7020 -13294
rect 6990 -13354 7020 -13334
rect 7080 -13334 7130 -13294
rect 7080 -13354 7110 -13334
rect 7190 -13394 7250 -13134
rect 6850 -13404 6930 -13394
rect 6850 -13464 6860 -13404
rect 6920 -13414 6930 -13404
rect 7170 -13404 7250 -13394
rect 7170 -13414 7180 -13404
rect 6920 -13464 7180 -13414
rect 7240 -13464 7250 -13404
rect 6850 -13474 7250 -13464
rect 7306 -13054 7706 -13044
rect 7306 -13114 7316 -13054
rect 7376 -13104 7636 -13054
rect 7376 -13114 7386 -13104
rect 7306 -13124 7386 -13114
rect 7626 -13114 7636 -13104
rect 7696 -13114 7706 -13054
rect 7626 -13124 7706 -13114
rect 7306 -13394 7366 -13124
rect 7636 -13134 7706 -13124
rect 7446 -13184 7476 -13164
rect 7426 -13224 7476 -13184
rect 7536 -13184 7566 -13164
rect 7536 -13224 7586 -13184
rect 7426 -13294 7586 -13224
rect 7426 -13334 7476 -13294
rect 7446 -13354 7476 -13334
rect 7536 -13334 7586 -13294
rect 7536 -13354 7566 -13334
rect 7646 -13394 7706 -13134
rect 7306 -13404 7386 -13394
rect 7306 -13464 7316 -13404
rect 7376 -13414 7386 -13404
rect 7626 -13404 7706 -13394
rect 7626 -13414 7636 -13404
rect 7376 -13464 7636 -13414
rect 7696 -13464 7706 -13404
rect 7306 -13474 7706 -13464
rect 7762 -13054 8162 -13044
rect 7762 -13114 7772 -13054
rect 7832 -13104 8092 -13054
rect 7832 -13114 7842 -13104
rect 7762 -13124 7842 -13114
rect 8082 -13114 8092 -13104
rect 8152 -13114 8162 -13054
rect 8082 -13124 8162 -13114
rect 7762 -13394 7822 -13124
rect 8092 -13134 8162 -13124
rect 7902 -13184 7932 -13164
rect 7882 -13224 7932 -13184
rect 7992 -13184 8022 -13164
rect 7992 -13224 8042 -13184
rect 7882 -13294 8042 -13224
rect 7882 -13334 7932 -13294
rect 7902 -13354 7932 -13334
rect 7992 -13334 8042 -13294
rect 7992 -13354 8022 -13334
rect 8102 -13394 8162 -13134
rect 7762 -13404 7842 -13394
rect 7762 -13464 7772 -13404
rect 7832 -13414 7842 -13404
rect 8082 -13404 8162 -13394
rect 8082 -13414 8092 -13404
rect 7832 -13464 8092 -13414
rect 8152 -13464 8162 -13404
rect 7762 -13474 8162 -13464
rect 8236 -13054 8636 -13044
rect 8236 -13114 8246 -13054
rect 8306 -13104 8566 -13054
rect 8306 -13114 8316 -13104
rect 8236 -13124 8316 -13114
rect 8556 -13114 8566 -13104
rect 8626 -13114 8636 -13054
rect 8556 -13124 8636 -13114
rect 8236 -13394 8296 -13124
rect 8566 -13134 8636 -13124
rect 8376 -13184 8406 -13164
rect 8356 -13224 8406 -13184
rect 8466 -13184 8496 -13164
rect 8466 -13224 8516 -13184
rect 8356 -13294 8516 -13224
rect 8356 -13334 8406 -13294
rect 8376 -13354 8406 -13334
rect 8466 -13334 8516 -13294
rect 8466 -13354 8496 -13334
rect 8576 -13394 8636 -13134
rect 8236 -13404 8316 -13394
rect 8236 -13464 8246 -13404
rect 8306 -13414 8316 -13404
rect 8556 -13404 8636 -13394
rect 8556 -13414 8566 -13404
rect 8306 -13464 8566 -13414
rect 8626 -13464 8636 -13404
rect 8236 -13474 8636 -13464
rect 8692 -13054 9092 -13044
rect 8692 -13114 8702 -13054
rect 8762 -13104 9022 -13054
rect 8762 -13114 8772 -13104
rect 8692 -13124 8772 -13114
rect 9012 -13114 9022 -13104
rect 9082 -13114 9092 -13054
rect 9012 -13124 9092 -13114
rect 8692 -13394 8752 -13124
rect 9022 -13134 9092 -13124
rect 8832 -13184 8862 -13164
rect 8812 -13224 8862 -13184
rect 8922 -13184 8952 -13164
rect 8922 -13224 8972 -13184
rect 8812 -13294 8972 -13224
rect 8812 -13334 8862 -13294
rect 8832 -13354 8862 -13334
rect 8922 -13334 8972 -13294
rect 8922 -13354 8952 -13334
rect 9032 -13394 9092 -13134
rect 8692 -13404 8772 -13394
rect 8692 -13464 8702 -13404
rect 8762 -13414 8772 -13404
rect 9012 -13404 9092 -13394
rect 9012 -13414 9022 -13404
rect 8762 -13464 9022 -13414
rect 9082 -13464 9092 -13404
rect 8692 -13474 9092 -13464
rect 9150 -13054 9550 -13044
rect 9150 -13114 9160 -13054
rect 9220 -13104 9480 -13054
rect 9220 -13114 9230 -13104
rect 9150 -13124 9230 -13114
rect 9470 -13114 9480 -13104
rect 9540 -13114 9550 -13054
rect 9470 -13124 9550 -13114
rect 9150 -13394 9210 -13124
rect 9480 -13134 9550 -13124
rect 9290 -13184 9320 -13164
rect 9270 -13224 9320 -13184
rect 9380 -13184 9410 -13164
rect 9380 -13224 9430 -13184
rect 9270 -13294 9430 -13224
rect 9270 -13334 9320 -13294
rect 9290 -13354 9320 -13334
rect 9380 -13334 9430 -13294
rect 9380 -13354 9410 -13334
rect 9490 -13394 9550 -13134
rect 9150 -13404 9230 -13394
rect 9150 -13464 9160 -13404
rect 9220 -13414 9230 -13404
rect 9470 -13404 9550 -13394
rect 9470 -13414 9480 -13404
rect 9220 -13464 9480 -13414
rect 9540 -13464 9550 -13404
rect 9150 -13474 9550 -13464
rect 9606 -13054 10006 -13044
rect 9606 -13114 9616 -13054
rect 9676 -13104 9936 -13054
rect 9676 -13114 9686 -13104
rect 9606 -13124 9686 -13114
rect 9926 -13114 9936 -13104
rect 9996 -13114 10006 -13054
rect 9926 -13124 10006 -13114
rect 9606 -13394 9666 -13124
rect 9936 -13134 10006 -13124
rect 9746 -13184 9776 -13164
rect 9726 -13224 9776 -13184
rect 9836 -13184 9866 -13164
rect 9836 -13224 9886 -13184
rect 9726 -13294 9886 -13224
rect 9726 -13334 9776 -13294
rect 9746 -13354 9776 -13334
rect 9836 -13334 9886 -13294
rect 9836 -13354 9866 -13334
rect 9946 -13394 10006 -13134
rect 9606 -13404 9686 -13394
rect 9606 -13464 9616 -13404
rect 9676 -13414 9686 -13404
rect 9926 -13404 10006 -13394
rect 9926 -13414 9936 -13404
rect 9676 -13464 9936 -13414
rect 9996 -13464 10006 -13404
rect 9606 -13474 10006 -13464
rect 10062 -13054 10462 -13044
rect 10062 -13114 10072 -13054
rect 10132 -13104 10392 -13054
rect 10132 -13114 10142 -13104
rect 10062 -13124 10142 -13114
rect 10382 -13114 10392 -13104
rect 10452 -13114 10462 -13054
rect 10382 -13124 10462 -13114
rect 10062 -13394 10122 -13124
rect 10392 -13134 10462 -13124
rect 10202 -13184 10232 -13164
rect 10182 -13224 10232 -13184
rect 10292 -13184 10322 -13164
rect 10292 -13224 10342 -13184
rect 10182 -13294 10342 -13224
rect 10182 -13334 10232 -13294
rect 10202 -13354 10232 -13334
rect 10292 -13334 10342 -13294
rect 10292 -13354 10322 -13334
rect 10402 -13394 10462 -13134
rect 10062 -13404 10142 -13394
rect 10062 -13464 10072 -13404
rect 10132 -13414 10142 -13404
rect 10382 -13404 10462 -13394
rect 10382 -13414 10392 -13404
rect 10132 -13464 10392 -13414
rect 10452 -13464 10462 -13404
rect 10062 -13474 10462 -13464
rect 10520 -13054 10920 -13044
rect 10520 -13114 10530 -13054
rect 10590 -13104 10850 -13054
rect 10590 -13114 10600 -13104
rect 10520 -13124 10600 -13114
rect 10840 -13114 10850 -13104
rect 10910 -13114 10920 -13054
rect 10840 -13124 10920 -13114
rect 10520 -13394 10580 -13124
rect 10850 -13134 10920 -13124
rect 10660 -13184 10690 -13164
rect 10640 -13224 10690 -13184
rect 10750 -13184 10780 -13164
rect 10750 -13224 10800 -13184
rect 10640 -13294 10800 -13224
rect 10640 -13334 10690 -13294
rect 10660 -13354 10690 -13334
rect 10750 -13334 10800 -13294
rect 10750 -13354 10780 -13334
rect 10860 -13394 10920 -13134
rect 10520 -13404 10600 -13394
rect 10520 -13464 10530 -13404
rect 10590 -13414 10600 -13404
rect 10840 -13404 10920 -13394
rect 10840 -13414 10850 -13404
rect 10590 -13464 10850 -13414
rect 10910 -13464 10920 -13404
rect 10520 -13474 10920 -13464
rect 10976 -13054 11376 -13044
rect 10976 -13114 10986 -13054
rect 11046 -13104 11306 -13054
rect 11046 -13114 11056 -13104
rect 10976 -13124 11056 -13114
rect 11296 -13114 11306 -13104
rect 11366 -13114 11376 -13054
rect 11296 -13124 11376 -13114
rect 10976 -13394 11036 -13124
rect 11306 -13134 11376 -13124
rect 11116 -13184 11146 -13164
rect 11096 -13224 11146 -13184
rect 11206 -13184 11236 -13164
rect 11206 -13224 11256 -13184
rect 11096 -13294 11256 -13224
rect 11096 -13334 11146 -13294
rect 11116 -13354 11146 -13334
rect 11206 -13334 11256 -13294
rect 11206 -13354 11236 -13334
rect 11316 -13394 11376 -13134
rect 10976 -13404 11056 -13394
rect 10976 -13464 10986 -13404
rect 11046 -13414 11056 -13404
rect 11296 -13404 11376 -13394
rect 11296 -13414 11306 -13404
rect 11046 -13464 11306 -13414
rect 11366 -13464 11376 -13404
rect 10976 -13474 11376 -13464
rect 11432 -13054 11832 -13044
rect 11432 -13114 11442 -13054
rect 11502 -13104 11762 -13054
rect 11502 -13114 11512 -13104
rect 11432 -13124 11512 -13114
rect 11752 -13114 11762 -13104
rect 11822 -13114 11832 -13054
rect 11752 -13124 11832 -13114
rect 11432 -13394 11492 -13124
rect 11762 -13134 11832 -13124
rect 11572 -13184 11602 -13164
rect 11552 -13224 11602 -13184
rect 11662 -13184 11692 -13164
rect 11662 -13224 11712 -13184
rect 11552 -13294 11712 -13224
rect 11552 -13334 11602 -13294
rect 11572 -13354 11602 -13334
rect 11662 -13334 11712 -13294
rect 11662 -13354 11692 -13334
rect 11772 -13394 11832 -13134
rect 11432 -13404 11512 -13394
rect 11432 -13464 11442 -13404
rect 11502 -13414 11512 -13404
rect 11752 -13404 11832 -13394
rect 11752 -13414 11762 -13404
rect 11502 -13464 11762 -13414
rect 11822 -13464 11832 -13404
rect 11432 -13474 11832 -13464
rect 11890 -13054 12290 -13044
rect 11890 -13114 11900 -13054
rect 11960 -13104 12220 -13054
rect 11960 -13114 11970 -13104
rect 11890 -13124 11970 -13114
rect 12210 -13114 12220 -13104
rect 12280 -13114 12290 -13054
rect 12210 -13124 12290 -13114
rect 11890 -13394 11950 -13124
rect 12220 -13134 12290 -13124
rect 12030 -13184 12060 -13164
rect 12010 -13224 12060 -13184
rect 12120 -13184 12150 -13164
rect 12120 -13224 12170 -13184
rect 12010 -13294 12170 -13224
rect 12010 -13334 12060 -13294
rect 12030 -13354 12060 -13334
rect 12120 -13334 12170 -13294
rect 12120 -13354 12150 -13334
rect 12230 -13394 12290 -13134
rect 11890 -13404 11970 -13394
rect 11890 -13464 11900 -13404
rect 11960 -13414 11970 -13404
rect 12210 -13404 12290 -13394
rect 12210 -13414 12220 -13404
rect 11960 -13464 12220 -13414
rect 12280 -13464 12290 -13404
rect 11890 -13474 12290 -13464
rect 12346 -13054 12746 -13044
rect 12346 -13114 12356 -13054
rect 12416 -13104 12676 -13054
rect 12416 -13114 12426 -13104
rect 12346 -13124 12426 -13114
rect 12666 -13114 12676 -13104
rect 12736 -13114 12746 -13054
rect 12666 -13124 12746 -13114
rect 12346 -13394 12406 -13124
rect 12676 -13134 12746 -13124
rect 12486 -13184 12516 -13164
rect 12466 -13224 12516 -13184
rect 12576 -13184 12606 -13164
rect 12576 -13224 12626 -13184
rect 12466 -13294 12626 -13224
rect 12466 -13334 12516 -13294
rect 12486 -13354 12516 -13334
rect 12576 -13334 12626 -13294
rect 12576 -13354 12606 -13334
rect 12686 -13394 12746 -13134
rect 12346 -13404 12426 -13394
rect 12346 -13464 12356 -13404
rect 12416 -13414 12426 -13404
rect 12666 -13404 12746 -13394
rect 12666 -13414 12676 -13404
rect 12416 -13464 12676 -13414
rect 12736 -13464 12746 -13404
rect 12346 -13474 12746 -13464
rect 12802 -13054 13202 -13044
rect 12802 -13114 12812 -13054
rect 12872 -13104 13132 -13054
rect 12872 -13114 12882 -13104
rect 12802 -13124 12882 -13114
rect 13122 -13114 13132 -13104
rect 13192 -13114 13202 -13054
rect 13122 -13124 13202 -13114
rect 12802 -13394 12862 -13124
rect 13132 -13134 13202 -13124
rect 12942 -13184 12972 -13164
rect 12922 -13224 12972 -13184
rect 13032 -13184 13062 -13164
rect 13032 -13224 13082 -13184
rect 12922 -13294 13082 -13224
rect 12922 -13334 12972 -13294
rect 12942 -13354 12972 -13334
rect 13032 -13334 13082 -13294
rect 13032 -13354 13062 -13334
rect 13142 -13394 13202 -13134
rect 12802 -13404 12882 -13394
rect 12802 -13464 12812 -13404
rect 12872 -13414 12882 -13404
rect 13122 -13404 13202 -13394
rect 13122 -13414 13132 -13404
rect 12872 -13464 13132 -13414
rect 13192 -13464 13202 -13404
rect 12802 -13474 13202 -13464
rect 13260 -13054 13660 -13044
rect 13260 -13114 13270 -13054
rect 13330 -13104 13590 -13054
rect 13330 -13114 13340 -13104
rect 13260 -13124 13340 -13114
rect 13580 -13114 13590 -13104
rect 13650 -13114 13660 -13054
rect 13580 -13124 13660 -13114
rect 13260 -13394 13320 -13124
rect 13590 -13134 13660 -13124
rect 13400 -13184 13430 -13164
rect 13380 -13224 13430 -13184
rect 13490 -13184 13520 -13164
rect 13490 -13224 13540 -13184
rect 13380 -13294 13540 -13224
rect 13380 -13334 13430 -13294
rect 13400 -13354 13430 -13334
rect 13490 -13334 13540 -13294
rect 13490 -13354 13520 -13334
rect 13600 -13394 13660 -13134
rect 13260 -13404 13340 -13394
rect 13260 -13464 13270 -13404
rect 13330 -13414 13340 -13404
rect 13580 -13404 13660 -13394
rect 13580 -13414 13590 -13404
rect 13330 -13464 13590 -13414
rect 13650 -13464 13660 -13404
rect 13260 -13474 13660 -13464
rect 13716 -13054 14116 -13044
rect 13716 -13114 13726 -13054
rect 13786 -13104 14046 -13054
rect 13786 -13114 13796 -13104
rect 13716 -13124 13796 -13114
rect 14036 -13114 14046 -13104
rect 14106 -13114 14116 -13054
rect 14036 -13124 14116 -13114
rect 13716 -13394 13776 -13124
rect 14046 -13134 14116 -13124
rect 13856 -13184 13886 -13164
rect 13836 -13224 13886 -13184
rect 13946 -13184 13976 -13164
rect 13946 -13224 13996 -13184
rect 13836 -13294 13996 -13224
rect 13836 -13334 13886 -13294
rect 13856 -13354 13886 -13334
rect 13946 -13334 13996 -13294
rect 13946 -13354 13976 -13334
rect 14056 -13394 14116 -13134
rect 13716 -13404 13796 -13394
rect 13716 -13464 13726 -13404
rect 13786 -13414 13796 -13404
rect 14036 -13404 14116 -13394
rect 14036 -13414 14046 -13404
rect 13786 -13464 14046 -13414
rect 14106 -13464 14116 -13404
rect 13716 -13474 14116 -13464
rect 14172 -13054 14572 -13044
rect 14172 -13114 14182 -13054
rect 14242 -13104 14502 -13054
rect 14242 -13114 14252 -13104
rect 14172 -13124 14252 -13114
rect 14492 -13114 14502 -13104
rect 14562 -13114 14572 -13054
rect 14492 -13124 14572 -13114
rect 14172 -13394 14232 -13124
rect 14502 -13134 14572 -13124
rect 14312 -13184 14342 -13164
rect 14292 -13224 14342 -13184
rect 14402 -13184 14432 -13164
rect 14402 -13224 14452 -13184
rect 14292 -13294 14452 -13224
rect 14292 -13334 14342 -13294
rect 14312 -13354 14342 -13334
rect 14402 -13334 14452 -13294
rect 14402 -13354 14432 -13334
rect 14512 -13394 14572 -13134
rect 14172 -13404 14252 -13394
rect 14172 -13464 14182 -13404
rect 14242 -13414 14252 -13404
rect 14492 -13404 14572 -13394
rect 14492 -13414 14502 -13404
rect 14242 -13464 14502 -13414
rect 14562 -13464 14572 -13404
rect 14172 -13474 14572 -13464
rect 14630 -13054 15030 -13044
rect 14630 -13114 14640 -13054
rect 14700 -13104 14960 -13054
rect 14700 -13114 14710 -13104
rect 14630 -13124 14710 -13114
rect 14950 -13114 14960 -13104
rect 15020 -13114 15030 -13054
rect 14950 -13124 15030 -13114
rect 14630 -13394 14690 -13124
rect 14960 -13134 15030 -13124
rect 14770 -13184 14800 -13164
rect 14750 -13224 14800 -13184
rect 14860 -13184 14890 -13164
rect 14860 -13224 14910 -13184
rect 14750 -13294 14910 -13224
rect 14750 -13334 14800 -13294
rect 14770 -13354 14800 -13334
rect 14860 -13334 14910 -13294
rect 14860 -13354 14890 -13334
rect 14970 -13394 15030 -13134
rect 14630 -13404 14710 -13394
rect 14630 -13464 14640 -13404
rect 14700 -13414 14710 -13404
rect 14950 -13404 15030 -13394
rect 14950 -13414 14960 -13404
rect 14700 -13464 14960 -13414
rect 15020 -13464 15030 -13404
rect 14630 -13474 15030 -13464
rect 15086 -13054 15486 -13044
rect 15086 -13114 15096 -13054
rect 15156 -13104 15416 -13054
rect 15156 -13114 15166 -13104
rect 15086 -13124 15166 -13114
rect 15406 -13114 15416 -13104
rect 15476 -13114 15486 -13054
rect 15406 -13124 15486 -13114
rect 15086 -13394 15146 -13124
rect 15416 -13134 15486 -13124
rect 15226 -13184 15256 -13164
rect 15206 -13224 15256 -13184
rect 15316 -13184 15346 -13164
rect 15316 -13224 15366 -13184
rect 15206 -13294 15366 -13224
rect 15206 -13334 15256 -13294
rect 15226 -13354 15256 -13334
rect 15316 -13334 15366 -13294
rect 15316 -13354 15346 -13334
rect 15426 -13394 15486 -13134
rect 15086 -13404 15166 -13394
rect 15086 -13464 15096 -13404
rect 15156 -13414 15166 -13404
rect 15406 -13404 15486 -13394
rect 15406 -13414 15416 -13404
rect 15156 -13464 15416 -13414
rect 15476 -13464 15486 -13404
rect 15086 -13474 15486 -13464
rect 0 -13546 400 -13536
rect 0 -13606 10 -13546
rect 70 -13596 330 -13546
rect 70 -13606 80 -13596
rect 0 -13616 80 -13606
rect 320 -13606 330 -13596
rect 390 -13606 400 -13546
rect 320 -13616 400 -13606
rect 0 -13886 60 -13616
rect 330 -13626 400 -13616
rect 140 -13676 170 -13656
rect 120 -13716 170 -13676
rect 230 -13676 260 -13656
rect 230 -13716 280 -13676
rect 120 -13786 280 -13716
rect 120 -13826 170 -13786
rect 140 -13846 170 -13826
rect 230 -13826 280 -13786
rect 230 -13846 260 -13826
rect 340 -13886 400 -13626
rect 0 -13896 80 -13886
rect 0 -13956 10 -13896
rect 70 -13906 80 -13896
rect 320 -13896 400 -13886
rect 320 -13906 330 -13896
rect 70 -13956 330 -13906
rect 390 -13956 400 -13896
rect 0 -13966 400 -13956
rect 456 -13546 856 -13536
rect 456 -13606 466 -13546
rect 526 -13596 786 -13546
rect 526 -13606 536 -13596
rect 456 -13616 536 -13606
rect 776 -13606 786 -13596
rect 846 -13606 856 -13546
rect 776 -13616 856 -13606
rect 456 -13886 516 -13616
rect 786 -13626 856 -13616
rect 596 -13676 626 -13656
rect 576 -13716 626 -13676
rect 686 -13676 716 -13656
rect 686 -13716 736 -13676
rect 576 -13786 736 -13716
rect 576 -13826 626 -13786
rect 596 -13846 626 -13826
rect 686 -13826 736 -13786
rect 686 -13846 716 -13826
rect 796 -13886 856 -13626
rect 456 -13896 536 -13886
rect 456 -13956 466 -13896
rect 526 -13906 536 -13896
rect 776 -13896 856 -13886
rect 776 -13906 786 -13896
rect 526 -13956 786 -13906
rect 846 -13956 856 -13896
rect 456 -13966 856 -13956
rect 912 -13546 1312 -13536
rect 912 -13606 922 -13546
rect 982 -13596 1242 -13546
rect 982 -13606 992 -13596
rect 912 -13616 992 -13606
rect 1232 -13606 1242 -13596
rect 1302 -13606 1312 -13546
rect 1232 -13616 1312 -13606
rect 912 -13886 972 -13616
rect 1242 -13626 1312 -13616
rect 1052 -13676 1082 -13656
rect 1032 -13716 1082 -13676
rect 1142 -13676 1172 -13656
rect 1142 -13716 1192 -13676
rect 1032 -13786 1192 -13716
rect 1032 -13826 1082 -13786
rect 1052 -13846 1082 -13826
rect 1142 -13826 1192 -13786
rect 1142 -13846 1172 -13826
rect 1252 -13886 1312 -13626
rect 912 -13896 992 -13886
rect 912 -13956 922 -13896
rect 982 -13906 992 -13896
rect 1232 -13896 1312 -13886
rect 1232 -13906 1242 -13896
rect 982 -13956 1242 -13906
rect 1302 -13956 1312 -13896
rect 912 -13966 1312 -13956
rect 1370 -13546 1770 -13536
rect 1370 -13606 1380 -13546
rect 1440 -13596 1700 -13546
rect 1440 -13606 1450 -13596
rect 1370 -13616 1450 -13606
rect 1690 -13606 1700 -13596
rect 1760 -13606 1770 -13546
rect 1690 -13616 1770 -13606
rect 1370 -13886 1430 -13616
rect 1700 -13626 1770 -13616
rect 1510 -13676 1540 -13656
rect 1490 -13716 1540 -13676
rect 1600 -13676 1630 -13656
rect 1600 -13716 1650 -13676
rect 1490 -13786 1650 -13716
rect 1490 -13826 1540 -13786
rect 1510 -13846 1540 -13826
rect 1600 -13826 1650 -13786
rect 1600 -13846 1630 -13826
rect 1710 -13886 1770 -13626
rect 1370 -13896 1450 -13886
rect 1370 -13956 1380 -13896
rect 1440 -13906 1450 -13896
rect 1690 -13896 1770 -13886
rect 1690 -13906 1700 -13896
rect 1440 -13956 1700 -13906
rect 1760 -13956 1770 -13896
rect 1370 -13966 1770 -13956
rect 1826 -13546 2226 -13536
rect 1826 -13606 1836 -13546
rect 1896 -13596 2156 -13546
rect 1896 -13606 1906 -13596
rect 1826 -13616 1906 -13606
rect 2146 -13606 2156 -13596
rect 2216 -13606 2226 -13546
rect 2146 -13616 2226 -13606
rect 1826 -13886 1886 -13616
rect 2156 -13626 2226 -13616
rect 1966 -13676 1996 -13656
rect 1946 -13716 1996 -13676
rect 2056 -13676 2086 -13656
rect 2056 -13716 2106 -13676
rect 1946 -13786 2106 -13716
rect 1946 -13826 1996 -13786
rect 1966 -13846 1996 -13826
rect 2056 -13826 2106 -13786
rect 2056 -13846 2086 -13826
rect 2166 -13886 2226 -13626
rect 1826 -13896 1906 -13886
rect 1826 -13956 1836 -13896
rect 1896 -13906 1906 -13896
rect 2146 -13896 2226 -13886
rect 2146 -13906 2156 -13896
rect 1896 -13956 2156 -13906
rect 2216 -13956 2226 -13896
rect 1826 -13966 2226 -13956
rect 2282 -13546 2682 -13536
rect 2282 -13606 2292 -13546
rect 2352 -13596 2612 -13546
rect 2352 -13606 2362 -13596
rect 2282 -13616 2362 -13606
rect 2602 -13606 2612 -13596
rect 2672 -13606 2682 -13546
rect 2602 -13616 2682 -13606
rect 2282 -13886 2342 -13616
rect 2612 -13626 2682 -13616
rect 2422 -13676 2452 -13656
rect 2402 -13716 2452 -13676
rect 2512 -13676 2542 -13656
rect 2512 -13716 2562 -13676
rect 2402 -13786 2562 -13716
rect 2402 -13826 2452 -13786
rect 2422 -13846 2452 -13826
rect 2512 -13826 2562 -13786
rect 2512 -13846 2542 -13826
rect 2622 -13886 2682 -13626
rect 2282 -13896 2362 -13886
rect 2282 -13956 2292 -13896
rect 2352 -13906 2362 -13896
rect 2602 -13896 2682 -13886
rect 2602 -13906 2612 -13896
rect 2352 -13956 2612 -13906
rect 2672 -13956 2682 -13896
rect 2282 -13966 2682 -13956
rect 2740 -13546 3140 -13536
rect 2740 -13606 2750 -13546
rect 2810 -13596 3070 -13546
rect 2810 -13606 2820 -13596
rect 2740 -13616 2820 -13606
rect 3060 -13606 3070 -13596
rect 3130 -13606 3140 -13546
rect 3060 -13616 3140 -13606
rect 2740 -13886 2800 -13616
rect 3070 -13626 3140 -13616
rect 2880 -13676 2910 -13656
rect 2860 -13716 2910 -13676
rect 2970 -13676 3000 -13656
rect 2970 -13716 3020 -13676
rect 2860 -13786 3020 -13716
rect 2860 -13826 2910 -13786
rect 2880 -13846 2910 -13826
rect 2970 -13826 3020 -13786
rect 2970 -13846 3000 -13826
rect 3080 -13886 3140 -13626
rect 2740 -13896 2820 -13886
rect 2740 -13956 2750 -13896
rect 2810 -13906 2820 -13896
rect 3060 -13896 3140 -13886
rect 3060 -13906 3070 -13896
rect 2810 -13956 3070 -13906
rect 3130 -13956 3140 -13896
rect 2740 -13966 3140 -13956
rect 3196 -13546 3596 -13536
rect 3196 -13606 3206 -13546
rect 3266 -13596 3526 -13546
rect 3266 -13606 3276 -13596
rect 3196 -13616 3276 -13606
rect 3516 -13606 3526 -13596
rect 3586 -13606 3596 -13546
rect 3516 -13616 3596 -13606
rect 3196 -13886 3256 -13616
rect 3526 -13626 3596 -13616
rect 3336 -13676 3366 -13656
rect 3316 -13716 3366 -13676
rect 3426 -13676 3456 -13656
rect 3426 -13716 3476 -13676
rect 3316 -13786 3476 -13716
rect 3316 -13826 3366 -13786
rect 3336 -13846 3366 -13826
rect 3426 -13826 3476 -13786
rect 3426 -13846 3456 -13826
rect 3536 -13886 3596 -13626
rect 3196 -13896 3276 -13886
rect 3196 -13956 3206 -13896
rect 3266 -13906 3276 -13896
rect 3516 -13896 3596 -13886
rect 3516 -13906 3526 -13896
rect 3266 -13956 3526 -13906
rect 3586 -13956 3596 -13896
rect 3196 -13966 3596 -13956
rect 3652 -13546 4052 -13536
rect 3652 -13606 3662 -13546
rect 3722 -13596 3982 -13546
rect 3722 -13606 3732 -13596
rect 3652 -13616 3732 -13606
rect 3972 -13606 3982 -13596
rect 4042 -13606 4052 -13546
rect 3972 -13616 4052 -13606
rect 3652 -13886 3712 -13616
rect 3982 -13626 4052 -13616
rect 3792 -13676 3822 -13656
rect 3772 -13716 3822 -13676
rect 3882 -13676 3912 -13656
rect 3882 -13716 3932 -13676
rect 3772 -13786 3932 -13716
rect 3772 -13826 3822 -13786
rect 3792 -13846 3822 -13826
rect 3882 -13826 3932 -13786
rect 3882 -13846 3912 -13826
rect 3992 -13886 4052 -13626
rect 3652 -13896 3732 -13886
rect 3652 -13956 3662 -13896
rect 3722 -13906 3732 -13896
rect 3972 -13896 4052 -13886
rect 3972 -13906 3982 -13896
rect 3722 -13956 3982 -13906
rect 4042 -13956 4052 -13896
rect 3652 -13966 4052 -13956
rect 4110 -13546 4510 -13536
rect 4110 -13606 4120 -13546
rect 4180 -13596 4440 -13546
rect 4180 -13606 4190 -13596
rect 4110 -13616 4190 -13606
rect 4430 -13606 4440 -13596
rect 4500 -13606 4510 -13546
rect 4430 -13616 4510 -13606
rect 4110 -13886 4170 -13616
rect 4440 -13626 4510 -13616
rect 4250 -13676 4280 -13656
rect 4230 -13716 4280 -13676
rect 4340 -13676 4370 -13656
rect 4340 -13716 4390 -13676
rect 4230 -13786 4390 -13716
rect 4230 -13826 4280 -13786
rect 4250 -13846 4280 -13826
rect 4340 -13826 4390 -13786
rect 4340 -13846 4370 -13826
rect 4450 -13886 4510 -13626
rect 4110 -13896 4190 -13886
rect 4110 -13956 4120 -13896
rect 4180 -13906 4190 -13896
rect 4430 -13896 4510 -13886
rect 4430 -13906 4440 -13896
rect 4180 -13956 4440 -13906
rect 4500 -13956 4510 -13896
rect 4110 -13966 4510 -13956
rect 4566 -13546 4966 -13536
rect 4566 -13606 4576 -13546
rect 4636 -13596 4896 -13546
rect 4636 -13606 4646 -13596
rect 4566 -13616 4646 -13606
rect 4886 -13606 4896 -13596
rect 4956 -13606 4966 -13546
rect 4886 -13616 4966 -13606
rect 4566 -13886 4626 -13616
rect 4896 -13626 4966 -13616
rect 4706 -13676 4736 -13656
rect 4686 -13716 4736 -13676
rect 4796 -13676 4826 -13656
rect 4796 -13716 4846 -13676
rect 4686 -13786 4846 -13716
rect 4686 -13826 4736 -13786
rect 4706 -13846 4736 -13826
rect 4796 -13826 4846 -13786
rect 4796 -13846 4826 -13826
rect 4906 -13886 4966 -13626
rect 4566 -13896 4646 -13886
rect 4566 -13956 4576 -13896
rect 4636 -13906 4646 -13896
rect 4886 -13896 4966 -13886
rect 4886 -13906 4896 -13896
rect 4636 -13956 4896 -13906
rect 4956 -13956 4966 -13896
rect 4566 -13966 4966 -13956
rect 5022 -13546 5422 -13536
rect 5022 -13606 5032 -13546
rect 5092 -13596 5352 -13546
rect 5092 -13606 5102 -13596
rect 5022 -13616 5102 -13606
rect 5342 -13606 5352 -13596
rect 5412 -13606 5422 -13546
rect 5342 -13616 5422 -13606
rect 5022 -13886 5082 -13616
rect 5352 -13626 5422 -13616
rect 5162 -13676 5192 -13656
rect 5142 -13716 5192 -13676
rect 5252 -13676 5282 -13656
rect 5252 -13716 5302 -13676
rect 5142 -13786 5302 -13716
rect 5142 -13826 5192 -13786
rect 5162 -13846 5192 -13826
rect 5252 -13826 5302 -13786
rect 5252 -13846 5282 -13826
rect 5362 -13886 5422 -13626
rect 5022 -13896 5102 -13886
rect 5022 -13956 5032 -13896
rect 5092 -13906 5102 -13896
rect 5342 -13896 5422 -13886
rect 5342 -13906 5352 -13896
rect 5092 -13956 5352 -13906
rect 5412 -13956 5422 -13896
rect 5022 -13966 5422 -13956
rect 5480 -13546 5880 -13536
rect 5480 -13606 5490 -13546
rect 5550 -13596 5810 -13546
rect 5550 -13606 5560 -13596
rect 5480 -13616 5560 -13606
rect 5800 -13606 5810 -13596
rect 5870 -13606 5880 -13546
rect 5800 -13616 5880 -13606
rect 5480 -13886 5540 -13616
rect 5810 -13626 5880 -13616
rect 5620 -13676 5650 -13656
rect 5600 -13716 5650 -13676
rect 5710 -13676 5740 -13656
rect 5710 -13716 5760 -13676
rect 5600 -13786 5760 -13716
rect 5600 -13826 5650 -13786
rect 5620 -13846 5650 -13826
rect 5710 -13826 5760 -13786
rect 5710 -13846 5740 -13826
rect 5820 -13886 5880 -13626
rect 5480 -13896 5560 -13886
rect 5480 -13956 5490 -13896
rect 5550 -13906 5560 -13896
rect 5800 -13896 5880 -13886
rect 5800 -13906 5810 -13896
rect 5550 -13956 5810 -13906
rect 5870 -13956 5880 -13896
rect 5480 -13966 5880 -13956
rect 5936 -13546 6336 -13536
rect 5936 -13606 5946 -13546
rect 6006 -13596 6266 -13546
rect 6006 -13606 6016 -13596
rect 5936 -13616 6016 -13606
rect 6256 -13606 6266 -13596
rect 6326 -13606 6336 -13546
rect 6256 -13616 6336 -13606
rect 5936 -13886 5996 -13616
rect 6266 -13626 6336 -13616
rect 6076 -13676 6106 -13656
rect 6056 -13716 6106 -13676
rect 6166 -13676 6196 -13656
rect 6166 -13716 6216 -13676
rect 6056 -13786 6216 -13716
rect 6056 -13826 6106 -13786
rect 6076 -13846 6106 -13826
rect 6166 -13826 6216 -13786
rect 6166 -13846 6196 -13826
rect 6276 -13886 6336 -13626
rect 5936 -13896 6016 -13886
rect 5936 -13956 5946 -13896
rect 6006 -13906 6016 -13896
rect 6256 -13896 6336 -13886
rect 6256 -13906 6266 -13896
rect 6006 -13956 6266 -13906
rect 6326 -13956 6336 -13896
rect 5936 -13966 6336 -13956
rect 6392 -13546 6792 -13536
rect 6392 -13606 6402 -13546
rect 6462 -13596 6722 -13546
rect 6462 -13606 6472 -13596
rect 6392 -13616 6472 -13606
rect 6712 -13606 6722 -13596
rect 6782 -13606 6792 -13546
rect 6712 -13616 6792 -13606
rect 6392 -13886 6452 -13616
rect 6722 -13626 6792 -13616
rect 6532 -13676 6562 -13656
rect 6512 -13716 6562 -13676
rect 6622 -13676 6652 -13656
rect 6622 -13716 6672 -13676
rect 6512 -13786 6672 -13716
rect 6512 -13826 6562 -13786
rect 6532 -13846 6562 -13826
rect 6622 -13826 6672 -13786
rect 6622 -13846 6652 -13826
rect 6732 -13886 6792 -13626
rect 6392 -13896 6472 -13886
rect 6392 -13956 6402 -13896
rect 6462 -13906 6472 -13896
rect 6712 -13896 6792 -13886
rect 6712 -13906 6722 -13896
rect 6462 -13956 6722 -13906
rect 6782 -13956 6792 -13896
rect 6392 -13966 6792 -13956
rect 6850 -13546 7250 -13536
rect 6850 -13606 6860 -13546
rect 6920 -13596 7180 -13546
rect 6920 -13606 6930 -13596
rect 6850 -13616 6930 -13606
rect 7170 -13606 7180 -13596
rect 7240 -13606 7250 -13546
rect 7170 -13616 7250 -13606
rect 6850 -13886 6910 -13616
rect 7180 -13626 7250 -13616
rect 6990 -13676 7020 -13656
rect 6970 -13716 7020 -13676
rect 7080 -13676 7110 -13656
rect 7080 -13716 7130 -13676
rect 6970 -13786 7130 -13716
rect 6970 -13826 7020 -13786
rect 6990 -13846 7020 -13826
rect 7080 -13826 7130 -13786
rect 7080 -13846 7110 -13826
rect 7190 -13886 7250 -13626
rect 6850 -13896 6930 -13886
rect 6850 -13956 6860 -13896
rect 6920 -13906 6930 -13896
rect 7170 -13896 7250 -13886
rect 7170 -13906 7180 -13896
rect 6920 -13956 7180 -13906
rect 7240 -13956 7250 -13896
rect 6850 -13966 7250 -13956
rect 7306 -13546 7706 -13536
rect 7306 -13606 7316 -13546
rect 7376 -13596 7636 -13546
rect 7376 -13606 7386 -13596
rect 7306 -13616 7386 -13606
rect 7626 -13606 7636 -13596
rect 7696 -13606 7706 -13546
rect 7626 -13616 7706 -13606
rect 7306 -13886 7366 -13616
rect 7636 -13626 7706 -13616
rect 7446 -13676 7476 -13656
rect 7426 -13716 7476 -13676
rect 7536 -13676 7566 -13656
rect 7536 -13716 7586 -13676
rect 7426 -13786 7586 -13716
rect 7426 -13826 7476 -13786
rect 7446 -13846 7476 -13826
rect 7536 -13826 7586 -13786
rect 7536 -13846 7566 -13826
rect 7646 -13886 7706 -13626
rect 7306 -13896 7386 -13886
rect 7306 -13956 7316 -13896
rect 7376 -13906 7386 -13896
rect 7626 -13896 7706 -13886
rect 7626 -13906 7636 -13896
rect 7376 -13956 7636 -13906
rect 7696 -13956 7706 -13896
rect 7306 -13966 7706 -13956
rect 7762 -13546 8162 -13536
rect 7762 -13606 7772 -13546
rect 7832 -13596 8092 -13546
rect 7832 -13606 7842 -13596
rect 7762 -13616 7842 -13606
rect 8082 -13606 8092 -13596
rect 8152 -13606 8162 -13546
rect 8082 -13616 8162 -13606
rect 7762 -13886 7822 -13616
rect 8092 -13626 8162 -13616
rect 7902 -13676 7932 -13656
rect 7882 -13716 7932 -13676
rect 7992 -13676 8022 -13656
rect 7992 -13716 8042 -13676
rect 7882 -13786 8042 -13716
rect 7882 -13826 7932 -13786
rect 7902 -13846 7932 -13826
rect 7992 -13826 8042 -13786
rect 7992 -13846 8022 -13826
rect 8102 -13886 8162 -13626
rect 7762 -13896 7842 -13886
rect 7762 -13956 7772 -13896
rect 7832 -13906 7842 -13896
rect 8082 -13896 8162 -13886
rect 8082 -13906 8092 -13896
rect 7832 -13956 8092 -13906
rect 8152 -13956 8162 -13896
rect 7762 -13966 8162 -13956
rect 8236 -13546 8636 -13536
rect 8236 -13606 8246 -13546
rect 8306 -13596 8566 -13546
rect 8306 -13606 8316 -13596
rect 8236 -13616 8316 -13606
rect 8556 -13606 8566 -13596
rect 8626 -13606 8636 -13546
rect 8556 -13616 8636 -13606
rect 8236 -13886 8296 -13616
rect 8566 -13626 8636 -13616
rect 8376 -13676 8406 -13656
rect 8356 -13716 8406 -13676
rect 8466 -13676 8496 -13656
rect 8466 -13716 8516 -13676
rect 8356 -13786 8516 -13716
rect 8356 -13826 8406 -13786
rect 8376 -13846 8406 -13826
rect 8466 -13826 8516 -13786
rect 8466 -13846 8496 -13826
rect 8576 -13886 8636 -13626
rect 8236 -13896 8316 -13886
rect 8236 -13956 8246 -13896
rect 8306 -13906 8316 -13896
rect 8556 -13896 8636 -13886
rect 8556 -13906 8566 -13896
rect 8306 -13956 8566 -13906
rect 8626 -13956 8636 -13896
rect 8236 -13966 8636 -13956
rect 8692 -13546 9092 -13536
rect 8692 -13606 8702 -13546
rect 8762 -13596 9022 -13546
rect 8762 -13606 8772 -13596
rect 8692 -13616 8772 -13606
rect 9012 -13606 9022 -13596
rect 9082 -13606 9092 -13546
rect 9012 -13616 9092 -13606
rect 8692 -13886 8752 -13616
rect 9022 -13626 9092 -13616
rect 8832 -13676 8862 -13656
rect 8812 -13716 8862 -13676
rect 8922 -13676 8952 -13656
rect 8922 -13716 8972 -13676
rect 8812 -13786 8972 -13716
rect 8812 -13826 8862 -13786
rect 8832 -13846 8862 -13826
rect 8922 -13826 8972 -13786
rect 8922 -13846 8952 -13826
rect 9032 -13886 9092 -13626
rect 8692 -13896 8772 -13886
rect 8692 -13956 8702 -13896
rect 8762 -13906 8772 -13896
rect 9012 -13896 9092 -13886
rect 9012 -13906 9022 -13896
rect 8762 -13956 9022 -13906
rect 9082 -13956 9092 -13896
rect 8692 -13966 9092 -13956
rect 9150 -13546 9550 -13536
rect 9150 -13606 9160 -13546
rect 9220 -13596 9480 -13546
rect 9220 -13606 9230 -13596
rect 9150 -13616 9230 -13606
rect 9470 -13606 9480 -13596
rect 9540 -13606 9550 -13546
rect 9470 -13616 9550 -13606
rect 9150 -13886 9210 -13616
rect 9480 -13626 9550 -13616
rect 9290 -13676 9320 -13656
rect 9270 -13716 9320 -13676
rect 9380 -13676 9410 -13656
rect 9380 -13716 9430 -13676
rect 9270 -13786 9430 -13716
rect 9270 -13826 9320 -13786
rect 9290 -13846 9320 -13826
rect 9380 -13826 9430 -13786
rect 9380 -13846 9410 -13826
rect 9490 -13886 9550 -13626
rect 9150 -13896 9230 -13886
rect 9150 -13956 9160 -13896
rect 9220 -13906 9230 -13896
rect 9470 -13896 9550 -13886
rect 9470 -13906 9480 -13896
rect 9220 -13956 9480 -13906
rect 9540 -13956 9550 -13896
rect 9150 -13966 9550 -13956
rect 9606 -13546 10006 -13536
rect 9606 -13606 9616 -13546
rect 9676 -13596 9936 -13546
rect 9676 -13606 9686 -13596
rect 9606 -13616 9686 -13606
rect 9926 -13606 9936 -13596
rect 9996 -13606 10006 -13546
rect 9926 -13616 10006 -13606
rect 9606 -13886 9666 -13616
rect 9936 -13626 10006 -13616
rect 9746 -13676 9776 -13656
rect 9726 -13716 9776 -13676
rect 9836 -13676 9866 -13656
rect 9836 -13716 9886 -13676
rect 9726 -13786 9886 -13716
rect 9726 -13826 9776 -13786
rect 9746 -13846 9776 -13826
rect 9836 -13826 9886 -13786
rect 9836 -13846 9866 -13826
rect 9946 -13886 10006 -13626
rect 9606 -13896 9686 -13886
rect 9606 -13956 9616 -13896
rect 9676 -13906 9686 -13896
rect 9926 -13896 10006 -13886
rect 9926 -13906 9936 -13896
rect 9676 -13956 9936 -13906
rect 9996 -13956 10006 -13896
rect 9606 -13966 10006 -13956
rect 10062 -13546 10462 -13536
rect 10062 -13606 10072 -13546
rect 10132 -13596 10392 -13546
rect 10132 -13606 10142 -13596
rect 10062 -13616 10142 -13606
rect 10382 -13606 10392 -13596
rect 10452 -13606 10462 -13546
rect 10382 -13616 10462 -13606
rect 10062 -13886 10122 -13616
rect 10392 -13626 10462 -13616
rect 10202 -13676 10232 -13656
rect 10182 -13716 10232 -13676
rect 10292 -13676 10322 -13656
rect 10292 -13716 10342 -13676
rect 10182 -13786 10342 -13716
rect 10182 -13826 10232 -13786
rect 10202 -13846 10232 -13826
rect 10292 -13826 10342 -13786
rect 10292 -13846 10322 -13826
rect 10402 -13886 10462 -13626
rect 10062 -13896 10142 -13886
rect 10062 -13956 10072 -13896
rect 10132 -13906 10142 -13896
rect 10382 -13896 10462 -13886
rect 10382 -13906 10392 -13896
rect 10132 -13956 10392 -13906
rect 10452 -13956 10462 -13896
rect 10062 -13966 10462 -13956
rect 10520 -13546 10920 -13536
rect 10520 -13606 10530 -13546
rect 10590 -13596 10850 -13546
rect 10590 -13606 10600 -13596
rect 10520 -13616 10600 -13606
rect 10840 -13606 10850 -13596
rect 10910 -13606 10920 -13546
rect 10840 -13616 10920 -13606
rect 10520 -13886 10580 -13616
rect 10850 -13626 10920 -13616
rect 10660 -13676 10690 -13656
rect 10640 -13716 10690 -13676
rect 10750 -13676 10780 -13656
rect 10750 -13716 10800 -13676
rect 10640 -13786 10800 -13716
rect 10640 -13826 10690 -13786
rect 10660 -13846 10690 -13826
rect 10750 -13826 10800 -13786
rect 10750 -13846 10780 -13826
rect 10860 -13886 10920 -13626
rect 10520 -13896 10600 -13886
rect 10520 -13956 10530 -13896
rect 10590 -13906 10600 -13896
rect 10840 -13896 10920 -13886
rect 10840 -13906 10850 -13896
rect 10590 -13956 10850 -13906
rect 10910 -13956 10920 -13896
rect 10520 -13966 10920 -13956
rect 10976 -13546 11376 -13536
rect 10976 -13606 10986 -13546
rect 11046 -13596 11306 -13546
rect 11046 -13606 11056 -13596
rect 10976 -13616 11056 -13606
rect 11296 -13606 11306 -13596
rect 11366 -13606 11376 -13546
rect 11296 -13616 11376 -13606
rect 10976 -13886 11036 -13616
rect 11306 -13626 11376 -13616
rect 11116 -13676 11146 -13656
rect 11096 -13716 11146 -13676
rect 11206 -13676 11236 -13656
rect 11206 -13716 11256 -13676
rect 11096 -13786 11256 -13716
rect 11096 -13826 11146 -13786
rect 11116 -13846 11146 -13826
rect 11206 -13826 11256 -13786
rect 11206 -13846 11236 -13826
rect 11316 -13886 11376 -13626
rect 10976 -13896 11056 -13886
rect 10976 -13956 10986 -13896
rect 11046 -13906 11056 -13896
rect 11296 -13896 11376 -13886
rect 11296 -13906 11306 -13896
rect 11046 -13956 11306 -13906
rect 11366 -13956 11376 -13896
rect 10976 -13966 11376 -13956
rect 11432 -13546 11832 -13536
rect 11432 -13606 11442 -13546
rect 11502 -13596 11762 -13546
rect 11502 -13606 11512 -13596
rect 11432 -13616 11512 -13606
rect 11752 -13606 11762 -13596
rect 11822 -13606 11832 -13546
rect 11752 -13616 11832 -13606
rect 11432 -13886 11492 -13616
rect 11762 -13626 11832 -13616
rect 11572 -13676 11602 -13656
rect 11552 -13716 11602 -13676
rect 11662 -13676 11692 -13656
rect 11662 -13716 11712 -13676
rect 11552 -13786 11712 -13716
rect 11552 -13826 11602 -13786
rect 11572 -13846 11602 -13826
rect 11662 -13826 11712 -13786
rect 11662 -13846 11692 -13826
rect 11772 -13886 11832 -13626
rect 11432 -13896 11512 -13886
rect 11432 -13956 11442 -13896
rect 11502 -13906 11512 -13896
rect 11752 -13896 11832 -13886
rect 11752 -13906 11762 -13896
rect 11502 -13956 11762 -13906
rect 11822 -13956 11832 -13896
rect 11432 -13966 11832 -13956
rect 11890 -13546 12290 -13536
rect 11890 -13606 11900 -13546
rect 11960 -13596 12220 -13546
rect 11960 -13606 11970 -13596
rect 11890 -13616 11970 -13606
rect 12210 -13606 12220 -13596
rect 12280 -13606 12290 -13546
rect 12210 -13616 12290 -13606
rect 11890 -13886 11950 -13616
rect 12220 -13626 12290 -13616
rect 12030 -13676 12060 -13656
rect 12010 -13716 12060 -13676
rect 12120 -13676 12150 -13656
rect 12120 -13716 12170 -13676
rect 12010 -13786 12170 -13716
rect 12010 -13826 12060 -13786
rect 12030 -13846 12060 -13826
rect 12120 -13826 12170 -13786
rect 12120 -13846 12150 -13826
rect 12230 -13886 12290 -13626
rect 11890 -13896 11970 -13886
rect 11890 -13956 11900 -13896
rect 11960 -13906 11970 -13896
rect 12210 -13896 12290 -13886
rect 12210 -13906 12220 -13896
rect 11960 -13956 12220 -13906
rect 12280 -13956 12290 -13896
rect 11890 -13966 12290 -13956
rect 12346 -13546 12746 -13536
rect 12346 -13606 12356 -13546
rect 12416 -13596 12676 -13546
rect 12416 -13606 12426 -13596
rect 12346 -13616 12426 -13606
rect 12666 -13606 12676 -13596
rect 12736 -13606 12746 -13546
rect 12666 -13616 12746 -13606
rect 12346 -13886 12406 -13616
rect 12676 -13626 12746 -13616
rect 12486 -13676 12516 -13656
rect 12466 -13716 12516 -13676
rect 12576 -13676 12606 -13656
rect 12576 -13716 12626 -13676
rect 12466 -13786 12626 -13716
rect 12466 -13826 12516 -13786
rect 12486 -13846 12516 -13826
rect 12576 -13826 12626 -13786
rect 12576 -13846 12606 -13826
rect 12686 -13886 12746 -13626
rect 12346 -13896 12426 -13886
rect 12346 -13956 12356 -13896
rect 12416 -13906 12426 -13896
rect 12666 -13896 12746 -13886
rect 12666 -13906 12676 -13896
rect 12416 -13956 12676 -13906
rect 12736 -13956 12746 -13896
rect 12346 -13966 12746 -13956
rect 12802 -13546 13202 -13536
rect 12802 -13606 12812 -13546
rect 12872 -13596 13132 -13546
rect 12872 -13606 12882 -13596
rect 12802 -13616 12882 -13606
rect 13122 -13606 13132 -13596
rect 13192 -13606 13202 -13546
rect 13122 -13616 13202 -13606
rect 12802 -13886 12862 -13616
rect 13132 -13626 13202 -13616
rect 12942 -13676 12972 -13656
rect 12922 -13716 12972 -13676
rect 13032 -13676 13062 -13656
rect 13032 -13716 13082 -13676
rect 12922 -13786 13082 -13716
rect 12922 -13826 12972 -13786
rect 12942 -13846 12972 -13826
rect 13032 -13826 13082 -13786
rect 13032 -13846 13062 -13826
rect 13142 -13886 13202 -13626
rect 12802 -13896 12882 -13886
rect 12802 -13956 12812 -13896
rect 12872 -13906 12882 -13896
rect 13122 -13896 13202 -13886
rect 13122 -13906 13132 -13896
rect 12872 -13956 13132 -13906
rect 13192 -13956 13202 -13896
rect 12802 -13966 13202 -13956
rect 13260 -13546 13660 -13536
rect 13260 -13606 13270 -13546
rect 13330 -13596 13590 -13546
rect 13330 -13606 13340 -13596
rect 13260 -13616 13340 -13606
rect 13580 -13606 13590 -13596
rect 13650 -13606 13660 -13546
rect 13580 -13616 13660 -13606
rect 13260 -13886 13320 -13616
rect 13590 -13626 13660 -13616
rect 13400 -13676 13430 -13656
rect 13380 -13716 13430 -13676
rect 13490 -13676 13520 -13656
rect 13490 -13716 13540 -13676
rect 13380 -13786 13540 -13716
rect 13380 -13826 13430 -13786
rect 13400 -13846 13430 -13826
rect 13490 -13826 13540 -13786
rect 13490 -13846 13520 -13826
rect 13600 -13886 13660 -13626
rect 13260 -13896 13340 -13886
rect 13260 -13956 13270 -13896
rect 13330 -13906 13340 -13896
rect 13580 -13896 13660 -13886
rect 13580 -13906 13590 -13896
rect 13330 -13956 13590 -13906
rect 13650 -13956 13660 -13896
rect 13260 -13966 13660 -13956
rect 13716 -13546 14116 -13536
rect 13716 -13606 13726 -13546
rect 13786 -13596 14046 -13546
rect 13786 -13606 13796 -13596
rect 13716 -13616 13796 -13606
rect 14036 -13606 14046 -13596
rect 14106 -13606 14116 -13546
rect 14036 -13616 14116 -13606
rect 13716 -13886 13776 -13616
rect 14046 -13626 14116 -13616
rect 13856 -13676 13886 -13656
rect 13836 -13716 13886 -13676
rect 13946 -13676 13976 -13656
rect 13946 -13716 13996 -13676
rect 13836 -13786 13996 -13716
rect 13836 -13826 13886 -13786
rect 13856 -13846 13886 -13826
rect 13946 -13826 13996 -13786
rect 13946 -13846 13976 -13826
rect 14056 -13886 14116 -13626
rect 13716 -13896 13796 -13886
rect 13716 -13956 13726 -13896
rect 13786 -13906 13796 -13896
rect 14036 -13896 14116 -13886
rect 14036 -13906 14046 -13896
rect 13786 -13956 14046 -13906
rect 14106 -13956 14116 -13896
rect 13716 -13966 14116 -13956
rect 14172 -13546 14572 -13536
rect 14172 -13606 14182 -13546
rect 14242 -13596 14502 -13546
rect 14242 -13606 14252 -13596
rect 14172 -13616 14252 -13606
rect 14492 -13606 14502 -13596
rect 14562 -13606 14572 -13546
rect 14492 -13616 14572 -13606
rect 14172 -13886 14232 -13616
rect 14502 -13626 14572 -13616
rect 14312 -13676 14342 -13656
rect 14292 -13716 14342 -13676
rect 14402 -13676 14432 -13656
rect 14402 -13716 14452 -13676
rect 14292 -13786 14452 -13716
rect 14292 -13826 14342 -13786
rect 14312 -13846 14342 -13826
rect 14402 -13826 14452 -13786
rect 14402 -13846 14432 -13826
rect 14512 -13886 14572 -13626
rect 14172 -13896 14252 -13886
rect 14172 -13956 14182 -13896
rect 14242 -13906 14252 -13896
rect 14492 -13896 14572 -13886
rect 14492 -13906 14502 -13896
rect 14242 -13956 14502 -13906
rect 14562 -13956 14572 -13896
rect 14172 -13966 14572 -13956
rect 14630 -13546 15030 -13536
rect 14630 -13606 14640 -13546
rect 14700 -13596 14960 -13546
rect 14700 -13606 14710 -13596
rect 14630 -13616 14710 -13606
rect 14950 -13606 14960 -13596
rect 15020 -13606 15030 -13546
rect 14950 -13616 15030 -13606
rect 14630 -13886 14690 -13616
rect 14960 -13626 15030 -13616
rect 14770 -13676 14800 -13656
rect 14750 -13716 14800 -13676
rect 14860 -13676 14890 -13656
rect 14860 -13716 14910 -13676
rect 14750 -13786 14910 -13716
rect 14750 -13826 14800 -13786
rect 14770 -13846 14800 -13826
rect 14860 -13826 14910 -13786
rect 14860 -13846 14890 -13826
rect 14970 -13886 15030 -13626
rect 14630 -13896 14710 -13886
rect 14630 -13956 14640 -13896
rect 14700 -13906 14710 -13896
rect 14950 -13896 15030 -13886
rect 14950 -13906 14960 -13896
rect 14700 -13956 14960 -13906
rect 15020 -13956 15030 -13896
rect 14630 -13966 15030 -13956
rect 15086 -13546 15486 -13536
rect 15086 -13606 15096 -13546
rect 15156 -13596 15416 -13546
rect 15156 -13606 15166 -13596
rect 15086 -13616 15166 -13606
rect 15406 -13606 15416 -13596
rect 15476 -13606 15486 -13546
rect 15406 -13616 15486 -13606
rect 15086 -13886 15146 -13616
rect 15416 -13626 15486 -13616
rect 15226 -13676 15256 -13656
rect 15206 -13716 15256 -13676
rect 15316 -13676 15346 -13656
rect 15316 -13716 15366 -13676
rect 15206 -13786 15366 -13716
rect 15206 -13826 15256 -13786
rect 15226 -13846 15256 -13826
rect 15316 -13826 15366 -13786
rect 15316 -13846 15346 -13826
rect 15426 -13886 15486 -13626
rect 15086 -13896 15166 -13886
rect 15086 -13956 15096 -13896
rect 15156 -13906 15166 -13896
rect 15406 -13896 15486 -13886
rect 15406 -13906 15416 -13896
rect 15156 -13956 15416 -13906
rect 15476 -13956 15486 -13896
rect 15086 -13966 15486 -13956
rect 0 -14040 400 -14030
rect 0 -14100 10 -14040
rect 70 -14090 330 -14040
rect 70 -14100 80 -14090
rect 0 -14110 80 -14100
rect 320 -14100 330 -14090
rect 390 -14100 400 -14040
rect 320 -14110 400 -14100
rect 0 -14380 60 -14110
rect 330 -14120 400 -14110
rect 140 -14170 170 -14150
rect 120 -14210 170 -14170
rect 230 -14170 260 -14150
rect 230 -14210 280 -14170
rect 120 -14280 280 -14210
rect 120 -14320 170 -14280
rect 140 -14340 170 -14320
rect 230 -14320 280 -14280
rect 230 -14340 260 -14320
rect 340 -14380 400 -14120
rect 0 -14390 80 -14380
rect 0 -14450 10 -14390
rect 70 -14400 80 -14390
rect 320 -14390 400 -14380
rect 320 -14400 330 -14390
rect 70 -14450 330 -14400
rect 390 -14450 400 -14390
rect 0 -14460 400 -14450
rect 456 -14040 856 -14030
rect 456 -14100 466 -14040
rect 526 -14090 786 -14040
rect 526 -14100 536 -14090
rect 456 -14110 536 -14100
rect 776 -14100 786 -14090
rect 846 -14100 856 -14040
rect 776 -14110 856 -14100
rect 456 -14380 516 -14110
rect 786 -14120 856 -14110
rect 596 -14170 626 -14150
rect 576 -14210 626 -14170
rect 686 -14170 716 -14150
rect 686 -14210 736 -14170
rect 576 -14280 736 -14210
rect 576 -14320 626 -14280
rect 596 -14340 626 -14320
rect 686 -14320 736 -14280
rect 686 -14340 716 -14320
rect 796 -14380 856 -14120
rect 456 -14390 536 -14380
rect 456 -14450 466 -14390
rect 526 -14400 536 -14390
rect 776 -14390 856 -14380
rect 776 -14400 786 -14390
rect 526 -14450 786 -14400
rect 846 -14450 856 -14390
rect 456 -14460 856 -14450
rect 912 -14040 1312 -14030
rect 912 -14100 922 -14040
rect 982 -14090 1242 -14040
rect 982 -14100 992 -14090
rect 912 -14110 992 -14100
rect 1232 -14100 1242 -14090
rect 1302 -14100 1312 -14040
rect 1232 -14110 1312 -14100
rect 912 -14380 972 -14110
rect 1242 -14120 1312 -14110
rect 1052 -14170 1082 -14150
rect 1032 -14210 1082 -14170
rect 1142 -14170 1172 -14150
rect 1142 -14210 1192 -14170
rect 1032 -14280 1192 -14210
rect 1032 -14320 1082 -14280
rect 1052 -14340 1082 -14320
rect 1142 -14320 1192 -14280
rect 1142 -14340 1172 -14320
rect 1252 -14380 1312 -14120
rect 912 -14390 992 -14380
rect 912 -14450 922 -14390
rect 982 -14400 992 -14390
rect 1232 -14390 1312 -14380
rect 1232 -14400 1242 -14390
rect 982 -14450 1242 -14400
rect 1302 -14450 1312 -14390
rect 912 -14460 1312 -14450
rect 1370 -14040 1770 -14030
rect 1370 -14100 1380 -14040
rect 1440 -14090 1700 -14040
rect 1440 -14100 1450 -14090
rect 1370 -14110 1450 -14100
rect 1690 -14100 1700 -14090
rect 1760 -14100 1770 -14040
rect 1690 -14110 1770 -14100
rect 1370 -14380 1430 -14110
rect 1700 -14120 1770 -14110
rect 1510 -14170 1540 -14150
rect 1490 -14210 1540 -14170
rect 1600 -14170 1630 -14150
rect 1600 -14210 1650 -14170
rect 1490 -14280 1650 -14210
rect 1490 -14320 1540 -14280
rect 1510 -14340 1540 -14320
rect 1600 -14320 1650 -14280
rect 1600 -14340 1630 -14320
rect 1710 -14380 1770 -14120
rect 1370 -14390 1450 -14380
rect 1370 -14450 1380 -14390
rect 1440 -14400 1450 -14390
rect 1690 -14390 1770 -14380
rect 1690 -14400 1700 -14390
rect 1440 -14450 1700 -14400
rect 1760 -14450 1770 -14390
rect 1370 -14460 1770 -14450
rect 1826 -14040 2226 -14030
rect 1826 -14100 1836 -14040
rect 1896 -14090 2156 -14040
rect 1896 -14100 1906 -14090
rect 1826 -14110 1906 -14100
rect 2146 -14100 2156 -14090
rect 2216 -14100 2226 -14040
rect 2146 -14110 2226 -14100
rect 1826 -14380 1886 -14110
rect 2156 -14120 2226 -14110
rect 1966 -14170 1996 -14150
rect 1946 -14210 1996 -14170
rect 2056 -14170 2086 -14150
rect 2056 -14210 2106 -14170
rect 1946 -14280 2106 -14210
rect 1946 -14320 1996 -14280
rect 1966 -14340 1996 -14320
rect 2056 -14320 2106 -14280
rect 2056 -14340 2086 -14320
rect 2166 -14380 2226 -14120
rect 1826 -14390 1906 -14380
rect 1826 -14450 1836 -14390
rect 1896 -14400 1906 -14390
rect 2146 -14390 2226 -14380
rect 2146 -14400 2156 -14390
rect 1896 -14450 2156 -14400
rect 2216 -14450 2226 -14390
rect 1826 -14460 2226 -14450
rect 2282 -14040 2682 -14030
rect 2282 -14100 2292 -14040
rect 2352 -14090 2612 -14040
rect 2352 -14100 2362 -14090
rect 2282 -14110 2362 -14100
rect 2602 -14100 2612 -14090
rect 2672 -14100 2682 -14040
rect 2602 -14110 2682 -14100
rect 2282 -14380 2342 -14110
rect 2612 -14120 2682 -14110
rect 2422 -14170 2452 -14150
rect 2402 -14210 2452 -14170
rect 2512 -14170 2542 -14150
rect 2512 -14210 2562 -14170
rect 2402 -14280 2562 -14210
rect 2402 -14320 2452 -14280
rect 2422 -14340 2452 -14320
rect 2512 -14320 2562 -14280
rect 2512 -14340 2542 -14320
rect 2622 -14380 2682 -14120
rect 2282 -14390 2362 -14380
rect 2282 -14450 2292 -14390
rect 2352 -14400 2362 -14390
rect 2602 -14390 2682 -14380
rect 2602 -14400 2612 -14390
rect 2352 -14450 2612 -14400
rect 2672 -14450 2682 -14390
rect 2282 -14460 2682 -14450
rect 2740 -14040 3140 -14030
rect 2740 -14100 2750 -14040
rect 2810 -14090 3070 -14040
rect 2810 -14100 2820 -14090
rect 2740 -14110 2820 -14100
rect 3060 -14100 3070 -14090
rect 3130 -14100 3140 -14040
rect 3060 -14110 3140 -14100
rect 2740 -14380 2800 -14110
rect 3070 -14120 3140 -14110
rect 2880 -14170 2910 -14150
rect 2860 -14210 2910 -14170
rect 2970 -14170 3000 -14150
rect 2970 -14210 3020 -14170
rect 2860 -14280 3020 -14210
rect 2860 -14320 2910 -14280
rect 2880 -14340 2910 -14320
rect 2970 -14320 3020 -14280
rect 2970 -14340 3000 -14320
rect 3080 -14380 3140 -14120
rect 2740 -14390 2820 -14380
rect 2740 -14450 2750 -14390
rect 2810 -14400 2820 -14390
rect 3060 -14390 3140 -14380
rect 3060 -14400 3070 -14390
rect 2810 -14450 3070 -14400
rect 3130 -14450 3140 -14390
rect 2740 -14460 3140 -14450
rect 3196 -14040 3596 -14030
rect 3196 -14100 3206 -14040
rect 3266 -14090 3526 -14040
rect 3266 -14100 3276 -14090
rect 3196 -14110 3276 -14100
rect 3516 -14100 3526 -14090
rect 3586 -14100 3596 -14040
rect 3516 -14110 3596 -14100
rect 3196 -14380 3256 -14110
rect 3526 -14120 3596 -14110
rect 3336 -14170 3366 -14150
rect 3316 -14210 3366 -14170
rect 3426 -14170 3456 -14150
rect 3426 -14210 3476 -14170
rect 3316 -14280 3476 -14210
rect 3316 -14320 3366 -14280
rect 3336 -14340 3366 -14320
rect 3426 -14320 3476 -14280
rect 3426 -14340 3456 -14320
rect 3536 -14380 3596 -14120
rect 3196 -14390 3276 -14380
rect 3196 -14450 3206 -14390
rect 3266 -14400 3276 -14390
rect 3516 -14390 3596 -14380
rect 3516 -14400 3526 -14390
rect 3266 -14450 3526 -14400
rect 3586 -14450 3596 -14390
rect 3196 -14460 3596 -14450
rect 3652 -14040 4052 -14030
rect 3652 -14100 3662 -14040
rect 3722 -14090 3982 -14040
rect 3722 -14100 3732 -14090
rect 3652 -14110 3732 -14100
rect 3972 -14100 3982 -14090
rect 4042 -14100 4052 -14040
rect 3972 -14110 4052 -14100
rect 3652 -14380 3712 -14110
rect 3982 -14120 4052 -14110
rect 3792 -14170 3822 -14150
rect 3772 -14210 3822 -14170
rect 3882 -14170 3912 -14150
rect 3882 -14210 3932 -14170
rect 3772 -14280 3932 -14210
rect 3772 -14320 3822 -14280
rect 3792 -14340 3822 -14320
rect 3882 -14320 3932 -14280
rect 3882 -14340 3912 -14320
rect 3992 -14380 4052 -14120
rect 3652 -14390 3732 -14380
rect 3652 -14450 3662 -14390
rect 3722 -14400 3732 -14390
rect 3972 -14390 4052 -14380
rect 3972 -14400 3982 -14390
rect 3722 -14450 3982 -14400
rect 4042 -14450 4052 -14390
rect 3652 -14460 4052 -14450
rect 4110 -14040 4510 -14030
rect 4110 -14100 4120 -14040
rect 4180 -14090 4440 -14040
rect 4180 -14100 4190 -14090
rect 4110 -14110 4190 -14100
rect 4430 -14100 4440 -14090
rect 4500 -14100 4510 -14040
rect 4430 -14110 4510 -14100
rect 4110 -14380 4170 -14110
rect 4440 -14120 4510 -14110
rect 4250 -14170 4280 -14150
rect 4230 -14210 4280 -14170
rect 4340 -14170 4370 -14150
rect 4340 -14210 4390 -14170
rect 4230 -14280 4390 -14210
rect 4230 -14320 4280 -14280
rect 4250 -14340 4280 -14320
rect 4340 -14320 4390 -14280
rect 4340 -14340 4370 -14320
rect 4450 -14380 4510 -14120
rect 4110 -14390 4190 -14380
rect 4110 -14450 4120 -14390
rect 4180 -14400 4190 -14390
rect 4430 -14390 4510 -14380
rect 4430 -14400 4440 -14390
rect 4180 -14450 4440 -14400
rect 4500 -14450 4510 -14390
rect 4110 -14460 4510 -14450
rect 4566 -14040 4966 -14030
rect 4566 -14100 4576 -14040
rect 4636 -14090 4896 -14040
rect 4636 -14100 4646 -14090
rect 4566 -14110 4646 -14100
rect 4886 -14100 4896 -14090
rect 4956 -14100 4966 -14040
rect 4886 -14110 4966 -14100
rect 4566 -14380 4626 -14110
rect 4896 -14120 4966 -14110
rect 4706 -14170 4736 -14150
rect 4686 -14210 4736 -14170
rect 4796 -14170 4826 -14150
rect 4796 -14210 4846 -14170
rect 4686 -14280 4846 -14210
rect 4686 -14320 4736 -14280
rect 4706 -14340 4736 -14320
rect 4796 -14320 4846 -14280
rect 4796 -14340 4826 -14320
rect 4906 -14380 4966 -14120
rect 4566 -14390 4646 -14380
rect 4566 -14450 4576 -14390
rect 4636 -14400 4646 -14390
rect 4886 -14390 4966 -14380
rect 4886 -14400 4896 -14390
rect 4636 -14450 4896 -14400
rect 4956 -14450 4966 -14390
rect 4566 -14460 4966 -14450
rect 5022 -14040 5422 -14030
rect 5022 -14100 5032 -14040
rect 5092 -14090 5352 -14040
rect 5092 -14100 5102 -14090
rect 5022 -14110 5102 -14100
rect 5342 -14100 5352 -14090
rect 5412 -14100 5422 -14040
rect 5342 -14110 5422 -14100
rect 5022 -14380 5082 -14110
rect 5352 -14120 5422 -14110
rect 5162 -14170 5192 -14150
rect 5142 -14210 5192 -14170
rect 5252 -14170 5282 -14150
rect 5252 -14210 5302 -14170
rect 5142 -14280 5302 -14210
rect 5142 -14320 5192 -14280
rect 5162 -14340 5192 -14320
rect 5252 -14320 5302 -14280
rect 5252 -14340 5282 -14320
rect 5362 -14380 5422 -14120
rect 5022 -14390 5102 -14380
rect 5022 -14450 5032 -14390
rect 5092 -14400 5102 -14390
rect 5342 -14390 5422 -14380
rect 5342 -14400 5352 -14390
rect 5092 -14450 5352 -14400
rect 5412 -14450 5422 -14390
rect 5022 -14460 5422 -14450
rect 5480 -14040 5880 -14030
rect 5480 -14100 5490 -14040
rect 5550 -14090 5810 -14040
rect 5550 -14100 5560 -14090
rect 5480 -14110 5560 -14100
rect 5800 -14100 5810 -14090
rect 5870 -14100 5880 -14040
rect 5800 -14110 5880 -14100
rect 5480 -14380 5540 -14110
rect 5810 -14120 5880 -14110
rect 5620 -14170 5650 -14150
rect 5600 -14210 5650 -14170
rect 5710 -14170 5740 -14150
rect 5710 -14210 5760 -14170
rect 5600 -14280 5760 -14210
rect 5600 -14320 5650 -14280
rect 5620 -14340 5650 -14320
rect 5710 -14320 5760 -14280
rect 5710 -14340 5740 -14320
rect 5820 -14380 5880 -14120
rect 5480 -14390 5560 -14380
rect 5480 -14450 5490 -14390
rect 5550 -14400 5560 -14390
rect 5800 -14390 5880 -14380
rect 5800 -14400 5810 -14390
rect 5550 -14450 5810 -14400
rect 5870 -14450 5880 -14390
rect 5480 -14460 5880 -14450
rect 5936 -14040 6336 -14030
rect 5936 -14100 5946 -14040
rect 6006 -14090 6266 -14040
rect 6006 -14100 6016 -14090
rect 5936 -14110 6016 -14100
rect 6256 -14100 6266 -14090
rect 6326 -14100 6336 -14040
rect 6256 -14110 6336 -14100
rect 5936 -14380 5996 -14110
rect 6266 -14120 6336 -14110
rect 6076 -14170 6106 -14150
rect 6056 -14210 6106 -14170
rect 6166 -14170 6196 -14150
rect 6166 -14210 6216 -14170
rect 6056 -14280 6216 -14210
rect 6056 -14320 6106 -14280
rect 6076 -14340 6106 -14320
rect 6166 -14320 6216 -14280
rect 6166 -14340 6196 -14320
rect 6276 -14380 6336 -14120
rect 5936 -14390 6016 -14380
rect 5936 -14450 5946 -14390
rect 6006 -14400 6016 -14390
rect 6256 -14390 6336 -14380
rect 6256 -14400 6266 -14390
rect 6006 -14450 6266 -14400
rect 6326 -14450 6336 -14390
rect 5936 -14460 6336 -14450
rect 6392 -14040 6792 -14030
rect 6392 -14100 6402 -14040
rect 6462 -14090 6722 -14040
rect 6462 -14100 6472 -14090
rect 6392 -14110 6472 -14100
rect 6712 -14100 6722 -14090
rect 6782 -14100 6792 -14040
rect 6712 -14110 6792 -14100
rect 6392 -14380 6452 -14110
rect 6722 -14120 6792 -14110
rect 6532 -14170 6562 -14150
rect 6512 -14210 6562 -14170
rect 6622 -14170 6652 -14150
rect 6622 -14210 6672 -14170
rect 6512 -14280 6672 -14210
rect 6512 -14320 6562 -14280
rect 6532 -14340 6562 -14320
rect 6622 -14320 6672 -14280
rect 6622 -14340 6652 -14320
rect 6732 -14380 6792 -14120
rect 6392 -14390 6472 -14380
rect 6392 -14450 6402 -14390
rect 6462 -14400 6472 -14390
rect 6712 -14390 6792 -14380
rect 6712 -14400 6722 -14390
rect 6462 -14450 6722 -14400
rect 6782 -14450 6792 -14390
rect 6392 -14460 6792 -14450
rect 6850 -14040 7250 -14030
rect 6850 -14100 6860 -14040
rect 6920 -14090 7180 -14040
rect 6920 -14100 6930 -14090
rect 6850 -14110 6930 -14100
rect 7170 -14100 7180 -14090
rect 7240 -14100 7250 -14040
rect 7170 -14110 7250 -14100
rect 6850 -14380 6910 -14110
rect 7180 -14120 7250 -14110
rect 6990 -14170 7020 -14150
rect 6970 -14210 7020 -14170
rect 7080 -14170 7110 -14150
rect 7080 -14210 7130 -14170
rect 6970 -14280 7130 -14210
rect 6970 -14320 7020 -14280
rect 6990 -14340 7020 -14320
rect 7080 -14320 7130 -14280
rect 7080 -14340 7110 -14320
rect 7190 -14380 7250 -14120
rect 6850 -14390 6930 -14380
rect 6850 -14450 6860 -14390
rect 6920 -14400 6930 -14390
rect 7170 -14390 7250 -14380
rect 7170 -14400 7180 -14390
rect 6920 -14450 7180 -14400
rect 7240 -14450 7250 -14390
rect 6850 -14460 7250 -14450
rect 7306 -14040 7706 -14030
rect 7306 -14100 7316 -14040
rect 7376 -14090 7636 -14040
rect 7376 -14100 7386 -14090
rect 7306 -14110 7386 -14100
rect 7626 -14100 7636 -14090
rect 7696 -14100 7706 -14040
rect 7626 -14110 7706 -14100
rect 7306 -14380 7366 -14110
rect 7636 -14120 7706 -14110
rect 7446 -14170 7476 -14150
rect 7426 -14210 7476 -14170
rect 7536 -14170 7566 -14150
rect 7536 -14210 7586 -14170
rect 7426 -14280 7586 -14210
rect 7426 -14320 7476 -14280
rect 7446 -14340 7476 -14320
rect 7536 -14320 7586 -14280
rect 7536 -14340 7566 -14320
rect 7646 -14380 7706 -14120
rect 7306 -14390 7386 -14380
rect 7306 -14450 7316 -14390
rect 7376 -14400 7386 -14390
rect 7626 -14390 7706 -14380
rect 7626 -14400 7636 -14390
rect 7376 -14450 7636 -14400
rect 7696 -14450 7706 -14390
rect 7306 -14460 7706 -14450
rect 7762 -14040 8162 -14030
rect 7762 -14100 7772 -14040
rect 7832 -14090 8092 -14040
rect 7832 -14100 7842 -14090
rect 7762 -14110 7842 -14100
rect 8082 -14100 8092 -14090
rect 8152 -14100 8162 -14040
rect 8082 -14110 8162 -14100
rect 7762 -14380 7822 -14110
rect 8092 -14120 8162 -14110
rect 7902 -14170 7932 -14150
rect 7882 -14210 7932 -14170
rect 7992 -14170 8022 -14150
rect 7992 -14210 8042 -14170
rect 7882 -14280 8042 -14210
rect 7882 -14320 7932 -14280
rect 7902 -14340 7932 -14320
rect 7992 -14320 8042 -14280
rect 7992 -14340 8022 -14320
rect 8102 -14380 8162 -14120
rect 7762 -14390 7842 -14380
rect 7762 -14450 7772 -14390
rect 7832 -14400 7842 -14390
rect 8082 -14390 8162 -14380
rect 8082 -14400 8092 -14390
rect 7832 -14450 8092 -14400
rect 8152 -14450 8162 -14390
rect 7762 -14460 8162 -14450
rect 8236 -14040 8636 -14030
rect 8236 -14100 8246 -14040
rect 8306 -14090 8566 -14040
rect 8306 -14100 8316 -14090
rect 8236 -14110 8316 -14100
rect 8556 -14100 8566 -14090
rect 8626 -14100 8636 -14040
rect 8556 -14110 8636 -14100
rect 8236 -14380 8296 -14110
rect 8566 -14120 8636 -14110
rect 8376 -14170 8406 -14150
rect 8356 -14210 8406 -14170
rect 8466 -14170 8496 -14150
rect 8466 -14210 8516 -14170
rect 8356 -14280 8516 -14210
rect 8356 -14320 8406 -14280
rect 8376 -14340 8406 -14320
rect 8466 -14320 8516 -14280
rect 8466 -14340 8496 -14320
rect 8576 -14380 8636 -14120
rect 8236 -14390 8316 -14380
rect 8236 -14450 8246 -14390
rect 8306 -14400 8316 -14390
rect 8556 -14390 8636 -14380
rect 8556 -14400 8566 -14390
rect 8306 -14450 8566 -14400
rect 8626 -14450 8636 -14390
rect 8236 -14460 8636 -14450
rect 8692 -14040 9092 -14030
rect 8692 -14100 8702 -14040
rect 8762 -14090 9022 -14040
rect 8762 -14100 8772 -14090
rect 8692 -14110 8772 -14100
rect 9012 -14100 9022 -14090
rect 9082 -14100 9092 -14040
rect 9012 -14110 9092 -14100
rect 8692 -14380 8752 -14110
rect 9022 -14120 9092 -14110
rect 8832 -14170 8862 -14150
rect 8812 -14210 8862 -14170
rect 8922 -14170 8952 -14150
rect 8922 -14210 8972 -14170
rect 8812 -14280 8972 -14210
rect 8812 -14320 8862 -14280
rect 8832 -14340 8862 -14320
rect 8922 -14320 8972 -14280
rect 8922 -14340 8952 -14320
rect 9032 -14380 9092 -14120
rect 8692 -14390 8772 -14380
rect 8692 -14450 8702 -14390
rect 8762 -14400 8772 -14390
rect 9012 -14390 9092 -14380
rect 9012 -14400 9022 -14390
rect 8762 -14450 9022 -14400
rect 9082 -14450 9092 -14390
rect 8692 -14460 9092 -14450
rect 9150 -14040 9550 -14030
rect 9150 -14100 9160 -14040
rect 9220 -14090 9480 -14040
rect 9220 -14100 9230 -14090
rect 9150 -14110 9230 -14100
rect 9470 -14100 9480 -14090
rect 9540 -14100 9550 -14040
rect 9470 -14110 9550 -14100
rect 9150 -14380 9210 -14110
rect 9480 -14120 9550 -14110
rect 9290 -14170 9320 -14150
rect 9270 -14210 9320 -14170
rect 9380 -14170 9410 -14150
rect 9380 -14210 9430 -14170
rect 9270 -14280 9430 -14210
rect 9270 -14320 9320 -14280
rect 9290 -14340 9320 -14320
rect 9380 -14320 9430 -14280
rect 9380 -14340 9410 -14320
rect 9490 -14380 9550 -14120
rect 9150 -14390 9230 -14380
rect 9150 -14450 9160 -14390
rect 9220 -14400 9230 -14390
rect 9470 -14390 9550 -14380
rect 9470 -14400 9480 -14390
rect 9220 -14450 9480 -14400
rect 9540 -14450 9550 -14390
rect 9150 -14460 9550 -14450
rect 9606 -14040 10006 -14030
rect 9606 -14100 9616 -14040
rect 9676 -14090 9936 -14040
rect 9676 -14100 9686 -14090
rect 9606 -14110 9686 -14100
rect 9926 -14100 9936 -14090
rect 9996 -14100 10006 -14040
rect 9926 -14110 10006 -14100
rect 9606 -14380 9666 -14110
rect 9936 -14120 10006 -14110
rect 9746 -14170 9776 -14150
rect 9726 -14210 9776 -14170
rect 9836 -14170 9866 -14150
rect 9836 -14210 9886 -14170
rect 9726 -14280 9886 -14210
rect 9726 -14320 9776 -14280
rect 9746 -14340 9776 -14320
rect 9836 -14320 9886 -14280
rect 9836 -14340 9866 -14320
rect 9946 -14380 10006 -14120
rect 9606 -14390 9686 -14380
rect 9606 -14450 9616 -14390
rect 9676 -14400 9686 -14390
rect 9926 -14390 10006 -14380
rect 9926 -14400 9936 -14390
rect 9676 -14450 9936 -14400
rect 9996 -14450 10006 -14390
rect 9606 -14460 10006 -14450
rect 10062 -14040 10462 -14030
rect 10062 -14100 10072 -14040
rect 10132 -14090 10392 -14040
rect 10132 -14100 10142 -14090
rect 10062 -14110 10142 -14100
rect 10382 -14100 10392 -14090
rect 10452 -14100 10462 -14040
rect 10382 -14110 10462 -14100
rect 10062 -14380 10122 -14110
rect 10392 -14120 10462 -14110
rect 10202 -14170 10232 -14150
rect 10182 -14210 10232 -14170
rect 10292 -14170 10322 -14150
rect 10292 -14210 10342 -14170
rect 10182 -14280 10342 -14210
rect 10182 -14320 10232 -14280
rect 10202 -14340 10232 -14320
rect 10292 -14320 10342 -14280
rect 10292 -14340 10322 -14320
rect 10402 -14380 10462 -14120
rect 10062 -14390 10142 -14380
rect 10062 -14450 10072 -14390
rect 10132 -14400 10142 -14390
rect 10382 -14390 10462 -14380
rect 10382 -14400 10392 -14390
rect 10132 -14450 10392 -14400
rect 10452 -14450 10462 -14390
rect 10062 -14460 10462 -14450
rect 10520 -14040 10920 -14030
rect 10520 -14100 10530 -14040
rect 10590 -14090 10850 -14040
rect 10590 -14100 10600 -14090
rect 10520 -14110 10600 -14100
rect 10840 -14100 10850 -14090
rect 10910 -14100 10920 -14040
rect 10840 -14110 10920 -14100
rect 10520 -14380 10580 -14110
rect 10850 -14120 10920 -14110
rect 10660 -14170 10690 -14150
rect 10640 -14210 10690 -14170
rect 10750 -14170 10780 -14150
rect 10750 -14210 10800 -14170
rect 10640 -14280 10800 -14210
rect 10640 -14320 10690 -14280
rect 10660 -14340 10690 -14320
rect 10750 -14320 10800 -14280
rect 10750 -14340 10780 -14320
rect 10860 -14380 10920 -14120
rect 10520 -14390 10600 -14380
rect 10520 -14450 10530 -14390
rect 10590 -14400 10600 -14390
rect 10840 -14390 10920 -14380
rect 10840 -14400 10850 -14390
rect 10590 -14450 10850 -14400
rect 10910 -14450 10920 -14390
rect 10520 -14460 10920 -14450
rect 10976 -14040 11376 -14030
rect 10976 -14100 10986 -14040
rect 11046 -14090 11306 -14040
rect 11046 -14100 11056 -14090
rect 10976 -14110 11056 -14100
rect 11296 -14100 11306 -14090
rect 11366 -14100 11376 -14040
rect 11296 -14110 11376 -14100
rect 10976 -14380 11036 -14110
rect 11306 -14120 11376 -14110
rect 11116 -14170 11146 -14150
rect 11096 -14210 11146 -14170
rect 11206 -14170 11236 -14150
rect 11206 -14210 11256 -14170
rect 11096 -14280 11256 -14210
rect 11096 -14320 11146 -14280
rect 11116 -14340 11146 -14320
rect 11206 -14320 11256 -14280
rect 11206 -14340 11236 -14320
rect 11316 -14380 11376 -14120
rect 10976 -14390 11056 -14380
rect 10976 -14450 10986 -14390
rect 11046 -14400 11056 -14390
rect 11296 -14390 11376 -14380
rect 11296 -14400 11306 -14390
rect 11046 -14450 11306 -14400
rect 11366 -14450 11376 -14390
rect 10976 -14460 11376 -14450
rect 11432 -14040 11832 -14030
rect 11432 -14100 11442 -14040
rect 11502 -14090 11762 -14040
rect 11502 -14100 11512 -14090
rect 11432 -14110 11512 -14100
rect 11752 -14100 11762 -14090
rect 11822 -14100 11832 -14040
rect 11752 -14110 11832 -14100
rect 11432 -14380 11492 -14110
rect 11762 -14120 11832 -14110
rect 11572 -14170 11602 -14150
rect 11552 -14210 11602 -14170
rect 11662 -14170 11692 -14150
rect 11662 -14210 11712 -14170
rect 11552 -14280 11712 -14210
rect 11552 -14320 11602 -14280
rect 11572 -14340 11602 -14320
rect 11662 -14320 11712 -14280
rect 11662 -14340 11692 -14320
rect 11772 -14380 11832 -14120
rect 11432 -14390 11512 -14380
rect 11432 -14450 11442 -14390
rect 11502 -14400 11512 -14390
rect 11752 -14390 11832 -14380
rect 11752 -14400 11762 -14390
rect 11502 -14450 11762 -14400
rect 11822 -14450 11832 -14390
rect 11432 -14460 11832 -14450
rect 11890 -14040 12290 -14030
rect 11890 -14100 11900 -14040
rect 11960 -14090 12220 -14040
rect 11960 -14100 11970 -14090
rect 11890 -14110 11970 -14100
rect 12210 -14100 12220 -14090
rect 12280 -14100 12290 -14040
rect 12210 -14110 12290 -14100
rect 11890 -14380 11950 -14110
rect 12220 -14120 12290 -14110
rect 12030 -14170 12060 -14150
rect 12010 -14210 12060 -14170
rect 12120 -14170 12150 -14150
rect 12120 -14210 12170 -14170
rect 12010 -14280 12170 -14210
rect 12010 -14320 12060 -14280
rect 12030 -14340 12060 -14320
rect 12120 -14320 12170 -14280
rect 12120 -14340 12150 -14320
rect 12230 -14380 12290 -14120
rect 11890 -14390 11970 -14380
rect 11890 -14450 11900 -14390
rect 11960 -14400 11970 -14390
rect 12210 -14390 12290 -14380
rect 12210 -14400 12220 -14390
rect 11960 -14450 12220 -14400
rect 12280 -14450 12290 -14390
rect 11890 -14460 12290 -14450
rect 12346 -14040 12746 -14030
rect 12346 -14100 12356 -14040
rect 12416 -14090 12676 -14040
rect 12416 -14100 12426 -14090
rect 12346 -14110 12426 -14100
rect 12666 -14100 12676 -14090
rect 12736 -14100 12746 -14040
rect 12666 -14110 12746 -14100
rect 12346 -14380 12406 -14110
rect 12676 -14120 12746 -14110
rect 12486 -14170 12516 -14150
rect 12466 -14210 12516 -14170
rect 12576 -14170 12606 -14150
rect 12576 -14210 12626 -14170
rect 12466 -14280 12626 -14210
rect 12466 -14320 12516 -14280
rect 12486 -14340 12516 -14320
rect 12576 -14320 12626 -14280
rect 12576 -14340 12606 -14320
rect 12686 -14380 12746 -14120
rect 12346 -14390 12426 -14380
rect 12346 -14450 12356 -14390
rect 12416 -14400 12426 -14390
rect 12666 -14390 12746 -14380
rect 12666 -14400 12676 -14390
rect 12416 -14450 12676 -14400
rect 12736 -14450 12746 -14390
rect 12346 -14460 12746 -14450
rect 12802 -14040 13202 -14030
rect 12802 -14100 12812 -14040
rect 12872 -14090 13132 -14040
rect 12872 -14100 12882 -14090
rect 12802 -14110 12882 -14100
rect 13122 -14100 13132 -14090
rect 13192 -14100 13202 -14040
rect 13122 -14110 13202 -14100
rect 12802 -14380 12862 -14110
rect 13132 -14120 13202 -14110
rect 12942 -14170 12972 -14150
rect 12922 -14210 12972 -14170
rect 13032 -14170 13062 -14150
rect 13032 -14210 13082 -14170
rect 12922 -14280 13082 -14210
rect 12922 -14320 12972 -14280
rect 12942 -14340 12972 -14320
rect 13032 -14320 13082 -14280
rect 13032 -14340 13062 -14320
rect 13142 -14380 13202 -14120
rect 12802 -14390 12882 -14380
rect 12802 -14450 12812 -14390
rect 12872 -14400 12882 -14390
rect 13122 -14390 13202 -14380
rect 13122 -14400 13132 -14390
rect 12872 -14450 13132 -14400
rect 13192 -14450 13202 -14390
rect 12802 -14460 13202 -14450
rect 13260 -14040 13660 -14030
rect 13260 -14100 13270 -14040
rect 13330 -14090 13590 -14040
rect 13330 -14100 13340 -14090
rect 13260 -14110 13340 -14100
rect 13580 -14100 13590 -14090
rect 13650 -14100 13660 -14040
rect 13580 -14110 13660 -14100
rect 13260 -14380 13320 -14110
rect 13590 -14120 13660 -14110
rect 13400 -14170 13430 -14150
rect 13380 -14210 13430 -14170
rect 13490 -14170 13520 -14150
rect 13490 -14210 13540 -14170
rect 13380 -14280 13540 -14210
rect 13380 -14320 13430 -14280
rect 13400 -14340 13430 -14320
rect 13490 -14320 13540 -14280
rect 13490 -14340 13520 -14320
rect 13600 -14380 13660 -14120
rect 13260 -14390 13340 -14380
rect 13260 -14450 13270 -14390
rect 13330 -14400 13340 -14390
rect 13580 -14390 13660 -14380
rect 13580 -14400 13590 -14390
rect 13330 -14450 13590 -14400
rect 13650 -14450 13660 -14390
rect 13260 -14460 13660 -14450
rect 13716 -14040 14116 -14030
rect 13716 -14100 13726 -14040
rect 13786 -14090 14046 -14040
rect 13786 -14100 13796 -14090
rect 13716 -14110 13796 -14100
rect 14036 -14100 14046 -14090
rect 14106 -14100 14116 -14040
rect 14036 -14110 14116 -14100
rect 13716 -14380 13776 -14110
rect 14046 -14120 14116 -14110
rect 13856 -14170 13886 -14150
rect 13836 -14210 13886 -14170
rect 13946 -14170 13976 -14150
rect 13946 -14210 13996 -14170
rect 13836 -14280 13996 -14210
rect 13836 -14320 13886 -14280
rect 13856 -14340 13886 -14320
rect 13946 -14320 13996 -14280
rect 13946 -14340 13976 -14320
rect 14056 -14380 14116 -14120
rect 13716 -14390 13796 -14380
rect 13716 -14450 13726 -14390
rect 13786 -14400 13796 -14390
rect 14036 -14390 14116 -14380
rect 14036 -14400 14046 -14390
rect 13786 -14450 14046 -14400
rect 14106 -14450 14116 -14390
rect 13716 -14460 14116 -14450
rect 14172 -14040 14572 -14030
rect 14172 -14100 14182 -14040
rect 14242 -14090 14502 -14040
rect 14242 -14100 14252 -14090
rect 14172 -14110 14252 -14100
rect 14492 -14100 14502 -14090
rect 14562 -14100 14572 -14040
rect 14492 -14110 14572 -14100
rect 14172 -14380 14232 -14110
rect 14502 -14120 14572 -14110
rect 14312 -14170 14342 -14150
rect 14292 -14210 14342 -14170
rect 14402 -14170 14432 -14150
rect 14402 -14210 14452 -14170
rect 14292 -14280 14452 -14210
rect 14292 -14320 14342 -14280
rect 14312 -14340 14342 -14320
rect 14402 -14320 14452 -14280
rect 14402 -14340 14432 -14320
rect 14512 -14380 14572 -14120
rect 14172 -14390 14252 -14380
rect 14172 -14450 14182 -14390
rect 14242 -14400 14252 -14390
rect 14492 -14390 14572 -14380
rect 14492 -14400 14502 -14390
rect 14242 -14450 14502 -14400
rect 14562 -14450 14572 -14390
rect 14172 -14460 14572 -14450
rect 14630 -14040 15030 -14030
rect 14630 -14100 14640 -14040
rect 14700 -14090 14960 -14040
rect 14700 -14100 14710 -14090
rect 14630 -14110 14710 -14100
rect 14950 -14100 14960 -14090
rect 15020 -14100 15030 -14040
rect 14950 -14110 15030 -14100
rect 14630 -14380 14690 -14110
rect 14960 -14120 15030 -14110
rect 14770 -14170 14800 -14150
rect 14750 -14210 14800 -14170
rect 14860 -14170 14890 -14150
rect 14860 -14210 14910 -14170
rect 14750 -14280 14910 -14210
rect 14750 -14320 14800 -14280
rect 14770 -14340 14800 -14320
rect 14860 -14320 14910 -14280
rect 14860 -14340 14890 -14320
rect 14970 -14380 15030 -14120
rect 14630 -14390 14710 -14380
rect 14630 -14450 14640 -14390
rect 14700 -14400 14710 -14390
rect 14950 -14390 15030 -14380
rect 14950 -14400 14960 -14390
rect 14700 -14450 14960 -14400
rect 15020 -14450 15030 -14390
rect 14630 -14460 15030 -14450
rect 15086 -14040 15486 -14030
rect 15086 -14100 15096 -14040
rect 15156 -14090 15416 -14040
rect 15156 -14100 15166 -14090
rect 15086 -14110 15166 -14100
rect 15406 -14100 15416 -14090
rect 15476 -14100 15486 -14040
rect 15406 -14110 15486 -14100
rect 15086 -14380 15146 -14110
rect 15416 -14120 15486 -14110
rect 15226 -14170 15256 -14150
rect 15206 -14210 15256 -14170
rect 15316 -14170 15346 -14150
rect 15316 -14210 15366 -14170
rect 15206 -14280 15366 -14210
rect 15206 -14320 15256 -14280
rect 15226 -14340 15256 -14320
rect 15316 -14320 15366 -14280
rect 15316 -14340 15346 -14320
rect 15426 -14380 15486 -14120
rect 15086 -14390 15166 -14380
rect 15086 -14450 15096 -14390
rect 15156 -14400 15166 -14390
rect 15406 -14390 15486 -14380
rect 15406 -14400 15416 -14390
rect 15156 -14450 15416 -14400
rect 15476 -14450 15486 -14390
rect 15086 -14460 15486 -14450
rect 0 -14542 400 -14532
rect 0 -14602 10 -14542
rect 70 -14592 330 -14542
rect 70 -14602 80 -14592
rect 0 -14612 80 -14602
rect 320 -14602 330 -14592
rect 390 -14602 400 -14542
rect 320 -14612 400 -14602
rect 0 -14882 60 -14612
rect 330 -14622 400 -14612
rect 140 -14672 170 -14652
rect 120 -14712 170 -14672
rect 230 -14672 260 -14652
rect 230 -14712 280 -14672
rect 120 -14782 280 -14712
rect 120 -14822 170 -14782
rect 140 -14842 170 -14822
rect 230 -14822 280 -14782
rect 230 -14842 260 -14822
rect 340 -14882 400 -14622
rect 0 -14892 80 -14882
rect 0 -14952 10 -14892
rect 70 -14902 80 -14892
rect 320 -14892 400 -14882
rect 320 -14902 330 -14892
rect 70 -14952 330 -14902
rect 390 -14952 400 -14892
rect 0 -14962 400 -14952
rect 456 -14542 856 -14532
rect 456 -14602 466 -14542
rect 526 -14592 786 -14542
rect 526 -14602 536 -14592
rect 456 -14612 536 -14602
rect 776 -14602 786 -14592
rect 846 -14602 856 -14542
rect 776 -14612 856 -14602
rect 456 -14882 516 -14612
rect 786 -14622 856 -14612
rect 596 -14672 626 -14652
rect 576 -14712 626 -14672
rect 686 -14672 716 -14652
rect 686 -14712 736 -14672
rect 576 -14782 736 -14712
rect 576 -14822 626 -14782
rect 596 -14842 626 -14822
rect 686 -14822 736 -14782
rect 686 -14842 716 -14822
rect 796 -14882 856 -14622
rect 456 -14892 536 -14882
rect 456 -14952 466 -14892
rect 526 -14902 536 -14892
rect 776 -14892 856 -14882
rect 776 -14902 786 -14892
rect 526 -14952 786 -14902
rect 846 -14952 856 -14892
rect 456 -14962 856 -14952
rect 912 -14542 1312 -14532
rect 912 -14602 922 -14542
rect 982 -14592 1242 -14542
rect 982 -14602 992 -14592
rect 912 -14612 992 -14602
rect 1232 -14602 1242 -14592
rect 1302 -14602 1312 -14542
rect 1232 -14612 1312 -14602
rect 912 -14882 972 -14612
rect 1242 -14622 1312 -14612
rect 1052 -14672 1082 -14652
rect 1032 -14712 1082 -14672
rect 1142 -14672 1172 -14652
rect 1142 -14712 1192 -14672
rect 1032 -14782 1192 -14712
rect 1032 -14822 1082 -14782
rect 1052 -14842 1082 -14822
rect 1142 -14822 1192 -14782
rect 1142 -14842 1172 -14822
rect 1252 -14882 1312 -14622
rect 912 -14892 992 -14882
rect 912 -14952 922 -14892
rect 982 -14902 992 -14892
rect 1232 -14892 1312 -14882
rect 1232 -14902 1242 -14892
rect 982 -14952 1242 -14902
rect 1302 -14952 1312 -14892
rect 912 -14962 1312 -14952
rect 1370 -14542 1770 -14532
rect 1370 -14602 1380 -14542
rect 1440 -14592 1700 -14542
rect 1440 -14602 1450 -14592
rect 1370 -14612 1450 -14602
rect 1690 -14602 1700 -14592
rect 1760 -14602 1770 -14542
rect 1690 -14612 1770 -14602
rect 1370 -14882 1430 -14612
rect 1700 -14622 1770 -14612
rect 1510 -14672 1540 -14652
rect 1490 -14712 1540 -14672
rect 1600 -14672 1630 -14652
rect 1600 -14712 1650 -14672
rect 1490 -14782 1650 -14712
rect 1490 -14822 1540 -14782
rect 1510 -14842 1540 -14822
rect 1600 -14822 1650 -14782
rect 1600 -14842 1630 -14822
rect 1710 -14882 1770 -14622
rect 1370 -14892 1450 -14882
rect 1370 -14952 1380 -14892
rect 1440 -14902 1450 -14892
rect 1690 -14892 1770 -14882
rect 1690 -14902 1700 -14892
rect 1440 -14952 1700 -14902
rect 1760 -14952 1770 -14892
rect 1370 -14962 1770 -14952
rect 1826 -14542 2226 -14532
rect 1826 -14602 1836 -14542
rect 1896 -14592 2156 -14542
rect 1896 -14602 1906 -14592
rect 1826 -14612 1906 -14602
rect 2146 -14602 2156 -14592
rect 2216 -14602 2226 -14542
rect 2146 -14612 2226 -14602
rect 1826 -14882 1886 -14612
rect 2156 -14622 2226 -14612
rect 1966 -14672 1996 -14652
rect 1946 -14712 1996 -14672
rect 2056 -14672 2086 -14652
rect 2056 -14712 2106 -14672
rect 1946 -14782 2106 -14712
rect 1946 -14822 1996 -14782
rect 1966 -14842 1996 -14822
rect 2056 -14822 2106 -14782
rect 2056 -14842 2086 -14822
rect 2166 -14882 2226 -14622
rect 1826 -14892 1906 -14882
rect 1826 -14952 1836 -14892
rect 1896 -14902 1906 -14892
rect 2146 -14892 2226 -14882
rect 2146 -14902 2156 -14892
rect 1896 -14952 2156 -14902
rect 2216 -14952 2226 -14892
rect 1826 -14962 2226 -14952
rect 2282 -14542 2682 -14532
rect 2282 -14602 2292 -14542
rect 2352 -14592 2612 -14542
rect 2352 -14602 2362 -14592
rect 2282 -14612 2362 -14602
rect 2602 -14602 2612 -14592
rect 2672 -14602 2682 -14542
rect 2602 -14612 2682 -14602
rect 2282 -14882 2342 -14612
rect 2612 -14622 2682 -14612
rect 2422 -14672 2452 -14652
rect 2402 -14712 2452 -14672
rect 2512 -14672 2542 -14652
rect 2512 -14712 2562 -14672
rect 2402 -14782 2562 -14712
rect 2402 -14822 2452 -14782
rect 2422 -14842 2452 -14822
rect 2512 -14822 2562 -14782
rect 2512 -14842 2542 -14822
rect 2622 -14882 2682 -14622
rect 2282 -14892 2362 -14882
rect 2282 -14952 2292 -14892
rect 2352 -14902 2362 -14892
rect 2602 -14892 2682 -14882
rect 2602 -14902 2612 -14892
rect 2352 -14952 2612 -14902
rect 2672 -14952 2682 -14892
rect 2282 -14962 2682 -14952
rect 2740 -14542 3140 -14532
rect 2740 -14602 2750 -14542
rect 2810 -14592 3070 -14542
rect 2810 -14602 2820 -14592
rect 2740 -14612 2820 -14602
rect 3060 -14602 3070 -14592
rect 3130 -14602 3140 -14542
rect 3060 -14612 3140 -14602
rect 2740 -14882 2800 -14612
rect 3070 -14622 3140 -14612
rect 2880 -14672 2910 -14652
rect 2860 -14712 2910 -14672
rect 2970 -14672 3000 -14652
rect 2970 -14712 3020 -14672
rect 2860 -14782 3020 -14712
rect 2860 -14822 2910 -14782
rect 2880 -14842 2910 -14822
rect 2970 -14822 3020 -14782
rect 2970 -14842 3000 -14822
rect 3080 -14882 3140 -14622
rect 2740 -14892 2820 -14882
rect 2740 -14952 2750 -14892
rect 2810 -14902 2820 -14892
rect 3060 -14892 3140 -14882
rect 3060 -14902 3070 -14892
rect 2810 -14952 3070 -14902
rect 3130 -14952 3140 -14892
rect 2740 -14962 3140 -14952
rect 3196 -14542 3596 -14532
rect 3196 -14602 3206 -14542
rect 3266 -14592 3526 -14542
rect 3266 -14602 3276 -14592
rect 3196 -14612 3276 -14602
rect 3516 -14602 3526 -14592
rect 3586 -14602 3596 -14542
rect 3516 -14612 3596 -14602
rect 3196 -14882 3256 -14612
rect 3526 -14622 3596 -14612
rect 3336 -14672 3366 -14652
rect 3316 -14712 3366 -14672
rect 3426 -14672 3456 -14652
rect 3426 -14712 3476 -14672
rect 3316 -14782 3476 -14712
rect 3316 -14822 3366 -14782
rect 3336 -14842 3366 -14822
rect 3426 -14822 3476 -14782
rect 3426 -14842 3456 -14822
rect 3536 -14882 3596 -14622
rect 3196 -14892 3276 -14882
rect 3196 -14952 3206 -14892
rect 3266 -14902 3276 -14892
rect 3516 -14892 3596 -14882
rect 3516 -14902 3526 -14892
rect 3266 -14952 3526 -14902
rect 3586 -14952 3596 -14892
rect 3196 -14962 3596 -14952
rect 3652 -14542 4052 -14532
rect 3652 -14602 3662 -14542
rect 3722 -14592 3982 -14542
rect 3722 -14602 3732 -14592
rect 3652 -14612 3732 -14602
rect 3972 -14602 3982 -14592
rect 4042 -14602 4052 -14542
rect 3972 -14612 4052 -14602
rect 3652 -14882 3712 -14612
rect 3982 -14622 4052 -14612
rect 3792 -14672 3822 -14652
rect 3772 -14712 3822 -14672
rect 3882 -14672 3912 -14652
rect 3882 -14712 3932 -14672
rect 3772 -14782 3932 -14712
rect 3772 -14822 3822 -14782
rect 3792 -14842 3822 -14822
rect 3882 -14822 3932 -14782
rect 3882 -14842 3912 -14822
rect 3992 -14882 4052 -14622
rect 3652 -14892 3732 -14882
rect 3652 -14952 3662 -14892
rect 3722 -14902 3732 -14892
rect 3972 -14892 4052 -14882
rect 3972 -14902 3982 -14892
rect 3722 -14952 3982 -14902
rect 4042 -14952 4052 -14892
rect 3652 -14962 4052 -14952
rect 4110 -14542 4510 -14532
rect 4110 -14602 4120 -14542
rect 4180 -14592 4440 -14542
rect 4180 -14602 4190 -14592
rect 4110 -14612 4190 -14602
rect 4430 -14602 4440 -14592
rect 4500 -14602 4510 -14542
rect 4430 -14612 4510 -14602
rect 4110 -14882 4170 -14612
rect 4440 -14622 4510 -14612
rect 4250 -14672 4280 -14652
rect 4230 -14712 4280 -14672
rect 4340 -14672 4370 -14652
rect 4340 -14712 4390 -14672
rect 4230 -14782 4390 -14712
rect 4230 -14822 4280 -14782
rect 4250 -14842 4280 -14822
rect 4340 -14822 4390 -14782
rect 4340 -14842 4370 -14822
rect 4450 -14882 4510 -14622
rect 4110 -14892 4190 -14882
rect 4110 -14952 4120 -14892
rect 4180 -14902 4190 -14892
rect 4430 -14892 4510 -14882
rect 4430 -14902 4440 -14892
rect 4180 -14952 4440 -14902
rect 4500 -14952 4510 -14892
rect 4110 -14962 4510 -14952
rect 4566 -14542 4966 -14532
rect 4566 -14602 4576 -14542
rect 4636 -14592 4896 -14542
rect 4636 -14602 4646 -14592
rect 4566 -14612 4646 -14602
rect 4886 -14602 4896 -14592
rect 4956 -14602 4966 -14542
rect 4886 -14612 4966 -14602
rect 4566 -14882 4626 -14612
rect 4896 -14622 4966 -14612
rect 4706 -14672 4736 -14652
rect 4686 -14712 4736 -14672
rect 4796 -14672 4826 -14652
rect 4796 -14712 4846 -14672
rect 4686 -14782 4846 -14712
rect 4686 -14822 4736 -14782
rect 4706 -14842 4736 -14822
rect 4796 -14822 4846 -14782
rect 4796 -14842 4826 -14822
rect 4906 -14882 4966 -14622
rect 4566 -14892 4646 -14882
rect 4566 -14952 4576 -14892
rect 4636 -14902 4646 -14892
rect 4886 -14892 4966 -14882
rect 4886 -14902 4896 -14892
rect 4636 -14952 4896 -14902
rect 4956 -14952 4966 -14892
rect 4566 -14962 4966 -14952
rect 5022 -14542 5422 -14532
rect 5022 -14602 5032 -14542
rect 5092 -14592 5352 -14542
rect 5092 -14602 5102 -14592
rect 5022 -14612 5102 -14602
rect 5342 -14602 5352 -14592
rect 5412 -14602 5422 -14542
rect 5342 -14612 5422 -14602
rect 5022 -14882 5082 -14612
rect 5352 -14622 5422 -14612
rect 5162 -14672 5192 -14652
rect 5142 -14712 5192 -14672
rect 5252 -14672 5282 -14652
rect 5252 -14712 5302 -14672
rect 5142 -14782 5302 -14712
rect 5142 -14822 5192 -14782
rect 5162 -14842 5192 -14822
rect 5252 -14822 5302 -14782
rect 5252 -14842 5282 -14822
rect 5362 -14882 5422 -14622
rect 5022 -14892 5102 -14882
rect 5022 -14952 5032 -14892
rect 5092 -14902 5102 -14892
rect 5342 -14892 5422 -14882
rect 5342 -14902 5352 -14892
rect 5092 -14952 5352 -14902
rect 5412 -14952 5422 -14892
rect 5022 -14962 5422 -14952
rect 5480 -14542 5880 -14532
rect 5480 -14602 5490 -14542
rect 5550 -14592 5810 -14542
rect 5550 -14602 5560 -14592
rect 5480 -14612 5560 -14602
rect 5800 -14602 5810 -14592
rect 5870 -14602 5880 -14542
rect 5800 -14612 5880 -14602
rect 5480 -14882 5540 -14612
rect 5810 -14622 5880 -14612
rect 5620 -14672 5650 -14652
rect 5600 -14712 5650 -14672
rect 5710 -14672 5740 -14652
rect 5710 -14712 5760 -14672
rect 5600 -14782 5760 -14712
rect 5600 -14822 5650 -14782
rect 5620 -14842 5650 -14822
rect 5710 -14822 5760 -14782
rect 5710 -14842 5740 -14822
rect 5820 -14882 5880 -14622
rect 5480 -14892 5560 -14882
rect 5480 -14952 5490 -14892
rect 5550 -14902 5560 -14892
rect 5800 -14892 5880 -14882
rect 5800 -14902 5810 -14892
rect 5550 -14952 5810 -14902
rect 5870 -14952 5880 -14892
rect 5480 -14962 5880 -14952
rect 5936 -14542 6336 -14532
rect 5936 -14602 5946 -14542
rect 6006 -14592 6266 -14542
rect 6006 -14602 6016 -14592
rect 5936 -14612 6016 -14602
rect 6256 -14602 6266 -14592
rect 6326 -14602 6336 -14542
rect 6256 -14612 6336 -14602
rect 5936 -14882 5996 -14612
rect 6266 -14622 6336 -14612
rect 6076 -14672 6106 -14652
rect 6056 -14712 6106 -14672
rect 6166 -14672 6196 -14652
rect 6166 -14712 6216 -14672
rect 6056 -14782 6216 -14712
rect 6056 -14822 6106 -14782
rect 6076 -14842 6106 -14822
rect 6166 -14822 6216 -14782
rect 6166 -14842 6196 -14822
rect 6276 -14882 6336 -14622
rect 5936 -14892 6016 -14882
rect 5936 -14952 5946 -14892
rect 6006 -14902 6016 -14892
rect 6256 -14892 6336 -14882
rect 6256 -14902 6266 -14892
rect 6006 -14952 6266 -14902
rect 6326 -14952 6336 -14892
rect 5936 -14962 6336 -14952
rect 6392 -14542 6792 -14532
rect 6392 -14602 6402 -14542
rect 6462 -14592 6722 -14542
rect 6462 -14602 6472 -14592
rect 6392 -14612 6472 -14602
rect 6712 -14602 6722 -14592
rect 6782 -14602 6792 -14542
rect 6712 -14612 6792 -14602
rect 6392 -14882 6452 -14612
rect 6722 -14622 6792 -14612
rect 6532 -14672 6562 -14652
rect 6512 -14712 6562 -14672
rect 6622 -14672 6652 -14652
rect 6622 -14712 6672 -14672
rect 6512 -14782 6672 -14712
rect 6512 -14822 6562 -14782
rect 6532 -14842 6562 -14822
rect 6622 -14822 6672 -14782
rect 6622 -14842 6652 -14822
rect 6732 -14882 6792 -14622
rect 6392 -14892 6472 -14882
rect 6392 -14952 6402 -14892
rect 6462 -14902 6472 -14892
rect 6712 -14892 6792 -14882
rect 6712 -14902 6722 -14892
rect 6462 -14952 6722 -14902
rect 6782 -14952 6792 -14892
rect 6392 -14962 6792 -14952
rect 6850 -14542 7250 -14532
rect 6850 -14602 6860 -14542
rect 6920 -14592 7180 -14542
rect 6920 -14602 6930 -14592
rect 6850 -14612 6930 -14602
rect 7170 -14602 7180 -14592
rect 7240 -14602 7250 -14542
rect 7170 -14612 7250 -14602
rect 6850 -14882 6910 -14612
rect 7180 -14622 7250 -14612
rect 6990 -14672 7020 -14652
rect 6970 -14712 7020 -14672
rect 7080 -14672 7110 -14652
rect 7080 -14712 7130 -14672
rect 6970 -14782 7130 -14712
rect 6970 -14822 7020 -14782
rect 6990 -14842 7020 -14822
rect 7080 -14822 7130 -14782
rect 7080 -14842 7110 -14822
rect 7190 -14882 7250 -14622
rect 6850 -14892 6930 -14882
rect 6850 -14952 6860 -14892
rect 6920 -14902 6930 -14892
rect 7170 -14892 7250 -14882
rect 7170 -14902 7180 -14892
rect 6920 -14952 7180 -14902
rect 7240 -14952 7250 -14892
rect 6850 -14962 7250 -14952
rect 7306 -14542 7706 -14532
rect 7306 -14602 7316 -14542
rect 7376 -14592 7636 -14542
rect 7376 -14602 7386 -14592
rect 7306 -14612 7386 -14602
rect 7626 -14602 7636 -14592
rect 7696 -14602 7706 -14542
rect 7626 -14612 7706 -14602
rect 7306 -14882 7366 -14612
rect 7636 -14622 7706 -14612
rect 7446 -14672 7476 -14652
rect 7426 -14712 7476 -14672
rect 7536 -14672 7566 -14652
rect 7536 -14712 7586 -14672
rect 7426 -14782 7586 -14712
rect 7426 -14822 7476 -14782
rect 7446 -14842 7476 -14822
rect 7536 -14822 7586 -14782
rect 7536 -14842 7566 -14822
rect 7646 -14882 7706 -14622
rect 7306 -14892 7386 -14882
rect 7306 -14952 7316 -14892
rect 7376 -14902 7386 -14892
rect 7626 -14892 7706 -14882
rect 7626 -14902 7636 -14892
rect 7376 -14952 7636 -14902
rect 7696 -14952 7706 -14892
rect 7306 -14962 7706 -14952
rect 7762 -14542 8162 -14532
rect 7762 -14602 7772 -14542
rect 7832 -14592 8092 -14542
rect 7832 -14602 7842 -14592
rect 7762 -14612 7842 -14602
rect 8082 -14602 8092 -14592
rect 8152 -14602 8162 -14542
rect 8082 -14612 8162 -14602
rect 7762 -14882 7822 -14612
rect 8092 -14622 8162 -14612
rect 7902 -14672 7932 -14652
rect 7882 -14712 7932 -14672
rect 7992 -14672 8022 -14652
rect 7992 -14712 8042 -14672
rect 7882 -14782 8042 -14712
rect 7882 -14822 7932 -14782
rect 7902 -14842 7932 -14822
rect 7992 -14822 8042 -14782
rect 7992 -14842 8022 -14822
rect 8102 -14882 8162 -14622
rect 7762 -14892 7842 -14882
rect 7762 -14952 7772 -14892
rect 7832 -14902 7842 -14892
rect 8082 -14892 8162 -14882
rect 8082 -14902 8092 -14892
rect 7832 -14952 8092 -14902
rect 8152 -14952 8162 -14892
rect 7762 -14962 8162 -14952
rect 8236 -14542 8636 -14532
rect 8236 -14602 8246 -14542
rect 8306 -14592 8566 -14542
rect 8306 -14602 8316 -14592
rect 8236 -14612 8316 -14602
rect 8556 -14602 8566 -14592
rect 8626 -14602 8636 -14542
rect 8556 -14612 8636 -14602
rect 8236 -14882 8296 -14612
rect 8566 -14622 8636 -14612
rect 8376 -14672 8406 -14652
rect 8356 -14712 8406 -14672
rect 8466 -14672 8496 -14652
rect 8466 -14712 8516 -14672
rect 8356 -14782 8516 -14712
rect 8356 -14822 8406 -14782
rect 8376 -14842 8406 -14822
rect 8466 -14822 8516 -14782
rect 8466 -14842 8496 -14822
rect 8576 -14882 8636 -14622
rect 8236 -14892 8316 -14882
rect 8236 -14952 8246 -14892
rect 8306 -14902 8316 -14892
rect 8556 -14892 8636 -14882
rect 8556 -14902 8566 -14892
rect 8306 -14952 8566 -14902
rect 8626 -14952 8636 -14892
rect 8236 -14962 8636 -14952
rect 8692 -14542 9092 -14532
rect 8692 -14602 8702 -14542
rect 8762 -14592 9022 -14542
rect 8762 -14602 8772 -14592
rect 8692 -14612 8772 -14602
rect 9012 -14602 9022 -14592
rect 9082 -14602 9092 -14542
rect 9012 -14612 9092 -14602
rect 8692 -14882 8752 -14612
rect 9022 -14622 9092 -14612
rect 8832 -14672 8862 -14652
rect 8812 -14712 8862 -14672
rect 8922 -14672 8952 -14652
rect 8922 -14712 8972 -14672
rect 8812 -14782 8972 -14712
rect 8812 -14822 8862 -14782
rect 8832 -14842 8862 -14822
rect 8922 -14822 8972 -14782
rect 8922 -14842 8952 -14822
rect 9032 -14882 9092 -14622
rect 8692 -14892 8772 -14882
rect 8692 -14952 8702 -14892
rect 8762 -14902 8772 -14892
rect 9012 -14892 9092 -14882
rect 9012 -14902 9022 -14892
rect 8762 -14952 9022 -14902
rect 9082 -14952 9092 -14892
rect 8692 -14962 9092 -14952
rect 9150 -14542 9550 -14532
rect 9150 -14602 9160 -14542
rect 9220 -14592 9480 -14542
rect 9220 -14602 9230 -14592
rect 9150 -14612 9230 -14602
rect 9470 -14602 9480 -14592
rect 9540 -14602 9550 -14542
rect 9470 -14612 9550 -14602
rect 9150 -14882 9210 -14612
rect 9480 -14622 9550 -14612
rect 9290 -14672 9320 -14652
rect 9270 -14712 9320 -14672
rect 9380 -14672 9410 -14652
rect 9380 -14712 9430 -14672
rect 9270 -14782 9430 -14712
rect 9270 -14822 9320 -14782
rect 9290 -14842 9320 -14822
rect 9380 -14822 9430 -14782
rect 9380 -14842 9410 -14822
rect 9490 -14882 9550 -14622
rect 9150 -14892 9230 -14882
rect 9150 -14952 9160 -14892
rect 9220 -14902 9230 -14892
rect 9470 -14892 9550 -14882
rect 9470 -14902 9480 -14892
rect 9220 -14952 9480 -14902
rect 9540 -14952 9550 -14892
rect 9150 -14962 9550 -14952
rect 9606 -14542 10006 -14532
rect 9606 -14602 9616 -14542
rect 9676 -14592 9936 -14542
rect 9676 -14602 9686 -14592
rect 9606 -14612 9686 -14602
rect 9926 -14602 9936 -14592
rect 9996 -14602 10006 -14542
rect 9926 -14612 10006 -14602
rect 9606 -14882 9666 -14612
rect 9936 -14622 10006 -14612
rect 9746 -14672 9776 -14652
rect 9726 -14712 9776 -14672
rect 9836 -14672 9866 -14652
rect 9836 -14712 9886 -14672
rect 9726 -14782 9886 -14712
rect 9726 -14822 9776 -14782
rect 9746 -14842 9776 -14822
rect 9836 -14822 9886 -14782
rect 9836 -14842 9866 -14822
rect 9946 -14882 10006 -14622
rect 9606 -14892 9686 -14882
rect 9606 -14952 9616 -14892
rect 9676 -14902 9686 -14892
rect 9926 -14892 10006 -14882
rect 9926 -14902 9936 -14892
rect 9676 -14952 9936 -14902
rect 9996 -14952 10006 -14892
rect 9606 -14962 10006 -14952
rect 10062 -14542 10462 -14532
rect 10062 -14602 10072 -14542
rect 10132 -14592 10392 -14542
rect 10132 -14602 10142 -14592
rect 10062 -14612 10142 -14602
rect 10382 -14602 10392 -14592
rect 10452 -14602 10462 -14542
rect 10382 -14612 10462 -14602
rect 10062 -14882 10122 -14612
rect 10392 -14622 10462 -14612
rect 10202 -14672 10232 -14652
rect 10182 -14712 10232 -14672
rect 10292 -14672 10322 -14652
rect 10292 -14712 10342 -14672
rect 10182 -14782 10342 -14712
rect 10182 -14822 10232 -14782
rect 10202 -14842 10232 -14822
rect 10292 -14822 10342 -14782
rect 10292 -14842 10322 -14822
rect 10402 -14882 10462 -14622
rect 10062 -14892 10142 -14882
rect 10062 -14952 10072 -14892
rect 10132 -14902 10142 -14892
rect 10382 -14892 10462 -14882
rect 10382 -14902 10392 -14892
rect 10132 -14952 10392 -14902
rect 10452 -14952 10462 -14892
rect 10062 -14962 10462 -14952
rect 10520 -14542 10920 -14532
rect 10520 -14602 10530 -14542
rect 10590 -14592 10850 -14542
rect 10590 -14602 10600 -14592
rect 10520 -14612 10600 -14602
rect 10840 -14602 10850 -14592
rect 10910 -14602 10920 -14542
rect 10840 -14612 10920 -14602
rect 10520 -14882 10580 -14612
rect 10850 -14622 10920 -14612
rect 10660 -14672 10690 -14652
rect 10640 -14712 10690 -14672
rect 10750 -14672 10780 -14652
rect 10750 -14712 10800 -14672
rect 10640 -14782 10800 -14712
rect 10640 -14822 10690 -14782
rect 10660 -14842 10690 -14822
rect 10750 -14822 10800 -14782
rect 10750 -14842 10780 -14822
rect 10860 -14882 10920 -14622
rect 10520 -14892 10600 -14882
rect 10520 -14952 10530 -14892
rect 10590 -14902 10600 -14892
rect 10840 -14892 10920 -14882
rect 10840 -14902 10850 -14892
rect 10590 -14952 10850 -14902
rect 10910 -14952 10920 -14892
rect 10520 -14962 10920 -14952
rect 10976 -14542 11376 -14532
rect 10976 -14602 10986 -14542
rect 11046 -14592 11306 -14542
rect 11046 -14602 11056 -14592
rect 10976 -14612 11056 -14602
rect 11296 -14602 11306 -14592
rect 11366 -14602 11376 -14542
rect 11296 -14612 11376 -14602
rect 10976 -14882 11036 -14612
rect 11306 -14622 11376 -14612
rect 11116 -14672 11146 -14652
rect 11096 -14712 11146 -14672
rect 11206 -14672 11236 -14652
rect 11206 -14712 11256 -14672
rect 11096 -14782 11256 -14712
rect 11096 -14822 11146 -14782
rect 11116 -14842 11146 -14822
rect 11206 -14822 11256 -14782
rect 11206 -14842 11236 -14822
rect 11316 -14882 11376 -14622
rect 10976 -14892 11056 -14882
rect 10976 -14952 10986 -14892
rect 11046 -14902 11056 -14892
rect 11296 -14892 11376 -14882
rect 11296 -14902 11306 -14892
rect 11046 -14952 11306 -14902
rect 11366 -14952 11376 -14892
rect 10976 -14962 11376 -14952
rect 11432 -14542 11832 -14532
rect 11432 -14602 11442 -14542
rect 11502 -14592 11762 -14542
rect 11502 -14602 11512 -14592
rect 11432 -14612 11512 -14602
rect 11752 -14602 11762 -14592
rect 11822 -14602 11832 -14542
rect 11752 -14612 11832 -14602
rect 11432 -14882 11492 -14612
rect 11762 -14622 11832 -14612
rect 11572 -14672 11602 -14652
rect 11552 -14712 11602 -14672
rect 11662 -14672 11692 -14652
rect 11662 -14712 11712 -14672
rect 11552 -14782 11712 -14712
rect 11552 -14822 11602 -14782
rect 11572 -14842 11602 -14822
rect 11662 -14822 11712 -14782
rect 11662 -14842 11692 -14822
rect 11772 -14882 11832 -14622
rect 11432 -14892 11512 -14882
rect 11432 -14952 11442 -14892
rect 11502 -14902 11512 -14892
rect 11752 -14892 11832 -14882
rect 11752 -14902 11762 -14892
rect 11502 -14952 11762 -14902
rect 11822 -14952 11832 -14892
rect 11432 -14962 11832 -14952
rect 11890 -14542 12290 -14532
rect 11890 -14602 11900 -14542
rect 11960 -14592 12220 -14542
rect 11960 -14602 11970 -14592
rect 11890 -14612 11970 -14602
rect 12210 -14602 12220 -14592
rect 12280 -14602 12290 -14542
rect 12210 -14612 12290 -14602
rect 11890 -14882 11950 -14612
rect 12220 -14622 12290 -14612
rect 12030 -14672 12060 -14652
rect 12010 -14712 12060 -14672
rect 12120 -14672 12150 -14652
rect 12120 -14712 12170 -14672
rect 12010 -14782 12170 -14712
rect 12010 -14822 12060 -14782
rect 12030 -14842 12060 -14822
rect 12120 -14822 12170 -14782
rect 12120 -14842 12150 -14822
rect 12230 -14882 12290 -14622
rect 11890 -14892 11970 -14882
rect 11890 -14952 11900 -14892
rect 11960 -14902 11970 -14892
rect 12210 -14892 12290 -14882
rect 12210 -14902 12220 -14892
rect 11960 -14952 12220 -14902
rect 12280 -14952 12290 -14892
rect 11890 -14962 12290 -14952
rect 12346 -14542 12746 -14532
rect 12346 -14602 12356 -14542
rect 12416 -14592 12676 -14542
rect 12416 -14602 12426 -14592
rect 12346 -14612 12426 -14602
rect 12666 -14602 12676 -14592
rect 12736 -14602 12746 -14542
rect 12666 -14612 12746 -14602
rect 12346 -14882 12406 -14612
rect 12676 -14622 12746 -14612
rect 12486 -14672 12516 -14652
rect 12466 -14712 12516 -14672
rect 12576 -14672 12606 -14652
rect 12576 -14712 12626 -14672
rect 12466 -14782 12626 -14712
rect 12466 -14822 12516 -14782
rect 12486 -14842 12516 -14822
rect 12576 -14822 12626 -14782
rect 12576 -14842 12606 -14822
rect 12686 -14882 12746 -14622
rect 12346 -14892 12426 -14882
rect 12346 -14952 12356 -14892
rect 12416 -14902 12426 -14892
rect 12666 -14892 12746 -14882
rect 12666 -14902 12676 -14892
rect 12416 -14952 12676 -14902
rect 12736 -14952 12746 -14892
rect 12346 -14962 12746 -14952
rect 12802 -14542 13202 -14532
rect 12802 -14602 12812 -14542
rect 12872 -14592 13132 -14542
rect 12872 -14602 12882 -14592
rect 12802 -14612 12882 -14602
rect 13122 -14602 13132 -14592
rect 13192 -14602 13202 -14542
rect 13122 -14612 13202 -14602
rect 12802 -14882 12862 -14612
rect 13132 -14622 13202 -14612
rect 12942 -14672 12972 -14652
rect 12922 -14712 12972 -14672
rect 13032 -14672 13062 -14652
rect 13032 -14712 13082 -14672
rect 12922 -14782 13082 -14712
rect 12922 -14822 12972 -14782
rect 12942 -14842 12972 -14822
rect 13032 -14822 13082 -14782
rect 13032 -14842 13062 -14822
rect 13142 -14882 13202 -14622
rect 12802 -14892 12882 -14882
rect 12802 -14952 12812 -14892
rect 12872 -14902 12882 -14892
rect 13122 -14892 13202 -14882
rect 13122 -14902 13132 -14892
rect 12872 -14952 13132 -14902
rect 13192 -14952 13202 -14892
rect 12802 -14962 13202 -14952
rect 13260 -14542 13660 -14532
rect 13260 -14602 13270 -14542
rect 13330 -14592 13590 -14542
rect 13330 -14602 13340 -14592
rect 13260 -14612 13340 -14602
rect 13580 -14602 13590 -14592
rect 13650 -14602 13660 -14542
rect 13580 -14612 13660 -14602
rect 13260 -14882 13320 -14612
rect 13590 -14622 13660 -14612
rect 13400 -14672 13430 -14652
rect 13380 -14712 13430 -14672
rect 13490 -14672 13520 -14652
rect 13490 -14712 13540 -14672
rect 13380 -14782 13540 -14712
rect 13380 -14822 13430 -14782
rect 13400 -14842 13430 -14822
rect 13490 -14822 13540 -14782
rect 13490 -14842 13520 -14822
rect 13600 -14882 13660 -14622
rect 13260 -14892 13340 -14882
rect 13260 -14952 13270 -14892
rect 13330 -14902 13340 -14892
rect 13580 -14892 13660 -14882
rect 13580 -14902 13590 -14892
rect 13330 -14952 13590 -14902
rect 13650 -14952 13660 -14892
rect 13260 -14962 13660 -14952
rect 13716 -14542 14116 -14532
rect 13716 -14602 13726 -14542
rect 13786 -14592 14046 -14542
rect 13786 -14602 13796 -14592
rect 13716 -14612 13796 -14602
rect 14036 -14602 14046 -14592
rect 14106 -14602 14116 -14542
rect 14036 -14612 14116 -14602
rect 13716 -14882 13776 -14612
rect 14046 -14622 14116 -14612
rect 13856 -14672 13886 -14652
rect 13836 -14712 13886 -14672
rect 13946 -14672 13976 -14652
rect 13946 -14712 13996 -14672
rect 13836 -14782 13996 -14712
rect 13836 -14822 13886 -14782
rect 13856 -14842 13886 -14822
rect 13946 -14822 13996 -14782
rect 13946 -14842 13976 -14822
rect 14056 -14882 14116 -14622
rect 13716 -14892 13796 -14882
rect 13716 -14952 13726 -14892
rect 13786 -14902 13796 -14892
rect 14036 -14892 14116 -14882
rect 14036 -14902 14046 -14892
rect 13786 -14952 14046 -14902
rect 14106 -14952 14116 -14892
rect 13716 -14962 14116 -14952
rect 14172 -14542 14572 -14532
rect 14172 -14602 14182 -14542
rect 14242 -14592 14502 -14542
rect 14242 -14602 14252 -14592
rect 14172 -14612 14252 -14602
rect 14492 -14602 14502 -14592
rect 14562 -14602 14572 -14542
rect 14492 -14612 14572 -14602
rect 14172 -14882 14232 -14612
rect 14502 -14622 14572 -14612
rect 14312 -14672 14342 -14652
rect 14292 -14712 14342 -14672
rect 14402 -14672 14432 -14652
rect 14402 -14712 14452 -14672
rect 14292 -14782 14452 -14712
rect 14292 -14822 14342 -14782
rect 14312 -14842 14342 -14822
rect 14402 -14822 14452 -14782
rect 14402 -14842 14432 -14822
rect 14512 -14882 14572 -14622
rect 14172 -14892 14252 -14882
rect 14172 -14952 14182 -14892
rect 14242 -14902 14252 -14892
rect 14492 -14892 14572 -14882
rect 14492 -14902 14502 -14892
rect 14242 -14952 14502 -14902
rect 14562 -14952 14572 -14892
rect 14172 -14962 14572 -14952
rect 14630 -14542 15030 -14532
rect 14630 -14602 14640 -14542
rect 14700 -14592 14960 -14542
rect 14700 -14602 14710 -14592
rect 14630 -14612 14710 -14602
rect 14950 -14602 14960 -14592
rect 15020 -14602 15030 -14542
rect 14950 -14612 15030 -14602
rect 14630 -14882 14690 -14612
rect 14960 -14622 15030 -14612
rect 14770 -14672 14800 -14652
rect 14750 -14712 14800 -14672
rect 14860 -14672 14890 -14652
rect 14860 -14712 14910 -14672
rect 14750 -14782 14910 -14712
rect 14750 -14822 14800 -14782
rect 14770 -14842 14800 -14822
rect 14860 -14822 14910 -14782
rect 14860 -14842 14890 -14822
rect 14970 -14882 15030 -14622
rect 14630 -14892 14710 -14882
rect 14630 -14952 14640 -14892
rect 14700 -14902 14710 -14892
rect 14950 -14892 15030 -14882
rect 14950 -14902 14960 -14892
rect 14700 -14952 14960 -14902
rect 15020 -14952 15030 -14892
rect 14630 -14962 15030 -14952
rect 15086 -14542 15486 -14532
rect 15086 -14602 15096 -14542
rect 15156 -14592 15416 -14542
rect 15156 -14602 15166 -14592
rect 15086 -14612 15166 -14602
rect 15406 -14602 15416 -14592
rect 15476 -14602 15486 -14542
rect 15406 -14612 15486 -14602
rect 15086 -14882 15146 -14612
rect 15416 -14622 15486 -14612
rect 15226 -14672 15256 -14652
rect 15206 -14712 15256 -14672
rect 15316 -14672 15346 -14652
rect 15316 -14712 15366 -14672
rect 15206 -14782 15366 -14712
rect 15206 -14822 15256 -14782
rect 15226 -14842 15256 -14822
rect 15316 -14822 15366 -14782
rect 15316 -14842 15346 -14822
rect 15426 -14882 15486 -14622
rect 15086 -14892 15166 -14882
rect 15086 -14952 15096 -14892
rect 15156 -14902 15166 -14892
rect 15406 -14892 15486 -14882
rect 15406 -14902 15416 -14892
rect 15156 -14952 15416 -14902
rect 15476 -14952 15486 -14892
rect 15086 -14962 15486 -14952
rect 0 -15034 400 -15024
rect 0 -15094 10 -15034
rect 70 -15084 330 -15034
rect 70 -15094 80 -15084
rect 0 -15104 80 -15094
rect 320 -15094 330 -15084
rect 390 -15094 400 -15034
rect 320 -15104 400 -15094
rect 0 -15374 60 -15104
rect 330 -15114 400 -15104
rect 140 -15164 170 -15144
rect 120 -15204 170 -15164
rect 230 -15164 260 -15144
rect 230 -15204 280 -15164
rect 120 -15274 280 -15204
rect 120 -15314 170 -15274
rect 140 -15334 170 -15314
rect 230 -15314 280 -15274
rect 230 -15334 260 -15314
rect 340 -15374 400 -15114
rect 0 -15384 80 -15374
rect 0 -15444 10 -15384
rect 70 -15394 80 -15384
rect 320 -15384 400 -15374
rect 320 -15394 330 -15384
rect 70 -15444 330 -15394
rect 390 -15444 400 -15384
rect 0 -15454 400 -15444
rect 456 -15034 856 -15024
rect 456 -15094 466 -15034
rect 526 -15084 786 -15034
rect 526 -15094 536 -15084
rect 456 -15104 536 -15094
rect 776 -15094 786 -15084
rect 846 -15094 856 -15034
rect 776 -15104 856 -15094
rect 456 -15374 516 -15104
rect 786 -15114 856 -15104
rect 596 -15164 626 -15144
rect 576 -15204 626 -15164
rect 686 -15164 716 -15144
rect 686 -15204 736 -15164
rect 576 -15274 736 -15204
rect 576 -15314 626 -15274
rect 596 -15334 626 -15314
rect 686 -15314 736 -15274
rect 686 -15334 716 -15314
rect 796 -15374 856 -15114
rect 456 -15384 536 -15374
rect 456 -15444 466 -15384
rect 526 -15394 536 -15384
rect 776 -15384 856 -15374
rect 776 -15394 786 -15384
rect 526 -15444 786 -15394
rect 846 -15444 856 -15384
rect 456 -15454 856 -15444
rect 912 -15034 1312 -15024
rect 912 -15094 922 -15034
rect 982 -15084 1242 -15034
rect 982 -15094 992 -15084
rect 912 -15104 992 -15094
rect 1232 -15094 1242 -15084
rect 1302 -15094 1312 -15034
rect 1232 -15104 1312 -15094
rect 912 -15374 972 -15104
rect 1242 -15114 1312 -15104
rect 1052 -15164 1082 -15144
rect 1032 -15204 1082 -15164
rect 1142 -15164 1172 -15144
rect 1142 -15204 1192 -15164
rect 1032 -15274 1192 -15204
rect 1032 -15314 1082 -15274
rect 1052 -15334 1082 -15314
rect 1142 -15314 1192 -15274
rect 1142 -15334 1172 -15314
rect 1252 -15374 1312 -15114
rect 912 -15384 992 -15374
rect 912 -15444 922 -15384
rect 982 -15394 992 -15384
rect 1232 -15384 1312 -15374
rect 1232 -15394 1242 -15384
rect 982 -15444 1242 -15394
rect 1302 -15444 1312 -15384
rect 912 -15454 1312 -15444
rect 1370 -15034 1770 -15024
rect 1370 -15094 1380 -15034
rect 1440 -15084 1700 -15034
rect 1440 -15094 1450 -15084
rect 1370 -15104 1450 -15094
rect 1690 -15094 1700 -15084
rect 1760 -15094 1770 -15034
rect 1690 -15104 1770 -15094
rect 1370 -15374 1430 -15104
rect 1700 -15114 1770 -15104
rect 1510 -15164 1540 -15144
rect 1490 -15204 1540 -15164
rect 1600 -15164 1630 -15144
rect 1600 -15204 1650 -15164
rect 1490 -15274 1650 -15204
rect 1490 -15314 1540 -15274
rect 1510 -15334 1540 -15314
rect 1600 -15314 1650 -15274
rect 1600 -15334 1630 -15314
rect 1710 -15374 1770 -15114
rect 1370 -15384 1450 -15374
rect 1370 -15444 1380 -15384
rect 1440 -15394 1450 -15384
rect 1690 -15384 1770 -15374
rect 1690 -15394 1700 -15384
rect 1440 -15444 1700 -15394
rect 1760 -15444 1770 -15384
rect 1370 -15454 1770 -15444
rect 1826 -15034 2226 -15024
rect 1826 -15094 1836 -15034
rect 1896 -15084 2156 -15034
rect 1896 -15094 1906 -15084
rect 1826 -15104 1906 -15094
rect 2146 -15094 2156 -15084
rect 2216 -15094 2226 -15034
rect 2146 -15104 2226 -15094
rect 1826 -15374 1886 -15104
rect 2156 -15114 2226 -15104
rect 1966 -15164 1996 -15144
rect 1946 -15204 1996 -15164
rect 2056 -15164 2086 -15144
rect 2056 -15204 2106 -15164
rect 1946 -15274 2106 -15204
rect 1946 -15314 1996 -15274
rect 1966 -15334 1996 -15314
rect 2056 -15314 2106 -15274
rect 2056 -15334 2086 -15314
rect 2166 -15374 2226 -15114
rect 1826 -15384 1906 -15374
rect 1826 -15444 1836 -15384
rect 1896 -15394 1906 -15384
rect 2146 -15384 2226 -15374
rect 2146 -15394 2156 -15384
rect 1896 -15444 2156 -15394
rect 2216 -15444 2226 -15384
rect 1826 -15454 2226 -15444
rect 2282 -15034 2682 -15024
rect 2282 -15094 2292 -15034
rect 2352 -15084 2612 -15034
rect 2352 -15094 2362 -15084
rect 2282 -15104 2362 -15094
rect 2602 -15094 2612 -15084
rect 2672 -15094 2682 -15034
rect 2602 -15104 2682 -15094
rect 2282 -15374 2342 -15104
rect 2612 -15114 2682 -15104
rect 2422 -15164 2452 -15144
rect 2402 -15204 2452 -15164
rect 2512 -15164 2542 -15144
rect 2512 -15204 2562 -15164
rect 2402 -15274 2562 -15204
rect 2402 -15314 2452 -15274
rect 2422 -15334 2452 -15314
rect 2512 -15314 2562 -15274
rect 2512 -15334 2542 -15314
rect 2622 -15374 2682 -15114
rect 2282 -15384 2362 -15374
rect 2282 -15444 2292 -15384
rect 2352 -15394 2362 -15384
rect 2602 -15384 2682 -15374
rect 2602 -15394 2612 -15384
rect 2352 -15444 2612 -15394
rect 2672 -15444 2682 -15384
rect 2282 -15454 2682 -15444
rect 2740 -15034 3140 -15024
rect 2740 -15094 2750 -15034
rect 2810 -15084 3070 -15034
rect 2810 -15094 2820 -15084
rect 2740 -15104 2820 -15094
rect 3060 -15094 3070 -15084
rect 3130 -15094 3140 -15034
rect 3060 -15104 3140 -15094
rect 2740 -15374 2800 -15104
rect 3070 -15114 3140 -15104
rect 2880 -15164 2910 -15144
rect 2860 -15204 2910 -15164
rect 2970 -15164 3000 -15144
rect 2970 -15204 3020 -15164
rect 2860 -15274 3020 -15204
rect 2860 -15314 2910 -15274
rect 2880 -15334 2910 -15314
rect 2970 -15314 3020 -15274
rect 2970 -15334 3000 -15314
rect 3080 -15374 3140 -15114
rect 2740 -15384 2820 -15374
rect 2740 -15444 2750 -15384
rect 2810 -15394 2820 -15384
rect 3060 -15384 3140 -15374
rect 3060 -15394 3070 -15384
rect 2810 -15444 3070 -15394
rect 3130 -15444 3140 -15384
rect 2740 -15454 3140 -15444
rect 3196 -15034 3596 -15024
rect 3196 -15094 3206 -15034
rect 3266 -15084 3526 -15034
rect 3266 -15094 3276 -15084
rect 3196 -15104 3276 -15094
rect 3516 -15094 3526 -15084
rect 3586 -15094 3596 -15034
rect 3516 -15104 3596 -15094
rect 3196 -15374 3256 -15104
rect 3526 -15114 3596 -15104
rect 3336 -15164 3366 -15144
rect 3316 -15204 3366 -15164
rect 3426 -15164 3456 -15144
rect 3426 -15204 3476 -15164
rect 3316 -15274 3476 -15204
rect 3316 -15314 3366 -15274
rect 3336 -15334 3366 -15314
rect 3426 -15314 3476 -15274
rect 3426 -15334 3456 -15314
rect 3536 -15374 3596 -15114
rect 3196 -15384 3276 -15374
rect 3196 -15444 3206 -15384
rect 3266 -15394 3276 -15384
rect 3516 -15384 3596 -15374
rect 3516 -15394 3526 -15384
rect 3266 -15444 3526 -15394
rect 3586 -15444 3596 -15384
rect 3196 -15454 3596 -15444
rect 3652 -15034 4052 -15024
rect 3652 -15094 3662 -15034
rect 3722 -15084 3982 -15034
rect 3722 -15094 3732 -15084
rect 3652 -15104 3732 -15094
rect 3972 -15094 3982 -15084
rect 4042 -15094 4052 -15034
rect 3972 -15104 4052 -15094
rect 3652 -15374 3712 -15104
rect 3982 -15114 4052 -15104
rect 3792 -15164 3822 -15144
rect 3772 -15204 3822 -15164
rect 3882 -15164 3912 -15144
rect 3882 -15204 3932 -15164
rect 3772 -15274 3932 -15204
rect 3772 -15314 3822 -15274
rect 3792 -15334 3822 -15314
rect 3882 -15314 3932 -15274
rect 3882 -15334 3912 -15314
rect 3992 -15374 4052 -15114
rect 3652 -15384 3732 -15374
rect 3652 -15444 3662 -15384
rect 3722 -15394 3732 -15384
rect 3972 -15384 4052 -15374
rect 3972 -15394 3982 -15384
rect 3722 -15444 3982 -15394
rect 4042 -15444 4052 -15384
rect 3652 -15454 4052 -15444
rect 4110 -15034 4510 -15024
rect 4110 -15094 4120 -15034
rect 4180 -15084 4440 -15034
rect 4180 -15094 4190 -15084
rect 4110 -15104 4190 -15094
rect 4430 -15094 4440 -15084
rect 4500 -15094 4510 -15034
rect 4430 -15104 4510 -15094
rect 4110 -15374 4170 -15104
rect 4440 -15114 4510 -15104
rect 4250 -15164 4280 -15144
rect 4230 -15204 4280 -15164
rect 4340 -15164 4370 -15144
rect 4340 -15204 4390 -15164
rect 4230 -15274 4390 -15204
rect 4230 -15314 4280 -15274
rect 4250 -15334 4280 -15314
rect 4340 -15314 4390 -15274
rect 4340 -15334 4370 -15314
rect 4450 -15374 4510 -15114
rect 4110 -15384 4190 -15374
rect 4110 -15444 4120 -15384
rect 4180 -15394 4190 -15384
rect 4430 -15384 4510 -15374
rect 4430 -15394 4440 -15384
rect 4180 -15444 4440 -15394
rect 4500 -15444 4510 -15384
rect 4110 -15454 4510 -15444
rect 4566 -15034 4966 -15024
rect 4566 -15094 4576 -15034
rect 4636 -15084 4896 -15034
rect 4636 -15094 4646 -15084
rect 4566 -15104 4646 -15094
rect 4886 -15094 4896 -15084
rect 4956 -15094 4966 -15034
rect 4886 -15104 4966 -15094
rect 4566 -15374 4626 -15104
rect 4896 -15114 4966 -15104
rect 4706 -15164 4736 -15144
rect 4686 -15204 4736 -15164
rect 4796 -15164 4826 -15144
rect 4796 -15204 4846 -15164
rect 4686 -15274 4846 -15204
rect 4686 -15314 4736 -15274
rect 4706 -15334 4736 -15314
rect 4796 -15314 4846 -15274
rect 4796 -15334 4826 -15314
rect 4906 -15374 4966 -15114
rect 4566 -15384 4646 -15374
rect 4566 -15444 4576 -15384
rect 4636 -15394 4646 -15384
rect 4886 -15384 4966 -15374
rect 4886 -15394 4896 -15384
rect 4636 -15444 4896 -15394
rect 4956 -15444 4966 -15384
rect 4566 -15454 4966 -15444
rect 5022 -15034 5422 -15024
rect 5022 -15094 5032 -15034
rect 5092 -15084 5352 -15034
rect 5092 -15094 5102 -15084
rect 5022 -15104 5102 -15094
rect 5342 -15094 5352 -15084
rect 5412 -15094 5422 -15034
rect 5342 -15104 5422 -15094
rect 5022 -15374 5082 -15104
rect 5352 -15114 5422 -15104
rect 5162 -15164 5192 -15144
rect 5142 -15204 5192 -15164
rect 5252 -15164 5282 -15144
rect 5252 -15204 5302 -15164
rect 5142 -15274 5302 -15204
rect 5142 -15314 5192 -15274
rect 5162 -15334 5192 -15314
rect 5252 -15314 5302 -15274
rect 5252 -15334 5282 -15314
rect 5362 -15374 5422 -15114
rect 5022 -15384 5102 -15374
rect 5022 -15444 5032 -15384
rect 5092 -15394 5102 -15384
rect 5342 -15384 5422 -15374
rect 5342 -15394 5352 -15384
rect 5092 -15444 5352 -15394
rect 5412 -15444 5422 -15384
rect 5022 -15454 5422 -15444
rect 5480 -15034 5880 -15024
rect 5480 -15094 5490 -15034
rect 5550 -15084 5810 -15034
rect 5550 -15094 5560 -15084
rect 5480 -15104 5560 -15094
rect 5800 -15094 5810 -15084
rect 5870 -15094 5880 -15034
rect 5800 -15104 5880 -15094
rect 5480 -15374 5540 -15104
rect 5810 -15114 5880 -15104
rect 5620 -15164 5650 -15144
rect 5600 -15204 5650 -15164
rect 5710 -15164 5740 -15144
rect 5710 -15204 5760 -15164
rect 5600 -15274 5760 -15204
rect 5600 -15314 5650 -15274
rect 5620 -15334 5650 -15314
rect 5710 -15314 5760 -15274
rect 5710 -15334 5740 -15314
rect 5820 -15374 5880 -15114
rect 5480 -15384 5560 -15374
rect 5480 -15444 5490 -15384
rect 5550 -15394 5560 -15384
rect 5800 -15384 5880 -15374
rect 5800 -15394 5810 -15384
rect 5550 -15444 5810 -15394
rect 5870 -15444 5880 -15384
rect 5480 -15454 5880 -15444
rect 5936 -15034 6336 -15024
rect 5936 -15094 5946 -15034
rect 6006 -15084 6266 -15034
rect 6006 -15094 6016 -15084
rect 5936 -15104 6016 -15094
rect 6256 -15094 6266 -15084
rect 6326 -15094 6336 -15034
rect 6256 -15104 6336 -15094
rect 5936 -15374 5996 -15104
rect 6266 -15114 6336 -15104
rect 6076 -15164 6106 -15144
rect 6056 -15204 6106 -15164
rect 6166 -15164 6196 -15144
rect 6166 -15204 6216 -15164
rect 6056 -15274 6216 -15204
rect 6056 -15314 6106 -15274
rect 6076 -15334 6106 -15314
rect 6166 -15314 6216 -15274
rect 6166 -15334 6196 -15314
rect 6276 -15374 6336 -15114
rect 5936 -15384 6016 -15374
rect 5936 -15444 5946 -15384
rect 6006 -15394 6016 -15384
rect 6256 -15384 6336 -15374
rect 6256 -15394 6266 -15384
rect 6006 -15444 6266 -15394
rect 6326 -15444 6336 -15384
rect 5936 -15454 6336 -15444
rect 6392 -15034 6792 -15024
rect 6392 -15094 6402 -15034
rect 6462 -15084 6722 -15034
rect 6462 -15094 6472 -15084
rect 6392 -15104 6472 -15094
rect 6712 -15094 6722 -15084
rect 6782 -15094 6792 -15034
rect 6712 -15104 6792 -15094
rect 6392 -15374 6452 -15104
rect 6722 -15114 6792 -15104
rect 6532 -15164 6562 -15144
rect 6512 -15204 6562 -15164
rect 6622 -15164 6652 -15144
rect 6622 -15204 6672 -15164
rect 6512 -15274 6672 -15204
rect 6512 -15314 6562 -15274
rect 6532 -15334 6562 -15314
rect 6622 -15314 6672 -15274
rect 6622 -15334 6652 -15314
rect 6732 -15374 6792 -15114
rect 6392 -15384 6472 -15374
rect 6392 -15444 6402 -15384
rect 6462 -15394 6472 -15384
rect 6712 -15384 6792 -15374
rect 6712 -15394 6722 -15384
rect 6462 -15444 6722 -15394
rect 6782 -15444 6792 -15384
rect 6392 -15454 6792 -15444
rect 6850 -15034 7250 -15024
rect 6850 -15094 6860 -15034
rect 6920 -15084 7180 -15034
rect 6920 -15094 6930 -15084
rect 6850 -15104 6930 -15094
rect 7170 -15094 7180 -15084
rect 7240 -15094 7250 -15034
rect 7170 -15104 7250 -15094
rect 6850 -15374 6910 -15104
rect 7180 -15114 7250 -15104
rect 6990 -15164 7020 -15144
rect 6970 -15204 7020 -15164
rect 7080 -15164 7110 -15144
rect 7080 -15204 7130 -15164
rect 6970 -15274 7130 -15204
rect 6970 -15314 7020 -15274
rect 6990 -15334 7020 -15314
rect 7080 -15314 7130 -15274
rect 7080 -15334 7110 -15314
rect 7190 -15374 7250 -15114
rect 6850 -15384 6930 -15374
rect 6850 -15444 6860 -15384
rect 6920 -15394 6930 -15384
rect 7170 -15384 7250 -15374
rect 7170 -15394 7180 -15384
rect 6920 -15444 7180 -15394
rect 7240 -15444 7250 -15384
rect 6850 -15454 7250 -15444
rect 7306 -15034 7706 -15024
rect 7306 -15094 7316 -15034
rect 7376 -15084 7636 -15034
rect 7376 -15094 7386 -15084
rect 7306 -15104 7386 -15094
rect 7626 -15094 7636 -15084
rect 7696 -15094 7706 -15034
rect 7626 -15104 7706 -15094
rect 7306 -15374 7366 -15104
rect 7636 -15114 7706 -15104
rect 7446 -15164 7476 -15144
rect 7426 -15204 7476 -15164
rect 7536 -15164 7566 -15144
rect 7536 -15204 7586 -15164
rect 7426 -15274 7586 -15204
rect 7426 -15314 7476 -15274
rect 7446 -15334 7476 -15314
rect 7536 -15314 7586 -15274
rect 7536 -15334 7566 -15314
rect 7646 -15374 7706 -15114
rect 7306 -15384 7386 -15374
rect 7306 -15444 7316 -15384
rect 7376 -15394 7386 -15384
rect 7626 -15384 7706 -15374
rect 7626 -15394 7636 -15384
rect 7376 -15444 7636 -15394
rect 7696 -15444 7706 -15384
rect 7306 -15454 7706 -15444
rect 7762 -15034 8162 -15024
rect 7762 -15094 7772 -15034
rect 7832 -15084 8092 -15034
rect 7832 -15094 7842 -15084
rect 7762 -15104 7842 -15094
rect 8082 -15094 8092 -15084
rect 8152 -15094 8162 -15034
rect 8082 -15104 8162 -15094
rect 7762 -15374 7822 -15104
rect 8092 -15114 8162 -15104
rect 7902 -15164 7932 -15144
rect 7882 -15204 7932 -15164
rect 7992 -15164 8022 -15144
rect 7992 -15204 8042 -15164
rect 7882 -15274 8042 -15204
rect 7882 -15314 7932 -15274
rect 7902 -15334 7932 -15314
rect 7992 -15314 8042 -15274
rect 7992 -15334 8022 -15314
rect 8102 -15374 8162 -15114
rect 7762 -15384 7842 -15374
rect 7762 -15444 7772 -15384
rect 7832 -15394 7842 -15384
rect 8082 -15384 8162 -15374
rect 8082 -15394 8092 -15384
rect 7832 -15444 8092 -15394
rect 8152 -15444 8162 -15384
rect 7762 -15454 8162 -15444
rect 8236 -15034 8636 -15024
rect 8236 -15094 8246 -15034
rect 8306 -15084 8566 -15034
rect 8306 -15094 8316 -15084
rect 8236 -15104 8316 -15094
rect 8556 -15094 8566 -15084
rect 8626 -15094 8636 -15034
rect 8556 -15104 8636 -15094
rect 8236 -15374 8296 -15104
rect 8566 -15114 8636 -15104
rect 8376 -15164 8406 -15144
rect 8356 -15204 8406 -15164
rect 8466 -15164 8496 -15144
rect 8466 -15204 8516 -15164
rect 8356 -15274 8516 -15204
rect 8356 -15314 8406 -15274
rect 8376 -15334 8406 -15314
rect 8466 -15314 8516 -15274
rect 8466 -15334 8496 -15314
rect 8576 -15374 8636 -15114
rect 8236 -15384 8316 -15374
rect 8236 -15444 8246 -15384
rect 8306 -15394 8316 -15384
rect 8556 -15384 8636 -15374
rect 8556 -15394 8566 -15384
rect 8306 -15444 8566 -15394
rect 8626 -15444 8636 -15384
rect 8236 -15454 8636 -15444
rect 8692 -15034 9092 -15024
rect 8692 -15094 8702 -15034
rect 8762 -15084 9022 -15034
rect 8762 -15094 8772 -15084
rect 8692 -15104 8772 -15094
rect 9012 -15094 9022 -15084
rect 9082 -15094 9092 -15034
rect 9012 -15104 9092 -15094
rect 8692 -15374 8752 -15104
rect 9022 -15114 9092 -15104
rect 8832 -15164 8862 -15144
rect 8812 -15204 8862 -15164
rect 8922 -15164 8952 -15144
rect 8922 -15204 8972 -15164
rect 8812 -15274 8972 -15204
rect 8812 -15314 8862 -15274
rect 8832 -15334 8862 -15314
rect 8922 -15314 8972 -15274
rect 8922 -15334 8952 -15314
rect 9032 -15374 9092 -15114
rect 8692 -15384 8772 -15374
rect 8692 -15444 8702 -15384
rect 8762 -15394 8772 -15384
rect 9012 -15384 9092 -15374
rect 9012 -15394 9022 -15384
rect 8762 -15444 9022 -15394
rect 9082 -15444 9092 -15384
rect 8692 -15454 9092 -15444
rect 9150 -15034 9550 -15024
rect 9150 -15094 9160 -15034
rect 9220 -15084 9480 -15034
rect 9220 -15094 9230 -15084
rect 9150 -15104 9230 -15094
rect 9470 -15094 9480 -15084
rect 9540 -15094 9550 -15034
rect 9470 -15104 9550 -15094
rect 9150 -15374 9210 -15104
rect 9480 -15114 9550 -15104
rect 9290 -15164 9320 -15144
rect 9270 -15204 9320 -15164
rect 9380 -15164 9410 -15144
rect 9380 -15204 9430 -15164
rect 9270 -15274 9430 -15204
rect 9270 -15314 9320 -15274
rect 9290 -15334 9320 -15314
rect 9380 -15314 9430 -15274
rect 9380 -15334 9410 -15314
rect 9490 -15374 9550 -15114
rect 9150 -15384 9230 -15374
rect 9150 -15444 9160 -15384
rect 9220 -15394 9230 -15384
rect 9470 -15384 9550 -15374
rect 9470 -15394 9480 -15384
rect 9220 -15444 9480 -15394
rect 9540 -15444 9550 -15384
rect 9150 -15454 9550 -15444
rect 9606 -15034 10006 -15024
rect 9606 -15094 9616 -15034
rect 9676 -15084 9936 -15034
rect 9676 -15094 9686 -15084
rect 9606 -15104 9686 -15094
rect 9926 -15094 9936 -15084
rect 9996 -15094 10006 -15034
rect 9926 -15104 10006 -15094
rect 9606 -15374 9666 -15104
rect 9936 -15114 10006 -15104
rect 9746 -15164 9776 -15144
rect 9726 -15204 9776 -15164
rect 9836 -15164 9866 -15144
rect 9836 -15204 9886 -15164
rect 9726 -15274 9886 -15204
rect 9726 -15314 9776 -15274
rect 9746 -15334 9776 -15314
rect 9836 -15314 9886 -15274
rect 9836 -15334 9866 -15314
rect 9946 -15374 10006 -15114
rect 9606 -15384 9686 -15374
rect 9606 -15444 9616 -15384
rect 9676 -15394 9686 -15384
rect 9926 -15384 10006 -15374
rect 9926 -15394 9936 -15384
rect 9676 -15444 9936 -15394
rect 9996 -15444 10006 -15384
rect 9606 -15454 10006 -15444
rect 10062 -15034 10462 -15024
rect 10062 -15094 10072 -15034
rect 10132 -15084 10392 -15034
rect 10132 -15094 10142 -15084
rect 10062 -15104 10142 -15094
rect 10382 -15094 10392 -15084
rect 10452 -15094 10462 -15034
rect 10382 -15104 10462 -15094
rect 10062 -15374 10122 -15104
rect 10392 -15114 10462 -15104
rect 10202 -15164 10232 -15144
rect 10182 -15204 10232 -15164
rect 10292 -15164 10322 -15144
rect 10292 -15204 10342 -15164
rect 10182 -15274 10342 -15204
rect 10182 -15314 10232 -15274
rect 10202 -15334 10232 -15314
rect 10292 -15314 10342 -15274
rect 10292 -15334 10322 -15314
rect 10402 -15374 10462 -15114
rect 10062 -15384 10142 -15374
rect 10062 -15444 10072 -15384
rect 10132 -15394 10142 -15384
rect 10382 -15384 10462 -15374
rect 10382 -15394 10392 -15384
rect 10132 -15444 10392 -15394
rect 10452 -15444 10462 -15384
rect 10062 -15454 10462 -15444
rect 10520 -15034 10920 -15024
rect 10520 -15094 10530 -15034
rect 10590 -15084 10850 -15034
rect 10590 -15094 10600 -15084
rect 10520 -15104 10600 -15094
rect 10840 -15094 10850 -15084
rect 10910 -15094 10920 -15034
rect 10840 -15104 10920 -15094
rect 10520 -15374 10580 -15104
rect 10850 -15114 10920 -15104
rect 10660 -15164 10690 -15144
rect 10640 -15204 10690 -15164
rect 10750 -15164 10780 -15144
rect 10750 -15204 10800 -15164
rect 10640 -15274 10800 -15204
rect 10640 -15314 10690 -15274
rect 10660 -15334 10690 -15314
rect 10750 -15314 10800 -15274
rect 10750 -15334 10780 -15314
rect 10860 -15374 10920 -15114
rect 10520 -15384 10600 -15374
rect 10520 -15444 10530 -15384
rect 10590 -15394 10600 -15384
rect 10840 -15384 10920 -15374
rect 10840 -15394 10850 -15384
rect 10590 -15444 10850 -15394
rect 10910 -15444 10920 -15384
rect 10520 -15454 10920 -15444
rect 10976 -15034 11376 -15024
rect 10976 -15094 10986 -15034
rect 11046 -15084 11306 -15034
rect 11046 -15094 11056 -15084
rect 10976 -15104 11056 -15094
rect 11296 -15094 11306 -15084
rect 11366 -15094 11376 -15034
rect 11296 -15104 11376 -15094
rect 10976 -15374 11036 -15104
rect 11306 -15114 11376 -15104
rect 11116 -15164 11146 -15144
rect 11096 -15204 11146 -15164
rect 11206 -15164 11236 -15144
rect 11206 -15204 11256 -15164
rect 11096 -15274 11256 -15204
rect 11096 -15314 11146 -15274
rect 11116 -15334 11146 -15314
rect 11206 -15314 11256 -15274
rect 11206 -15334 11236 -15314
rect 11316 -15374 11376 -15114
rect 10976 -15384 11056 -15374
rect 10976 -15444 10986 -15384
rect 11046 -15394 11056 -15384
rect 11296 -15384 11376 -15374
rect 11296 -15394 11306 -15384
rect 11046 -15444 11306 -15394
rect 11366 -15444 11376 -15384
rect 10976 -15454 11376 -15444
rect 11432 -15034 11832 -15024
rect 11432 -15094 11442 -15034
rect 11502 -15084 11762 -15034
rect 11502 -15094 11512 -15084
rect 11432 -15104 11512 -15094
rect 11752 -15094 11762 -15084
rect 11822 -15094 11832 -15034
rect 11752 -15104 11832 -15094
rect 11432 -15374 11492 -15104
rect 11762 -15114 11832 -15104
rect 11572 -15164 11602 -15144
rect 11552 -15204 11602 -15164
rect 11662 -15164 11692 -15144
rect 11662 -15204 11712 -15164
rect 11552 -15274 11712 -15204
rect 11552 -15314 11602 -15274
rect 11572 -15334 11602 -15314
rect 11662 -15314 11712 -15274
rect 11662 -15334 11692 -15314
rect 11772 -15374 11832 -15114
rect 11432 -15384 11512 -15374
rect 11432 -15444 11442 -15384
rect 11502 -15394 11512 -15384
rect 11752 -15384 11832 -15374
rect 11752 -15394 11762 -15384
rect 11502 -15444 11762 -15394
rect 11822 -15444 11832 -15384
rect 11432 -15454 11832 -15444
rect 11890 -15034 12290 -15024
rect 11890 -15094 11900 -15034
rect 11960 -15084 12220 -15034
rect 11960 -15094 11970 -15084
rect 11890 -15104 11970 -15094
rect 12210 -15094 12220 -15084
rect 12280 -15094 12290 -15034
rect 12210 -15104 12290 -15094
rect 11890 -15374 11950 -15104
rect 12220 -15114 12290 -15104
rect 12030 -15164 12060 -15144
rect 12010 -15204 12060 -15164
rect 12120 -15164 12150 -15144
rect 12120 -15204 12170 -15164
rect 12010 -15274 12170 -15204
rect 12010 -15314 12060 -15274
rect 12030 -15334 12060 -15314
rect 12120 -15314 12170 -15274
rect 12120 -15334 12150 -15314
rect 12230 -15374 12290 -15114
rect 11890 -15384 11970 -15374
rect 11890 -15444 11900 -15384
rect 11960 -15394 11970 -15384
rect 12210 -15384 12290 -15374
rect 12210 -15394 12220 -15384
rect 11960 -15444 12220 -15394
rect 12280 -15444 12290 -15384
rect 11890 -15454 12290 -15444
rect 12346 -15034 12746 -15024
rect 12346 -15094 12356 -15034
rect 12416 -15084 12676 -15034
rect 12416 -15094 12426 -15084
rect 12346 -15104 12426 -15094
rect 12666 -15094 12676 -15084
rect 12736 -15094 12746 -15034
rect 12666 -15104 12746 -15094
rect 12346 -15374 12406 -15104
rect 12676 -15114 12746 -15104
rect 12486 -15164 12516 -15144
rect 12466 -15204 12516 -15164
rect 12576 -15164 12606 -15144
rect 12576 -15204 12626 -15164
rect 12466 -15274 12626 -15204
rect 12466 -15314 12516 -15274
rect 12486 -15334 12516 -15314
rect 12576 -15314 12626 -15274
rect 12576 -15334 12606 -15314
rect 12686 -15374 12746 -15114
rect 12346 -15384 12426 -15374
rect 12346 -15444 12356 -15384
rect 12416 -15394 12426 -15384
rect 12666 -15384 12746 -15374
rect 12666 -15394 12676 -15384
rect 12416 -15444 12676 -15394
rect 12736 -15444 12746 -15384
rect 12346 -15454 12746 -15444
rect 12802 -15034 13202 -15024
rect 12802 -15094 12812 -15034
rect 12872 -15084 13132 -15034
rect 12872 -15094 12882 -15084
rect 12802 -15104 12882 -15094
rect 13122 -15094 13132 -15084
rect 13192 -15094 13202 -15034
rect 13122 -15104 13202 -15094
rect 12802 -15374 12862 -15104
rect 13132 -15114 13202 -15104
rect 12942 -15164 12972 -15144
rect 12922 -15204 12972 -15164
rect 13032 -15164 13062 -15144
rect 13032 -15204 13082 -15164
rect 12922 -15274 13082 -15204
rect 12922 -15314 12972 -15274
rect 12942 -15334 12972 -15314
rect 13032 -15314 13082 -15274
rect 13032 -15334 13062 -15314
rect 13142 -15374 13202 -15114
rect 12802 -15384 12882 -15374
rect 12802 -15444 12812 -15384
rect 12872 -15394 12882 -15384
rect 13122 -15384 13202 -15374
rect 13122 -15394 13132 -15384
rect 12872 -15444 13132 -15394
rect 13192 -15444 13202 -15384
rect 12802 -15454 13202 -15444
rect 13260 -15034 13660 -15024
rect 13260 -15094 13270 -15034
rect 13330 -15084 13590 -15034
rect 13330 -15094 13340 -15084
rect 13260 -15104 13340 -15094
rect 13580 -15094 13590 -15084
rect 13650 -15094 13660 -15034
rect 13580 -15104 13660 -15094
rect 13260 -15374 13320 -15104
rect 13590 -15114 13660 -15104
rect 13400 -15164 13430 -15144
rect 13380 -15204 13430 -15164
rect 13490 -15164 13520 -15144
rect 13490 -15204 13540 -15164
rect 13380 -15274 13540 -15204
rect 13380 -15314 13430 -15274
rect 13400 -15334 13430 -15314
rect 13490 -15314 13540 -15274
rect 13490 -15334 13520 -15314
rect 13600 -15374 13660 -15114
rect 13260 -15384 13340 -15374
rect 13260 -15444 13270 -15384
rect 13330 -15394 13340 -15384
rect 13580 -15384 13660 -15374
rect 13580 -15394 13590 -15384
rect 13330 -15444 13590 -15394
rect 13650 -15444 13660 -15384
rect 13260 -15454 13660 -15444
rect 13716 -15034 14116 -15024
rect 13716 -15094 13726 -15034
rect 13786 -15084 14046 -15034
rect 13786 -15094 13796 -15084
rect 13716 -15104 13796 -15094
rect 14036 -15094 14046 -15084
rect 14106 -15094 14116 -15034
rect 14036 -15104 14116 -15094
rect 13716 -15374 13776 -15104
rect 14046 -15114 14116 -15104
rect 13856 -15164 13886 -15144
rect 13836 -15204 13886 -15164
rect 13946 -15164 13976 -15144
rect 13946 -15204 13996 -15164
rect 13836 -15274 13996 -15204
rect 13836 -15314 13886 -15274
rect 13856 -15334 13886 -15314
rect 13946 -15314 13996 -15274
rect 13946 -15334 13976 -15314
rect 14056 -15374 14116 -15114
rect 13716 -15384 13796 -15374
rect 13716 -15444 13726 -15384
rect 13786 -15394 13796 -15384
rect 14036 -15384 14116 -15374
rect 14036 -15394 14046 -15384
rect 13786 -15444 14046 -15394
rect 14106 -15444 14116 -15384
rect 13716 -15454 14116 -15444
rect 14172 -15034 14572 -15024
rect 14172 -15094 14182 -15034
rect 14242 -15084 14502 -15034
rect 14242 -15094 14252 -15084
rect 14172 -15104 14252 -15094
rect 14492 -15094 14502 -15084
rect 14562 -15094 14572 -15034
rect 14492 -15104 14572 -15094
rect 14172 -15374 14232 -15104
rect 14502 -15114 14572 -15104
rect 14312 -15164 14342 -15144
rect 14292 -15204 14342 -15164
rect 14402 -15164 14432 -15144
rect 14402 -15204 14452 -15164
rect 14292 -15274 14452 -15204
rect 14292 -15314 14342 -15274
rect 14312 -15334 14342 -15314
rect 14402 -15314 14452 -15274
rect 14512 -15200 14572 -15114
rect 14630 -15034 15030 -15024
rect 14630 -15094 14640 -15034
rect 14700 -15084 14960 -15034
rect 14700 -15094 14710 -15084
rect 14630 -15104 14710 -15094
rect 14950 -15094 14960 -15084
rect 15020 -15094 15030 -15034
rect 14950 -15104 15030 -15094
rect 14512 -15275 14571 -15200
rect 14402 -15334 14432 -15314
rect 14512 -15374 14572 -15275
rect 14172 -15384 14252 -15374
rect 14172 -15444 14182 -15384
rect 14242 -15394 14252 -15384
rect 14492 -15384 14572 -15374
rect 14492 -15394 14502 -15384
rect 14242 -15444 14502 -15394
rect 14562 -15444 14572 -15384
rect 14172 -15454 14572 -15444
rect 14630 -15374 14690 -15104
rect 14960 -15114 15030 -15104
rect 14770 -15164 14800 -15144
rect 14750 -15204 14800 -15164
rect 14860 -15164 14890 -15144
rect 14860 -15204 14910 -15164
rect 14750 -15274 14910 -15204
rect 14750 -15314 14800 -15274
rect 14770 -15334 14800 -15314
rect 14860 -15314 14910 -15274
rect 14860 -15334 14890 -15314
rect 14970 -15374 15030 -15114
rect 14630 -15384 14710 -15374
rect 14630 -15444 14640 -15384
rect 14700 -15394 14710 -15384
rect 14950 -15384 15030 -15374
rect 14950 -15394 14960 -15384
rect 14700 -15444 14960 -15394
rect 15020 -15444 15030 -15384
rect 14630 -15454 15030 -15444
rect 15086 -15034 15486 -15024
rect 15086 -15094 15096 -15034
rect 15156 -15084 15416 -15034
rect 15156 -15094 15166 -15084
rect 15086 -15104 15166 -15094
rect 15406 -15094 15416 -15084
rect 15476 -15094 15486 -15034
rect 15406 -15104 15486 -15094
rect 15086 -15374 15146 -15104
rect 15416 -15114 15486 -15104
rect 15226 -15164 15256 -15144
rect 15206 -15204 15256 -15164
rect 15316 -15164 15346 -15144
rect 15316 -15204 15366 -15164
rect 15206 -15274 15366 -15204
rect 15206 -15314 15256 -15274
rect 15226 -15334 15256 -15314
rect 15316 -15314 15366 -15274
rect 15316 -15334 15346 -15314
rect 15426 -15374 15486 -15114
rect 15086 -15384 15166 -15374
rect 15086 -15444 15096 -15384
rect 15156 -15394 15166 -15384
rect 15406 -15384 15486 -15374
rect 15406 -15394 15416 -15384
rect 15156 -15444 15416 -15394
rect 15476 -15444 15486 -15384
rect 15086 -15454 15486 -15444
rect 0 -15550 400 -15540
rect 0 -15610 10 -15550
rect 70 -15600 330 -15550
rect 70 -15610 80 -15600
rect 0 -15620 80 -15610
rect 320 -15610 330 -15600
rect 390 -15610 400 -15550
rect 320 -15620 400 -15610
rect 0 -15890 60 -15620
rect 330 -15630 400 -15620
rect 140 -15680 170 -15660
rect 120 -15720 170 -15680
rect 230 -15680 260 -15660
rect 230 -15720 280 -15680
rect 120 -15790 280 -15720
rect 120 -15830 170 -15790
rect 140 -15850 170 -15830
rect 230 -15830 280 -15790
rect 230 -15850 260 -15830
rect 340 -15890 400 -15630
rect 0 -15900 80 -15890
rect 0 -15960 10 -15900
rect 70 -15910 80 -15900
rect 320 -15900 400 -15890
rect 320 -15910 330 -15900
rect 70 -15960 330 -15910
rect 390 -15960 400 -15900
rect 0 -15970 400 -15960
rect 456 -15550 856 -15540
rect 456 -15610 466 -15550
rect 526 -15600 786 -15550
rect 526 -15610 536 -15600
rect 456 -15620 536 -15610
rect 776 -15610 786 -15600
rect 846 -15610 856 -15550
rect 776 -15620 856 -15610
rect 456 -15890 516 -15620
rect 786 -15630 856 -15620
rect 596 -15680 626 -15660
rect 576 -15720 626 -15680
rect 686 -15680 716 -15660
rect 686 -15720 736 -15680
rect 576 -15790 736 -15720
rect 576 -15830 626 -15790
rect 596 -15850 626 -15830
rect 686 -15830 736 -15790
rect 686 -15850 716 -15830
rect 796 -15890 856 -15630
rect 456 -15900 536 -15890
rect 456 -15960 466 -15900
rect 526 -15910 536 -15900
rect 776 -15900 856 -15890
rect 776 -15910 786 -15900
rect 526 -15960 786 -15910
rect 846 -15960 856 -15900
rect 456 -15970 856 -15960
rect 912 -15550 1312 -15540
rect 912 -15610 922 -15550
rect 982 -15600 1242 -15550
rect 982 -15610 992 -15600
rect 912 -15620 992 -15610
rect 1232 -15610 1242 -15600
rect 1302 -15610 1312 -15550
rect 1232 -15620 1312 -15610
rect 912 -15890 972 -15620
rect 1242 -15630 1312 -15620
rect 1052 -15680 1082 -15660
rect 1032 -15720 1082 -15680
rect 1142 -15680 1172 -15660
rect 1142 -15720 1192 -15680
rect 1032 -15790 1192 -15720
rect 1032 -15830 1082 -15790
rect 1052 -15850 1082 -15830
rect 1142 -15830 1192 -15790
rect 1142 -15850 1172 -15830
rect 1252 -15890 1312 -15630
rect 912 -15900 992 -15890
rect 912 -15960 922 -15900
rect 982 -15910 992 -15900
rect 1232 -15900 1312 -15890
rect 1232 -15910 1242 -15900
rect 982 -15960 1242 -15910
rect 1302 -15960 1312 -15900
rect 912 -15970 1312 -15960
rect 1370 -15550 1770 -15540
rect 1370 -15610 1380 -15550
rect 1440 -15600 1700 -15550
rect 1440 -15610 1450 -15600
rect 1370 -15620 1450 -15610
rect 1690 -15610 1700 -15600
rect 1760 -15610 1770 -15550
rect 1690 -15620 1770 -15610
rect 1370 -15890 1430 -15620
rect 1700 -15630 1770 -15620
rect 1510 -15680 1540 -15660
rect 1490 -15720 1540 -15680
rect 1600 -15680 1630 -15660
rect 1600 -15720 1650 -15680
rect 1490 -15790 1650 -15720
rect 1490 -15830 1540 -15790
rect 1510 -15850 1540 -15830
rect 1600 -15830 1650 -15790
rect 1600 -15850 1630 -15830
rect 1710 -15890 1770 -15630
rect 1370 -15900 1450 -15890
rect 1370 -15960 1380 -15900
rect 1440 -15910 1450 -15900
rect 1690 -15900 1770 -15890
rect 1690 -15910 1700 -15900
rect 1440 -15960 1700 -15910
rect 1760 -15960 1770 -15900
rect 1370 -15970 1770 -15960
rect 1826 -15550 2226 -15540
rect 1826 -15610 1836 -15550
rect 1896 -15600 2156 -15550
rect 1896 -15610 1906 -15600
rect 1826 -15620 1906 -15610
rect 2146 -15610 2156 -15600
rect 2216 -15610 2226 -15550
rect 2146 -15620 2226 -15610
rect 1826 -15890 1886 -15620
rect 2156 -15630 2226 -15620
rect 1966 -15680 1996 -15660
rect 1946 -15720 1996 -15680
rect 2056 -15680 2086 -15660
rect 2056 -15720 2106 -15680
rect 1946 -15790 2106 -15720
rect 1946 -15830 1996 -15790
rect 1966 -15850 1996 -15830
rect 2056 -15830 2106 -15790
rect 2056 -15850 2086 -15830
rect 2166 -15890 2226 -15630
rect 1826 -15900 1906 -15890
rect 1826 -15960 1836 -15900
rect 1896 -15910 1906 -15900
rect 2146 -15900 2226 -15890
rect 2146 -15910 2156 -15900
rect 1896 -15960 2156 -15910
rect 2216 -15960 2226 -15900
rect 1826 -15970 2226 -15960
rect 2282 -15550 2682 -15540
rect 2282 -15610 2292 -15550
rect 2352 -15600 2612 -15550
rect 2352 -15610 2362 -15600
rect 2282 -15620 2362 -15610
rect 2602 -15610 2612 -15600
rect 2672 -15610 2682 -15550
rect 2602 -15620 2682 -15610
rect 2282 -15890 2342 -15620
rect 2612 -15630 2682 -15620
rect 2422 -15680 2452 -15660
rect 2402 -15720 2452 -15680
rect 2512 -15680 2542 -15660
rect 2512 -15720 2562 -15680
rect 2402 -15790 2562 -15720
rect 2402 -15830 2452 -15790
rect 2422 -15850 2452 -15830
rect 2512 -15830 2562 -15790
rect 2512 -15850 2542 -15830
rect 2622 -15890 2682 -15630
rect 2282 -15900 2362 -15890
rect 2282 -15960 2292 -15900
rect 2352 -15910 2362 -15900
rect 2602 -15900 2682 -15890
rect 2602 -15910 2612 -15900
rect 2352 -15960 2612 -15910
rect 2672 -15960 2682 -15900
rect 2282 -15970 2682 -15960
rect 2740 -15550 3140 -15540
rect 2740 -15610 2750 -15550
rect 2810 -15600 3070 -15550
rect 2810 -15610 2820 -15600
rect 2740 -15620 2820 -15610
rect 3060 -15610 3070 -15600
rect 3130 -15610 3140 -15550
rect 3060 -15620 3140 -15610
rect 2740 -15890 2800 -15620
rect 3070 -15630 3140 -15620
rect 2880 -15680 2910 -15660
rect 2860 -15720 2910 -15680
rect 2970 -15680 3000 -15660
rect 2970 -15720 3020 -15680
rect 2860 -15790 3020 -15720
rect 2860 -15830 2910 -15790
rect 2880 -15850 2910 -15830
rect 2970 -15830 3020 -15790
rect 2970 -15850 3000 -15830
rect 3080 -15890 3140 -15630
rect 2740 -15900 2820 -15890
rect 2740 -15960 2750 -15900
rect 2810 -15910 2820 -15900
rect 3060 -15900 3140 -15890
rect 3060 -15910 3070 -15900
rect 2810 -15960 3070 -15910
rect 3130 -15960 3140 -15900
rect 2740 -15970 3140 -15960
rect 3196 -15550 3596 -15540
rect 3196 -15610 3206 -15550
rect 3266 -15600 3526 -15550
rect 3266 -15610 3276 -15600
rect 3196 -15620 3276 -15610
rect 3516 -15610 3526 -15600
rect 3586 -15610 3596 -15550
rect 3516 -15620 3596 -15610
rect 3196 -15890 3256 -15620
rect 3526 -15630 3596 -15620
rect 3336 -15680 3366 -15660
rect 3316 -15720 3366 -15680
rect 3426 -15680 3456 -15660
rect 3426 -15720 3476 -15680
rect 3316 -15790 3476 -15720
rect 3316 -15830 3366 -15790
rect 3336 -15850 3366 -15830
rect 3426 -15830 3476 -15790
rect 3426 -15850 3456 -15830
rect 3536 -15890 3596 -15630
rect 3196 -15900 3276 -15890
rect 3196 -15960 3206 -15900
rect 3266 -15910 3276 -15900
rect 3516 -15900 3596 -15890
rect 3516 -15910 3526 -15900
rect 3266 -15960 3526 -15910
rect 3586 -15960 3596 -15900
rect 3196 -15970 3596 -15960
rect 3652 -15550 4052 -15540
rect 3652 -15610 3662 -15550
rect 3722 -15600 3982 -15550
rect 3722 -15610 3732 -15600
rect 3652 -15620 3732 -15610
rect 3972 -15610 3982 -15600
rect 4042 -15610 4052 -15550
rect 3972 -15620 4052 -15610
rect 3652 -15890 3712 -15620
rect 3982 -15630 4052 -15620
rect 3792 -15680 3822 -15660
rect 3772 -15720 3822 -15680
rect 3882 -15680 3912 -15660
rect 3882 -15720 3932 -15680
rect 3772 -15790 3932 -15720
rect 3772 -15830 3822 -15790
rect 3792 -15850 3822 -15830
rect 3882 -15830 3932 -15790
rect 3882 -15850 3912 -15830
rect 3992 -15890 4052 -15630
rect 3652 -15900 3732 -15890
rect 3652 -15960 3662 -15900
rect 3722 -15910 3732 -15900
rect 3972 -15900 4052 -15890
rect 3972 -15910 3982 -15900
rect 3722 -15960 3982 -15910
rect 4042 -15960 4052 -15900
rect 3652 -15970 4052 -15960
rect 4110 -15550 4510 -15540
rect 4110 -15610 4120 -15550
rect 4180 -15600 4440 -15550
rect 4180 -15610 4190 -15600
rect 4110 -15620 4190 -15610
rect 4430 -15610 4440 -15600
rect 4500 -15610 4510 -15550
rect 4430 -15620 4510 -15610
rect 4110 -15890 4170 -15620
rect 4440 -15630 4510 -15620
rect 4250 -15680 4280 -15660
rect 4230 -15720 4280 -15680
rect 4340 -15680 4370 -15660
rect 4340 -15720 4390 -15680
rect 4230 -15790 4390 -15720
rect 4230 -15830 4280 -15790
rect 4250 -15850 4280 -15830
rect 4340 -15830 4390 -15790
rect 4340 -15850 4370 -15830
rect 4450 -15890 4510 -15630
rect 4110 -15900 4190 -15890
rect 4110 -15960 4120 -15900
rect 4180 -15910 4190 -15900
rect 4430 -15900 4510 -15890
rect 4430 -15910 4440 -15900
rect 4180 -15960 4440 -15910
rect 4500 -15960 4510 -15900
rect 4110 -15970 4510 -15960
rect 4566 -15550 4966 -15540
rect 4566 -15610 4576 -15550
rect 4636 -15600 4896 -15550
rect 4636 -15610 4646 -15600
rect 4566 -15620 4646 -15610
rect 4886 -15610 4896 -15600
rect 4956 -15610 4966 -15550
rect 4886 -15620 4966 -15610
rect 4566 -15890 4626 -15620
rect 4896 -15630 4966 -15620
rect 4706 -15680 4736 -15660
rect 4686 -15720 4736 -15680
rect 4796 -15680 4826 -15660
rect 4796 -15720 4846 -15680
rect 4686 -15790 4846 -15720
rect 4686 -15830 4736 -15790
rect 4706 -15850 4736 -15830
rect 4796 -15830 4846 -15790
rect 4796 -15850 4826 -15830
rect 4906 -15890 4966 -15630
rect 4566 -15900 4646 -15890
rect 4566 -15960 4576 -15900
rect 4636 -15910 4646 -15900
rect 4886 -15900 4966 -15890
rect 4886 -15910 4896 -15900
rect 4636 -15960 4896 -15910
rect 4956 -15960 4966 -15900
rect 4566 -15970 4966 -15960
rect 5022 -15550 5422 -15540
rect 5022 -15610 5032 -15550
rect 5092 -15600 5352 -15550
rect 5092 -15610 5102 -15600
rect 5022 -15620 5102 -15610
rect 5342 -15610 5352 -15600
rect 5412 -15610 5422 -15550
rect 5342 -15620 5422 -15610
rect 5022 -15890 5082 -15620
rect 5352 -15630 5422 -15620
rect 5162 -15680 5192 -15660
rect 5142 -15720 5192 -15680
rect 5252 -15680 5282 -15660
rect 5252 -15720 5302 -15680
rect 5142 -15790 5302 -15720
rect 5142 -15830 5192 -15790
rect 5162 -15850 5192 -15830
rect 5252 -15830 5302 -15790
rect 5252 -15850 5282 -15830
rect 5362 -15890 5422 -15630
rect 5022 -15900 5102 -15890
rect 5022 -15960 5032 -15900
rect 5092 -15910 5102 -15900
rect 5342 -15900 5422 -15890
rect 5342 -15910 5352 -15900
rect 5092 -15960 5352 -15910
rect 5412 -15960 5422 -15900
rect 5022 -15970 5422 -15960
rect 5480 -15550 5880 -15540
rect 5480 -15610 5490 -15550
rect 5550 -15600 5810 -15550
rect 5550 -15610 5560 -15600
rect 5480 -15620 5560 -15610
rect 5800 -15610 5810 -15600
rect 5870 -15610 5880 -15550
rect 5800 -15620 5880 -15610
rect 5480 -15890 5540 -15620
rect 5810 -15630 5880 -15620
rect 5620 -15680 5650 -15660
rect 5600 -15720 5650 -15680
rect 5710 -15680 5740 -15660
rect 5710 -15720 5760 -15680
rect 5600 -15790 5760 -15720
rect 5600 -15830 5650 -15790
rect 5620 -15850 5650 -15830
rect 5710 -15830 5760 -15790
rect 5710 -15850 5740 -15830
rect 5820 -15890 5880 -15630
rect 5480 -15900 5560 -15890
rect 5480 -15960 5490 -15900
rect 5550 -15910 5560 -15900
rect 5800 -15900 5880 -15890
rect 5800 -15910 5810 -15900
rect 5550 -15960 5810 -15910
rect 5870 -15960 5880 -15900
rect 5480 -15970 5880 -15960
rect 5936 -15550 6336 -15540
rect 5936 -15610 5946 -15550
rect 6006 -15600 6266 -15550
rect 6006 -15610 6016 -15600
rect 5936 -15620 6016 -15610
rect 6256 -15610 6266 -15600
rect 6326 -15610 6336 -15550
rect 6256 -15620 6336 -15610
rect 5936 -15890 5996 -15620
rect 6266 -15630 6336 -15620
rect 6076 -15680 6106 -15660
rect 6056 -15720 6106 -15680
rect 6166 -15680 6196 -15660
rect 6166 -15720 6216 -15680
rect 6056 -15790 6216 -15720
rect 6056 -15830 6106 -15790
rect 6076 -15850 6106 -15830
rect 6166 -15830 6216 -15790
rect 6166 -15850 6196 -15830
rect 6276 -15890 6336 -15630
rect 5936 -15900 6016 -15890
rect 5936 -15960 5946 -15900
rect 6006 -15910 6016 -15900
rect 6256 -15900 6336 -15890
rect 6256 -15910 6266 -15900
rect 6006 -15960 6266 -15910
rect 6326 -15960 6336 -15900
rect 5936 -15970 6336 -15960
rect 6392 -15550 6792 -15540
rect 6392 -15610 6402 -15550
rect 6462 -15600 6722 -15550
rect 6462 -15610 6472 -15600
rect 6392 -15620 6472 -15610
rect 6712 -15610 6722 -15600
rect 6782 -15610 6792 -15550
rect 6712 -15620 6792 -15610
rect 6392 -15890 6452 -15620
rect 6722 -15630 6792 -15620
rect 6532 -15680 6562 -15660
rect 6512 -15720 6562 -15680
rect 6622 -15680 6652 -15660
rect 6622 -15720 6672 -15680
rect 6512 -15790 6672 -15720
rect 6512 -15830 6562 -15790
rect 6532 -15850 6562 -15830
rect 6622 -15830 6672 -15790
rect 6622 -15850 6652 -15830
rect 6732 -15890 6792 -15630
rect 6392 -15900 6472 -15890
rect 6392 -15960 6402 -15900
rect 6462 -15910 6472 -15900
rect 6712 -15900 6792 -15890
rect 6712 -15910 6722 -15900
rect 6462 -15960 6722 -15910
rect 6782 -15960 6792 -15900
rect 6392 -15970 6792 -15960
rect 6850 -15550 7250 -15540
rect 6850 -15610 6860 -15550
rect 6920 -15600 7180 -15550
rect 6920 -15610 6930 -15600
rect 6850 -15620 6930 -15610
rect 7170 -15610 7180 -15600
rect 7240 -15610 7250 -15550
rect 7170 -15620 7250 -15610
rect 6850 -15890 6910 -15620
rect 7180 -15630 7250 -15620
rect 6990 -15680 7020 -15660
rect 6970 -15720 7020 -15680
rect 7080 -15680 7110 -15660
rect 7080 -15720 7130 -15680
rect 6970 -15790 7130 -15720
rect 6970 -15830 7020 -15790
rect 6990 -15850 7020 -15830
rect 7080 -15830 7130 -15790
rect 7080 -15850 7110 -15830
rect 7190 -15890 7250 -15630
rect 6850 -15900 6930 -15890
rect 6850 -15960 6860 -15900
rect 6920 -15910 6930 -15900
rect 7170 -15900 7250 -15890
rect 7170 -15910 7180 -15900
rect 6920 -15960 7180 -15910
rect 7240 -15960 7250 -15900
rect 6850 -15970 7250 -15960
rect 7306 -15550 7706 -15540
rect 7306 -15610 7316 -15550
rect 7376 -15600 7636 -15550
rect 7376 -15610 7386 -15600
rect 7306 -15620 7386 -15610
rect 7626 -15610 7636 -15600
rect 7696 -15610 7706 -15550
rect 7626 -15620 7706 -15610
rect 7306 -15890 7366 -15620
rect 7636 -15630 7706 -15620
rect 7446 -15680 7476 -15660
rect 7426 -15720 7476 -15680
rect 7536 -15680 7566 -15660
rect 7536 -15720 7586 -15680
rect 7426 -15790 7586 -15720
rect 7426 -15830 7476 -15790
rect 7446 -15850 7476 -15830
rect 7536 -15830 7586 -15790
rect 7536 -15850 7566 -15830
rect 7646 -15890 7706 -15630
rect 7306 -15900 7386 -15890
rect 7306 -15960 7316 -15900
rect 7376 -15910 7386 -15900
rect 7626 -15900 7706 -15890
rect 7626 -15910 7636 -15900
rect 7376 -15960 7636 -15910
rect 7696 -15960 7706 -15900
rect 7306 -15970 7706 -15960
rect 7762 -15550 8162 -15540
rect 7762 -15610 7772 -15550
rect 7832 -15600 8092 -15550
rect 7832 -15610 7842 -15600
rect 7762 -15620 7842 -15610
rect 8082 -15610 8092 -15600
rect 8152 -15610 8162 -15550
rect 8082 -15620 8162 -15610
rect 7762 -15890 7822 -15620
rect 8092 -15630 8162 -15620
rect 7902 -15680 7932 -15660
rect 7882 -15720 7932 -15680
rect 7992 -15680 8022 -15660
rect 7992 -15720 8042 -15680
rect 7882 -15790 8042 -15720
rect 7882 -15830 7932 -15790
rect 7902 -15850 7932 -15830
rect 7992 -15830 8042 -15790
rect 7992 -15850 8022 -15830
rect 8102 -15890 8162 -15630
rect 7762 -15900 7842 -15890
rect 7762 -15960 7772 -15900
rect 7832 -15910 7842 -15900
rect 8082 -15900 8162 -15890
rect 8082 -15910 8092 -15900
rect 7832 -15960 8092 -15910
rect 8152 -15960 8162 -15900
rect 7762 -15970 8162 -15960
rect 8236 -15550 8636 -15540
rect 8236 -15610 8246 -15550
rect 8306 -15600 8566 -15550
rect 8306 -15610 8316 -15600
rect 8236 -15620 8316 -15610
rect 8556 -15610 8566 -15600
rect 8626 -15610 8636 -15550
rect 8556 -15620 8636 -15610
rect 8236 -15890 8296 -15620
rect 8566 -15630 8636 -15620
rect 8376 -15680 8406 -15660
rect 8356 -15720 8406 -15680
rect 8466 -15680 8496 -15660
rect 8466 -15720 8516 -15680
rect 8356 -15790 8516 -15720
rect 8356 -15830 8406 -15790
rect 8376 -15850 8406 -15830
rect 8466 -15830 8516 -15790
rect 8466 -15850 8496 -15830
rect 8576 -15890 8636 -15630
rect 8236 -15900 8316 -15890
rect 8236 -15960 8246 -15900
rect 8306 -15910 8316 -15900
rect 8556 -15900 8636 -15890
rect 8556 -15910 8566 -15900
rect 8306 -15960 8566 -15910
rect 8626 -15960 8636 -15900
rect 8236 -15970 8636 -15960
rect 8692 -15550 9092 -15540
rect 8692 -15610 8702 -15550
rect 8762 -15600 9022 -15550
rect 8762 -15610 8772 -15600
rect 8692 -15620 8772 -15610
rect 9012 -15610 9022 -15600
rect 9082 -15610 9092 -15550
rect 9012 -15620 9092 -15610
rect 8692 -15890 8752 -15620
rect 9022 -15630 9092 -15620
rect 8832 -15680 8862 -15660
rect 8812 -15720 8862 -15680
rect 8922 -15680 8952 -15660
rect 8922 -15720 8972 -15680
rect 8812 -15790 8972 -15720
rect 8812 -15830 8862 -15790
rect 8832 -15850 8862 -15830
rect 8922 -15830 8972 -15790
rect 8922 -15850 8952 -15830
rect 9032 -15890 9092 -15630
rect 8692 -15900 8772 -15890
rect 8692 -15960 8702 -15900
rect 8762 -15910 8772 -15900
rect 9012 -15900 9092 -15890
rect 9012 -15910 9022 -15900
rect 8762 -15960 9022 -15910
rect 9082 -15960 9092 -15900
rect 8692 -15970 9092 -15960
rect 9150 -15550 9550 -15540
rect 9150 -15610 9160 -15550
rect 9220 -15600 9480 -15550
rect 9220 -15610 9230 -15600
rect 9150 -15620 9230 -15610
rect 9470 -15610 9480 -15600
rect 9540 -15610 9550 -15550
rect 9470 -15620 9550 -15610
rect 9150 -15890 9210 -15620
rect 9480 -15630 9550 -15620
rect 9290 -15680 9320 -15660
rect 9270 -15720 9320 -15680
rect 9380 -15680 9410 -15660
rect 9380 -15720 9430 -15680
rect 9270 -15790 9430 -15720
rect 9270 -15830 9320 -15790
rect 9290 -15850 9320 -15830
rect 9380 -15830 9430 -15790
rect 9380 -15850 9410 -15830
rect 9490 -15890 9550 -15630
rect 9150 -15900 9230 -15890
rect 9150 -15960 9160 -15900
rect 9220 -15910 9230 -15900
rect 9470 -15900 9550 -15890
rect 9470 -15910 9480 -15900
rect 9220 -15960 9480 -15910
rect 9540 -15960 9550 -15900
rect 9150 -15970 9550 -15960
rect 9606 -15550 10006 -15540
rect 9606 -15610 9616 -15550
rect 9676 -15600 9936 -15550
rect 9676 -15610 9686 -15600
rect 9606 -15620 9686 -15610
rect 9926 -15610 9936 -15600
rect 9996 -15610 10006 -15550
rect 9926 -15620 10006 -15610
rect 9606 -15890 9666 -15620
rect 9936 -15630 10006 -15620
rect 9746 -15680 9776 -15660
rect 9726 -15720 9776 -15680
rect 9836 -15680 9866 -15660
rect 9836 -15720 9886 -15680
rect 9726 -15790 9886 -15720
rect 9726 -15830 9776 -15790
rect 9746 -15850 9776 -15830
rect 9836 -15830 9886 -15790
rect 9836 -15850 9866 -15830
rect 9946 -15890 10006 -15630
rect 9606 -15900 9686 -15890
rect 9606 -15960 9616 -15900
rect 9676 -15910 9686 -15900
rect 9926 -15900 10006 -15890
rect 9926 -15910 9936 -15900
rect 9676 -15960 9936 -15910
rect 9996 -15960 10006 -15900
rect 9606 -15970 10006 -15960
rect 10062 -15550 10462 -15540
rect 10062 -15610 10072 -15550
rect 10132 -15600 10392 -15550
rect 10132 -15610 10142 -15600
rect 10062 -15620 10142 -15610
rect 10382 -15610 10392 -15600
rect 10452 -15610 10462 -15550
rect 10382 -15620 10462 -15610
rect 10062 -15890 10122 -15620
rect 10392 -15630 10462 -15620
rect 10202 -15680 10232 -15660
rect 10182 -15720 10232 -15680
rect 10292 -15680 10322 -15660
rect 10292 -15720 10342 -15680
rect 10182 -15790 10342 -15720
rect 10182 -15830 10232 -15790
rect 10202 -15850 10232 -15830
rect 10292 -15830 10342 -15790
rect 10292 -15850 10322 -15830
rect 10402 -15890 10462 -15630
rect 10062 -15900 10142 -15890
rect 10062 -15960 10072 -15900
rect 10132 -15910 10142 -15900
rect 10382 -15900 10462 -15890
rect 10382 -15910 10392 -15900
rect 10132 -15960 10392 -15910
rect 10452 -15960 10462 -15900
rect 10062 -15970 10462 -15960
rect 10520 -15550 10920 -15540
rect 10520 -15610 10530 -15550
rect 10590 -15600 10850 -15550
rect 10590 -15610 10600 -15600
rect 10520 -15620 10600 -15610
rect 10840 -15610 10850 -15600
rect 10910 -15610 10920 -15550
rect 10840 -15620 10920 -15610
rect 10520 -15890 10580 -15620
rect 10850 -15630 10920 -15620
rect 10660 -15680 10690 -15660
rect 10640 -15720 10690 -15680
rect 10750 -15680 10780 -15660
rect 10750 -15720 10800 -15680
rect 10640 -15790 10800 -15720
rect 10640 -15830 10690 -15790
rect 10660 -15850 10690 -15830
rect 10750 -15830 10800 -15790
rect 10750 -15850 10780 -15830
rect 10860 -15890 10920 -15630
rect 10520 -15900 10600 -15890
rect 10520 -15960 10530 -15900
rect 10590 -15910 10600 -15900
rect 10840 -15900 10920 -15890
rect 10840 -15910 10850 -15900
rect 10590 -15960 10850 -15910
rect 10910 -15960 10920 -15900
rect 10520 -15970 10920 -15960
rect 10976 -15550 11376 -15540
rect 10976 -15610 10986 -15550
rect 11046 -15600 11306 -15550
rect 11046 -15610 11056 -15600
rect 10976 -15620 11056 -15610
rect 11296 -15610 11306 -15600
rect 11366 -15610 11376 -15550
rect 11296 -15620 11376 -15610
rect 10976 -15890 11036 -15620
rect 11306 -15630 11376 -15620
rect 11116 -15680 11146 -15660
rect 11096 -15720 11146 -15680
rect 11206 -15680 11236 -15660
rect 11206 -15720 11256 -15680
rect 11096 -15790 11256 -15720
rect 11096 -15830 11146 -15790
rect 11116 -15850 11146 -15830
rect 11206 -15830 11256 -15790
rect 11206 -15850 11236 -15830
rect 11316 -15890 11376 -15630
rect 10976 -15900 11056 -15890
rect 10976 -15960 10986 -15900
rect 11046 -15910 11056 -15900
rect 11296 -15900 11376 -15890
rect 11296 -15910 11306 -15900
rect 11046 -15960 11306 -15910
rect 11366 -15960 11376 -15900
rect 10976 -15970 11376 -15960
rect 11432 -15550 11832 -15540
rect 11432 -15610 11442 -15550
rect 11502 -15600 11762 -15550
rect 11502 -15610 11512 -15600
rect 11432 -15620 11512 -15610
rect 11752 -15610 11762 -15600
rect 11822 -15610 11832 -15550
rect 11752 -15620 11832 -15610
rect 11432 -15890 11492 -15620
rect 11762 -15630 11832 -15620
rect 11572 -15680 11602 -15660
rect 11552 -15720 11602 -15680
rect 11662 -15680 11692 -15660
rect 11662 -15720 11712 -15680
rect 11552 -15790 11712 -15720
rect 11552 -15830 11602 -15790
rect 11572 -15850 11602 -15830
rect 11662 -15830 11712 -15790
rect 11662 -15850 11692 -15830
rect 11772 -15890 11832 -15630
rect 11432 -15900 11512 -15890
rect 11432 -15960 11442 -15900
rect 11502 -15910 11512 -15900
rect 11752 -15900 11832 -15890
rect 11752 -15910 11762 -15900
rect 11502 -15960 11762 -15910
rect 11822 -15960 11832 -15900
rect 11432 -15970 11832 -15960
rect 11890 -15550 12290 -15540
rect 11890 -15610 11900 -15550
rect 11960 -15600 12220 -15550
rect 11960 -15610 11970 -15600
rect 11890 -15620 11970 -15610
rect 12210 -15610 12220 -15600
rect 12280 -15610 12290 -15550
rect 12210 -15620 12290 -15610
rect 11890 -15890 11950 -15620
rect 12220 -15630 12290 -15620
rect 12030 -15680 12060 -15660
rect 12010 -15720 12060 -15680
rect 12120 -15680 12150 -15660
rect 12120 -15720 12170 -15680
rect 12010 -15790 12170 -15720
rect 12010 -15830 12060 -15790
rect 12030 -15850 12060 -15830
rect 12120 -15830 12170 -15790
rect 12120 -15850 12150 -15830
rect 12230 -15890 12290 -15630
rect 11890 -15900 11970 -15890
rect 11890 -15960 11900 -15900
rect 11960 -15910 11970 -15900
rect 12210 -15900 12290 -15890
rect 12210 -15910 12220 -15900
rect 11960 -15960 12220 -15910
rect 12280 -15960 12290 -15900
rect 11890 -15970 12290 -15960
rect 12346 -15550 12746 -15540
rect 12346 -15610 12356 -15550
rect 12416 -15600 12676 -15550
rect 12416 -15610 12426 -15600
rect 12346 -15620 12426 -15610
rect 12666 -15610 12676 -15600
rect 12736 -15610 12746 -15550
rect 12666 -15620 12746 -15610
rect 12346 -15890 12406 -15620
rect 12676 -15630 12746 -15620
rect 12486 -15680 12516 -15660
rect 12466 -15720 12516 -15680
rect 12576 -15680 12606 -15660
rect 12576 -15720 12626 -15680
rect 12466 -15790 12626 -15720
rect 12466 -15830 12516 -15790
rect 12486 -15850 12516 -15830
rect 12576 -15830 12626 -15790
rect 12576 -15850 12606 -15830
rect 12686 -15890 12746 -15630
rect 12346 -15900 12426 -15890
rect 12346 -15960 12356 -15900
rect 12416 -15910 12426 -15900
rect 12666 -15900 12746 -15890
rect 12666 -15910 12676 -15900
rect 12416 -15960 12676 -15910
rect 12736 -15960 12746 -15900
rect 12346 -15970 12746 -15960
rect 12802 -15550 13202 -15540
rect 12802 -15610 12812 -15550
rect 12872 -15600 13132 -15550
rect 12872 -15610 12882 -15600
rect 12802 -15620 12882 -15610
rect 13122 -15610 13132 -15600
rect 13192 -15610 13202 -15550
rect 13122 -15620 13202 -15610
rect 12802 -15890 12862 -15620
rect 13132 -15630 13202 -15620
rect 12942 -15680 12972 -15660
rect 12922 -15720 12972 -15680
rect 13032 -15680 13062 -15660
rect 13032 -15720 13082 -15680
rect 12922 -15790 13082 -15720
rect 12922 -15830 12972 -15790
rect 12942 -15850 12972 -15830
rect 13032 -15830 13082 -15790
rect 13032 -15850 13062 -15830
rect 13142 -15890 13202 -15630
rect 12802 -15900 12882 -15890
rect 12802 -15960 12812 -15900
rect 12872 -15910 12882 -15900
rect 13122 -15900 13202 -15890
rect 13122 -15910 13132 -15900
rect 12872 -15960 13132 -15910
rect 13192 -15960 13202 -15900
rect 12802 -15970 13202 -15960
rect 13260 -15550 13660 -15540
rect 13260 -15610 13270 -15550
rect 13330 -15600 13590 -15550
rect 13330 -15610 13340 -15600
rect 13260 -15620 13340 -15610
rect 13580 -15610 13590 -15600
rect 13650 -15610 13660 -15550
rect 13580 -15620 13660 -15610
rect 13260 -15890 13320 -15620
rect 13590 -15630 13660 -15620
rect 13400 -15680 13430 -15660
rect 13380 -15720 13430 -15680
rect 13490 -15680 13520 -15660
rect 13490 -15720 13540 -15680
rect 13380 -15790 13540 -15720
rect 13380 -15830 13430 -15790
rect 13400 -15850 13430 -15830
rect 13490 -15830 13540 -15790
rect 13490 -15850 13520 -15830
rect 13600 -15890 13660 -15630
rect 13260 -15900 13340 -15890
rect 13260 -15960 13270 -15900
rect 13330 -15910 13340 -15900
rect 13580 -15900 13660 -15890
rect 13580 -15910 13590 -15900
rect 13330 -15960 13590 -15910
rect 13650 -15960 13660 -15900
rect 13260 -15970 13660 -15960
rect 13716 -15550 14116 -15540
rect 13716 -15610 13726 -15550
rect 13786 -15600 14046 -15550
rect 13786 -15610 13796 -15600
rect 13716 -15620 13796 -15610
rect 14036 -15610 14046 -15600
rect 14106 -15610 14116 -15550
rect 14036 -15620 14116 -15610
rect 13716 -15890 13776 -15620
rect 14046 -15630 14116 -15620
rect 13856 -15680 13886 -15660
rect 13836 -15720 13886 -15680
rect 13946 -15680 13976 -15660
rect 13946 -15720 13996 -15680
rect 13836 -15790 13996 -15720
rect 13836 -15830 13886 -15790
rect 13856 -15850 13886 -15830
rect 13946 -15830 13996 -15790
rect 13946 -15850 13976 -15830
rect 14056 -15890 14116 -15630
rect 13716 -15900 13796 -15890
rect 13716 -15960 13726 -15900
rect 13786 -15910 13796 -15900
rect 14036 -15900 14116 -15890
rect 14036 -15910 14046 -15900
rect 13786 -15960 14046 -15910
rect 14106 -15960 14116 -15900
rect 13716 -15970 14116 -15960
rect 14172 -15550 14572 -15540
rect 14172 -15610 14182 -15550
rect 14242 -15600 14502 -15550
rect 14242 -15610 14252 -15600
rect 14172 -15620 14252 -15610
rect 14492 -15610 14502 -15600
rect 14562 -15610 14572 -15550
rect 14492 -15620 14572 -15610
rect 14172 -15890 14232 -15620
rect 14502 -15630 14572 -15620
rect 14312 -15680 14342 -15660
rect 14292 -15720 14342 -15680
rect 14402 -15680 14432 -15660
rect 14402 -15720 14452 -15680
rect 14292 -15790 14452 -15720
rect 14292 -15830 14342 -15790
rect 14312 -15850 14342 -15830
rect 14402 -15830 14452 -15790
rect 14402 -15850 14432 -15830
rect 14512 -15890 14572 -15630
rect 14172 -15900 14252 -15890
rect 14172 -15960 14182 -15900
rect 14242 -15910 14252 -15900
rect 14492 -15900 14572 -15890
rect 14492 -15910 14502 -15900
rect 14242 -15960 14502 -15910
rect 14562 -15960 14572 -15900
rect 14172 -15970 14572 -15960
rect 14630 -15550 15030 -15540
rect 14630 -15610 14640 -15550
rect 14700 -15600 14960 -15550
rect 14700 -15610 14710 -15600
rect 14630 -15620 14710 -15610
rect 14950 -15610 14960 -15600
rect 15020 -15610 15030 -15550
rect 14950 -15620 15030 -15610
rect 14630 -15890 14690 -15620
rect 14960 -15630 15030 -15620
rect 14770 -15680 14800 -15660
rect 14750 -15720 14800 -15680
rect 14860 -15680 14890 -15660
rect 14860 -15720 14910 -15680
rect 14750 -15790 14910 -15720
rect 14750 -15830 14800 -15790
rect 14770 -15850 14800 -15830
rect 14860 -15830 14910 -15790
rect 14860 -15850 14890 -15830
rect 14970 -15890 15030 -15630
rect 14630 -15900 14710 -15890
rect 14630 -15960 14640 -15900
rect 14700 -15910 14710 -15900
rect 14950 -15900 15030 -15890
rect 14950 -15910 14960 -15900
rect 14700 -15960 14960 -15910
rect 15020 -15960 15030 -15900
rect 14630 -15970 15030 -15960
rect 15086 -15550 15486 -15540
rect 15086 -15610 15096 -15550
rect 15156 -15600 15416 -15550
rect 15156 -15610 15166 -15600
rect 15086 -15620 15166 -15610
rect 15406 -15610 15416 -15600
rect 15476 -15610 15486 -15550
rect 15406 -15620 15486 -15610
rect 15086 -15890 15146 -15620
rect 15416 -15630 15486 -15620
rect 15226 -15680 15256 -15660
rect 15206 -15720 15256 -15680
rect 15316 -15680 15346 -15660
rect 15316 -15720 15366 -15680
rect 15206 -15790 15366 -15720
rect 15206 -15830 15256 -15790
rect 15226 -15850 15256 -15830
rect 15316 -15830 15366 -15790
rect 15316 -15850 15346 -15830
rect 15426 -15890 15486 -15630
rect 15086 -15900 15166 -15890
rect 15086 -15960 15096 -15900
rect 15156 -15910 15166 -15900
rect 15406 -15900 15486 -15890
rect 15406 -15910 15416 -15900
rect 15156 -15960 15416 -15910
rect 15476 -15960 15486 -15900
rect 15086 -15970 15486 -15960
rect 0 -16052 400 -16042
rect 0 -16112 10 -16052
rect 70 -16102 330 -16052
rect 70 -16112 80 -16102
rect 0 -16122 80 -16112
rect 320 -16112 330 -16102
rect 390 -16112 400 -16052
rect 320 -16122 400 -16112
rect 0 -16392 60 -16122
rect 330 -16132 400 -16122
rect 140 -16182 170 -16162
rect 120 -16222 170 -16182
rect 230 -16182 260 -16162
rect 230 -16222 280 -16182
rect 120 -16292 280 -16222
rect 120 -16332 170 -16292
rect 140 -16352 170 -16332
rect 230 -16332 280 -16292
rect 230 -16352 260 -16332
rect 340 -16392 400 -16132
rect 0 -16402 80 -16392
rect 0 -16462 10 -16402
rect 70 -16412 80 -16402
rect 320 -16402 400 -16392
rect 320 -16412 330 -16402
rect 70 -16462 330 -16412
rect 390 -16462 400 -16402
rect 0 -16472 400 -16462
rect 456 -16052 856 -16042
rect 456 -16112 466 -16052
rect 526 -16102 786 -16052
rect 526 -16112 536 -16102
rect 456 -16122 536 -16112
rect 776 -16112 786 -16102
rect 846 -16112 856 -16052
rect 776 -16122 856 -16112
rect 456 -16392 516 -16122
rect 786 -16132 856 -16122
rect 596 -16182 626 -16162
rect 576 -16222 626 -16182
rect 686 -16182 716 -16162
rect 686 -16222 736 -16182
rect 576 -16292 736 -16222
rect 576 -16332 626 -16292
rect 596 -16352 626 -16332
rect 686 -16332 736 -16292
rect 686 -16352 716 -16332
rect 796 -16392 856 -16132
rect 456 -16402 536 -16392
rect 456 -16462 466 -16402
rect 526 -16412 536 -16402
rect 776 -16402 856 -16392
rect 776 -16412 786 -16402
rect 526 -16462 786 -16412
rect 846 -16462 856 -16402
rect 456 -16472 856 -16462
rect 912 -16052 1312 -16042
rect 912 -16112 922 -16052
rect 982 -16102 1242 -16052
rect 982 -16112 992 -16102
rect 912 -16122 992 -16112
rect 1232 -16112 1242 -16102
rect 1302 -16112 1312 -16052
rect 1232 -16122 1312 -16112
rect 912 -16392 972 -16122
rect 1242 -16132 1312 -16122
rect 1052 -16182 1082 -16162
rect 1032 -16222 1082 -16182
rect 1142 -16182 1172 -16162
rect 1142 -16222 1192 -16182
rect 1032 -16292 1192 -16222
rect 1032 -16332 1082 -16292
rect 1052 -16352 1082 -16332
rect 1142 -16332 1192 -16292
rect 1142 -16352 1172 -16332
rect 1252 -16392 1312 -16132
rect 912 -16402 992 -16392
rect 912 -16462 922 -16402
rect 982 -16412 992 -16402
rect 1232 -16402 1312 -16392
rect 1232 -16412 1242 -16402
rect 982 -16462 1242 -16412
rect 1302 -16462 1312 -16402
rect 912 -16472 1312 -16462
rect 1370 -16052 1770 -16042
rect 1370 -16112 1380 -16052
rect 1440 -16102 1700 -16052
rect 1440 -16112 1450 -16102
rect 1370 -16122 1450 -16112
rect 1690 -16112 1700 -16102
rect 1760 -16112 1770 -16052
rect 1690 -16122 1770 -16112
rect 1370 -16392 1430 -16122
rect 1700 -16132 1770 -16122
rect 1510 -16182 1540 -16162
rect 1490 -16222 1540 -16182
rect 1600 -16182 1630 -16162
rect 1600 -16222 1650 -16182
rect 1490 -16292 1650 -16222
rect 1490 -16332 1540 -16292
rect 1510 -16352 1540 -16332
rect 1600 -16332 1650 -16292
rect 1600 -16352 1630 -16332
rect 1710 -16392 1770 -16132
rect 1370 -16402 1450 -16392
rect 1370 -16462 1380 -16402
rect 1440 -16412 1450 -16402
rect 1690 -16402 1770 -16392
rect 1690 -16412 1700 -16402
rect 1440 -16462 1700 -16412
rect 1760 -16462 1770 -16402
rect 1370 -16472 1770 -16462
rect 1826 -16052 2226 -16042
rect 1826 -16112 1836 -16052
rect 1896 -16102 2156 -16052
rect 1896 -16112 1906 -16102
rect 1826 -16122 1906 -16112
rect 2146 -16112 2156 -16102
rect 2216 -16112 2226 -16052
rect 2146 -16122 2226 -16112
rect 1826 -16392 1886 -16122
rect 2156 -16132 2226 -16122
rect 1966 -16182 1996 -16162
rect 1946 -16222 1996 -16182
rect 2056 -16182 2086 -16162
rect 2056 -16222 2106 -16182
rect 1946 -16292 2106 -16222
rect 1946 -16332 1996 -16292
rect 1966 -16352 1996 -16332
rect 2056 -16332 2106 -16292
rect 2056 -16352 2086 -16332
rect 2166 -16392 2226 -16132
rect 1826 -16402 1906 -16392
rect 1826 -16462 1836 -16402
rect 1896 -16412 1906 -16402
rect 2146 -16402 2226 -16392
rect 2146 -16412 2156 -16402
rect 1896 -16462 2156 -16412
rect 2216 -16462 2226 -16402
rect 1826 -16472 2226 -16462
rect 2282 -16052 2682 -16042
rect 2282 -16112 2292 -16052
rect 2352 -16102 2612 -16052
rect 2352 -16112 2362 -16102
rect 2282 -16122 2362 -16112
rect 2602 -16112 2612 -16102
rect 2672 -16112 2682 -16052
rect 2602 -16122 2682 -16112
rect 2282 -16392 2342 -16122
rect 2612 -16132 2682 -16122
rect 2422 -16182 2452 -16162
rect 2402 -16222 2452 -16182
rect 2512 -16182 2542 -16162
rect 2512 -16222 2562 -16182
rect 2402 -16292 2562 -16222
rect 2402 -16332 2452 -16292
rect 2422 -16352 2452 -16332
rect 2512 -16332 2562 -16292
rect 2512 -16352 2542 -16332
rect 2622 -16392 2682 -16132
rect 2282 -16402 2362 -16392
rect 2282 -16462 2292 -16402
rect 2352 -16412 2362 -16402
rect 2602 -16402 2682 -16392
rect 2602 -16412 2612 -16402
rect 2352 -16462 2612 -16412
rect 2672 -16462 2682 -16402
rect 2282 -16472 2682 -16462
rect 2740 -16052 3140 -16042
rect 2740 -16112 2750 -16052
rect 2810 -16102 3070 -16052
rect 2810 -16112 2820 -16102
rect 2740 -16122 2820 -16112
rect 3060 -16112 3070 -16102
rect 3130 -16112 3140 -16052
rect 3060 -16122 3140 -16112
rect 2740 -16392 2800 -16122
rect 3070 -16132 3140 -16122
rect 2880 -16182 2910 -16162
rect 2860 -16222 2910 -16182
rect 2970 -16182 3000 -16162
rect 2970 -16222 3020 -16182
rect 2860 -16292 3020 -16222
rect 2860 -16332 2910 -16292
rect 2880 -16352 2910 -16332
rect 2970 -16332 3020 -16292
rect 2970 -16352 3000 -16332
rect 3080 -16392 3140 -16132
rect 2740 -16402 2820 -16392
rect 2740 -16462 2750 -16402
rect 2810 -16412 2820 -16402
rect 3060 -16402 3140 -16392
rect 3060 -16412 3070 -16402
rect 2810 -16462 3070 -16412
rect 3130 -16462 3140 -16402
rect 2740 -16472 3140 -16462
rect 3196 -16052 3596 -16042
rect 3196 -16112 3206 -16052
rect 3266 -16102 3526 -16052
rect 3266 -16112 3276 -16102
rect 3196 -16122 3276 -16112
rect 3516 -16112 3526 -16102
rect 3586 -16112 3596 -16052
rect 3516 -16122 3596 -16112
rect 3196 -16392 3256 -16122
rect 3526 -16132 3596 -16122
rect 3336 -16182 3366 -16162
rect 3316 -16222 3366 -16182
rect 3426 -16182 3456 -16162
rect 3426 -16222 3476 -16182
rect 3316 -16292 3476 -16222
rect 3316 -16332 3366 -16292
rect 3336 -16352 3366 -16332
rect 3426 -16332 3476 -16292
rect 3426 -16352 3456 -16332
rect 3536 -16392 3596 -16132
rect 3196 -16402 3276 -16392
rect 3196 -16462 3206 -16402
rect 3266 -16412 3276 -16402
rect 3516 -16402 3596 -16392
rect 3516 -16412 3526 -16402
rect 3266 -16462 3526 -16412
rect 3586 -16462 3596 -16402
rect 3196 -16472 3596 -16462
rect 3652 -16052 4052 -16042
rect 3652 -16112 3662 -16052
rect 3722 -16102 3982 -16052
rect 3722 -16112 3732 -16102
rect 3652 -16122 3732 -16112
rect 3972 -16112 3982 -16102
rect 4042 -16112 4052 -16052
rect 3972 -16122 4052 -16112
rect 3652 -16392 3712 -16122
rect 3982 -16132 4052 -16122
rect 3792 -16182 3822 -16162
rect 3772 -16222 3822 -16182
rect 3882 -16182 3912 -16162
rect 3882 -16222 3932 -16182
rect 3772 -16292 3932 -16222
rect 3772 -16332 3822 -16292
rect 3792 -16352 3822 -16332
rect 3882 -16332 3932 -16292
rect 3882 -16352 3912 -16332
rect 3992 -16392 4052 -16132
rect 3652 -16402 3732 -16392
rect 3652 -16462 3662 -16402
rect 3722 -16412 3732 -16402
rect 3972 -16402 4052 -16392
rect 3972 -16412 3982 -16402
rect 3722 -16462 3982 -16412
rect 4042 -16462 4052 -16402
rect 3652 -16472 4052 -16462
rect 4110 -16052 4510 -16042
rect 4110 -16112 4120 -16052
rect 4180 -16102 4440 -16052
rect 4180 -16112 4190 -16102
rect 4110 -16122 4190 -16112
rect 4430 -16112 4440 -16102
rect 4500 -16112 4510 -16052
rect 4430 -16122 4510 -16112
rect 4110 -16392 4170 -16122
rect 4440 -16132 4510 -16122
rect 4250 -16182 4280 -16162
rect 4230 -16222 4280 -16182
rect 4340 -16182 4370 -16162
rect 4340 -16222 4390 -16182
rect 4230 -16292 4390 -16222
rect 4230 -16332 4280 -16292
rect 4250 -16352 4280 -16332
rect 4340 -16332 4390 -16292
rect 4340 -16352 4370 -16332
rect 4450 -16392 4510 -16132
rect 4110 -16402 4190 -16392
rect 4110 -16462 4120 -16402
rect 4180 -16412 4190 -16402
rect 4430 -16402 4510 -16392
rect 4430 -16412 4440 -16402
rect 4180 -16462 4440 -16412
rect 4500 -16462 4510 -16402
rect 4110 -16472 4510 -16462
rect 4566 -16052 4966 -16042
rect 4566 -16112 4576 -16052
rect 4636 -16102 4896 -16052
rect 4636 -16112 4646 -16102
rect 4566 -16122 4646 -16112
rect 4886 -16112 4896 -16102
rect 4956 -16112 4966 -16052
rect 4886 -16122 4966 -16112
rect 4566 -16392 4626 -16122
rect 4896 -16132 4966 -16122
rect 4706 -16182 4736 -16162
rect 4686 -16222 4736 -16182
rect 4796 -16182 4826 -16162
rect 4796 -16222 4846 -16182
rect 4686 -16292 4846 -16222
rect 4686 -16332 4736 -16292
rect 4706 -16352 4736 -16332
rect 4796 -16332 4846 -16292
rect 4796 -16352 4826 -16332
rect 4906 -16392 4966 -16132
rect 4566 -16402 4646 -16392
rect 4566 -16462 4576 -16402
rect 4636 -16412 4646 -16402
rect 4886 -16402 4966 -16392
rect 4886 -16412 4896 -16402
rect 4636 -16462 4896 -16412
rect 4956 -16462 4966 -16402
rect 4566 -16472 4966 -16462
rect 5022 -16052 5422 -16042
rect 5022 -16112 5032 -16052
rect 5092 -16102 5352 -16052
rect 5092 -16112 5102 -16102
rect 5022 -16122 5102 -16112
rect 5342 -16112 5352 -16102
rect 5412 -16112 5422 -16052
rect 5342 -16122 5422 -16112
rect 5022 -16392 5082 -16122
rect 5352 -16132 5422 -16122
rect 5162 -16182 5192 -16162
rect 5142 -16222 5192 -16182
rect 5252 -16182 5282 -16162
rect 5252 -16222 5302 -16182
rect 5142 -16292 5302 -16222
rect 5142 -16332 5192 -16292
rect 5162 -16352 5192 -16332
rect 5252 -16332 5302 -16292
rect 5252 -16352 5282 -16332
rect 5362 -16392 5422 -16132
rect 5022 -16402 5102 -16392
rect 5022 -16462 5032 -16402
rect 5092 -16412 5102 -16402
rect 5342 -16402 5422 -16392
rect 5342 -16412 5352 -16402
rect 5092 -16462 5352 -16412
rect 5412 -16462 5422 -16402
rect 5022 -16472 5422 -16462
rect 5480 -16052 5880 -16042
rect 5480 -16112 5490 -16052
rect 5550 -16102 5810 -16052
rect 5550 -16112 5560 -16102
rect 5480 -16122 5560 -16112
rect 5800 -16112 5810 -16102
rect 5870 -16112 5880 -16052
rect 5800 -16122 5880 -16112
rect 5480 -16392 5540 -16122
rect 5810 -16132 5880 -16122
rect 5620 -16182 5650 -16162
rect 5600 -16222 5650 -16182
rect 5710 -16182 5740 -16162
rect 5710 -16222 5760 -16182
rect 5600 -16292 5760 -16222
rect 5600 -16332 5650 -16292
rect 5620 -16352 5650 -16332
rect 5710 -16332 5760 -16292
rect 5710 -16352 5740 -16332
rect 5820 -16392 5880 -16132
rect 5480 -16402 5560 -16392
rect 5480 -16462 5490 -16402
rect 5550 -16412 5560 -16402
rect 5800 -16402 5880 -16392
rect 5800 -16412 5810 -16402
rect 5550 -16462 5810 -16412
rect 5870 -16462 5880 -16402
rect 5480 -16472 5880 -16462
rect 5936 -16052 6336 -16042
rect 5936 -16112 5946 -16052
rect 6006 -16102 6266 -16052
rect 6006 -16112 6016 -16102
rect 5936 -16122 6016 -16112
rect 6256 -16112 6266 -16102
rect 6326 -16112 6336 -16052
rect 6256 -16122 6336 -16112
rect 5936 -16392 5996 -16122
rect 6266 -16132 6336 -16122
rect 6076 -16182 6106 -16162
rect 6056 -16222 6106 -16182
rect 6166 -16182 6196 -16162
rect 6166 -16222 6216 -16182
rect 6056 -16292 6216 -16222
rect 6056 -16332 6106 -16292
rect 6076 -16352 6106 -16332
rect 6166 -16332 6216 -16292
rect 6166 -16352 6196 -16332
rect 6276 -16392 6336 -16132
rect 5936 -16402 6016 -16392
rect 5936 -16462 5946 -16402
rect 6006 -16412 6016 -16402
rect 6256 -16402 6336 -16392
rect 6256 -16412 6266 -16402
rect 6006 -16462 6266 -16412
rect 6326 -16462 6336 -16402
rect 5936 -16472 6336 -16462
rect 6392 -16052 6792 -16042
rect 6392 -16112 6402 -16052
rect 6462 -16102 6722 -16052
rect 6462 -16112 6472 -16102
rect 6392 -16122 6472 -16112
rect 6712 -16112 6722 -16102
rect 6782 -16112 6792 -16052
rect 6712 -16122 6792 -16112
rect 6392 -16392 6452 -16122
rect 6722 -16132 6792 -16122
rect 6532 -16182 6562 -16162
rect 6512 -16222 6562 -16182
rect 6622 -16182 6652 -16162
rect 6622 -16222 6672 -16182
rect 6512 -16292 6672 -16222
rect 6512 -16332 6562 -16292
rect 6532 -16352 6562 -16332
rect 6622 -16332 6672 -16292
rect 6622 -16352 6652 -16332
rect 6732 -16392 6792 -16132
rect 6392 -16402 6472 -16392
rect 6392 -16462 6402 -16402
rect 6462 -16412 6472 -16402
rect 6712 -16402 6792 -16392
rect 6712 -16412 6722 -16402
rect 6462 -16462 6722 -16412
rect 6782 -16462 6792 -16402
rect 6392 -16472 6792 -16462
rect 6850 -16052 7250 -16042
rect 6850 -16112 6860 -16052
rect 6920 -16102 7180 -16052
rect 6920 -16112 6930 -16102
rect 6850 -16122 6930 -16112
rect 7170 -16112 7180 -16102
rect 7240 -16112 7250 -16052
rect 7170 -16122 7250 -16112
rect 6850 -16392 6910 -16122
rect 7180 -16132 7250 -16122
rect 6990 -16182 7020 -16162
rect 6970 -16222 7020 -16182
rect 7080 -16182 7110 -16162
rect 7080 -16222 7130 -16182
rect 6970 -16292 7130 -16222
rect 6970 -16332 7020 -16292
rect 6990 -16352 7020 -16332
rect 7080 -16332 7130 -16292
rect 7080 -16352 7110 -16332
rect 7190 -16392 7250 -16132
rect 6850 -16402 6930 -16392
rect 6850 -16462 6860 -16402
rect 6920 -16412 6930 -16402
rect 7170 -16402 7250 -16392
rect 7170 -16412 7180 -16402
rect 6920 -16462 7180 -16412
rect 7240 -16462 7250 -16402
rect 6850 -16472 7250 -16462
rect 7306 -16052 7706 -16042
rect 7306 -16112 7316 -16052
rect 7376 -16102 7636 -16052
rect 7376 -16112 7386 -16102
rect 7306 -16122 7386 -16112
rect 7626 -16112 7636 -16102
rect 7696 -16112 7706 -16052
rect 7626 -16122 7706 -16112
rect 7306 -16392 7366 -16122
rect 7636 -16132 7706 -16122
rect 7446 -16182 7476 -16162
rect 7426 -16222 7476 -16182
rect 7536 -16182 7566 -16162
rect 7536 -16222 7586 -16182
rect 7426 -16292 7586 -16222
rect 7426 -16332 7476 -16292
rect 7446 -16352 7476 -16332
rect 7536 -16332 7586 -16292
rect 7536 -16352 7566 -16332
rect 7646 -16392 7706 -16132
rect 7306 -16402 7386 -16392
rect 7306 -16462 7316 -16402
rect 7376 -16412 7386 -16402
rect 7626 -16402 7706 -16392
rect 7626 -16412 7636 -16402
rect 7376 -16462 7636 -16412
rect 7696 -16462 7706 -16402
rect 7306 -16472 7706 -16462
rect 7762 -16052 8162 -16042
rect 7762 -16112 7772 -16052
rect 7832 -16102 8092 -16052
rect 7832 -16112 7842 -16102
rect 7762 -16122 7842 -16112
rect 8082 -16112 8092 -16102
rect 8152 -16112 8162 -16052
rect 8082 -16122 8162 -16112
rect 7762 -16392 7822 -16122
rect 8092 -16132 8162 -16122
rect 7902 -16182 7932 -16162
rect 7882 -16222 7932 -16182
rect 7992 -16182 8022 -16162
rect 7992 -16222 8042 -16182
rect 7882 -16292 8042 -16222
rect 7882 -16332 7932 -16292
rect 7902 -16352 7932 -16332
rect 7992 -16332 8042 -16292
rect 7992 -16352 8022 -16332
rect 8102 -16392 8162 -16132
rect 7762 -16402 7842 -16392
rect 7762 -16462 7772 -16402
rect 7832 -16412 7842 -16402
rect 8082 -16402 8162 -16392
rect 8082 -16412 8092 -16402
rect 7832 -16462 8092 -16412
rect 8152 -16462 8162 -16402
rect 7762 -16472 8162 -16462
rect 8236 -16052 8636 -16042
rect 8236 -16112 8246 -16052
rect 8306 -16102 8566 -16052
rect 8306 -16112 8316 -16102
rect 8236 -16122 8316 -16112
rect 8556 -16112 8566 -16102
rect 8626 -16112 8636 -16052
rect 8556 -16122 8636 -16112
rect 8236 -16392 8296 -16122
rect 8566 -16132 8636 -16122
rect 8376 -16182 8406 -16162
rect 8356 -16222 8406 -16182
rect 8466 -16182 8496 -16162
rect 8466 -16222 8516 -16182
rect 8356 -16292 8516 -16222
rect 8356 -16332 8406 -16292
rect 8376 -16352 8406 -16332
rect 8466 -16332 8516 -16292
rect 8466 -16352 8496 -16332
rect 8576 -16392 8636 -16132
rect 8236 -16402 8316 -16392
rect 8236 -16462 8246 -16402
rect 8306 -16412 8316 -16402
rect 8556 -16402 8636 -16392
rect 8556 -16412 8566 -16402
rect 8306 -16462 8566 -16412
rect 8626 -16462 8636 -16402
rect 8236 -16472 8636 -16462
rect 8692 -16052 9092 -16042
rect 8692 -16112 8702 -16052
rect 8762 -16102 9022 -16052
rect 8762 -16112 8772 -16102
rect 8692 -16122 8772 -16112
rect 9012 -16112 9022 -16102
rect 9082 -16112 9092 -16052
rect 9012 -16122 9092 -16112
rect 8692 -16392 8752 -16122
rect 9022 -16132 9092 -16122
rect 8832 -16182 8862 -16162
rect 8812 -16222 8862 -16182
rect 8922 -16182 8952 -16162
rect 8922 -16222 8972 -16182
rect 8812 -16292 8972 -16222
rect 8812 -16332 8862 -16292
rect 8832 -16352 8862 -16332
rect 8922 -16332 8972 -16292
rect 8922 -16352 8952 -16332
rect 9032 -16392 9092 -16132
rect 8692 -16402 8772 -16392
rect 8692 -16462 8702 -16402
rect 8762 -16412 8772 -16402
rect 9012 -16402 9092 -16392
rect 9012 -16412 9022 -16402
rect 8762 -16462 9022 -16412
rect 9082 -16462 9092 -16402
rect 8692 -16472 9092 -16462
rect 9150 -16052 9550 -16042
rect 9150 -16112 9160 -16052
rect 9220 -16102 9480 -16052
rect 9220 -16112 9230 -16102
rect 9150 -16122 9230 -16112
rect 9470 -16112 9480 -16102
rect 9540 -16112 9550 -16052
rect 9470 -16122 9550 -16112
rect 9150 -16392 9210 -16122
rect 9480 -16132 9550 -16122
rect 9290 -16182 9320 -16162
rect 9270 -16222 9320 -16182
rect 9380 -16182 9410 -16162
rect 9380 -16222 9430 -16182
rect 9270 -16292 9430 -16222
rect 9270 -16332 9320 -16292
rect 9290 -16352 9320 -16332
rect 9380 -16332 9430 -16292
rect 9380 -16352 9410 -16332
rect 9490 -16392 9550 -16132
rect 9150 -16402 9230 -16392
rect 9150 -16462 9160 -16402
rect 9220 -16412 9230 -16402
rect 9470 -16402 9550 -16392
rect 9470 -16412 9480 -16402
rect 9220 -16462 9480 -16412
rect 9540 -16462 9550 -16402
rect 9150 -16472 9550 -16462
rect 9606 -16052 10006 -16042
rect 9606 -16112 9616 -16052
rect 9676 -16102 9936 -16052
rect 9676 -16112 9686 -16102
rect 9606 -16122 9686 -16112
rect 9926 -16112 9936 -16102
rect 9996 -16112 10006 -16052
rect 9926 -16122 10006 -16112
rect 9606 -16392 9666 -16122
rect 9936 -16132 10006 -16122
rect 9746 -16182 9776 -16162
rect 9726 -16222 9776 -16182
rect 9836 -16182 9866 -16162
rect 9836 -16222 9886 -16182
rect 9726 -16292 9886 -16222
rect 9726 -16332 9776 -16292
rect 9746 -16352 9776 -16332
rect 9836 -16332 9886 -16292
rect 9836 -16352 9866 -16332
rect 9946 -16392 10006 -16132
rect 9606 -16402 9686 -16392
rect 9606 -16462 9616 -16402
rect 9676 -16412 9686 -16402
rect 9926 -16402 10006 -16392
rect 9926 -16412 9936 -16402
rect 9676 -16462 9936 -16412
rect 9996 -16462 10006 -16402
rect 9606 -16472 10006 -16462
rect 10062 -16052 10462 -16042
rect 10062 -16112 10072 -16052
rect 10132 -16102 10392 -16052
rect 10132 -16112 10142 -16102
rect 10062 -16122 10142 -16112
rect 10382 -16112 10392 -16102
rect 10452 -16112 10462 -16052
rect 10382 -16122 10462 -16112
rect 10062 -16392 10122 -16122
rect 10392 -16132 10462 -16122
rect 10202 -16182 10232 -16162
rect 10182 -16222 10232 -16182
rect 10292 -16182 10322 -16162
rect 10292 -16222 10342 -16182
rect 10182 -16292 10342 -16222
rect 10182 -16332 10232 -16292
rect 10202 -16352 10232 -16332
rect 10292 -16332 10342 -16292
rect 10292 -16352 10322 -16332
rect 10402 -16392 10462 -16132
rect 10062 -16402 10142 -16392
rect 10062 -16462 10072 -16402
rect 10132 -16412 10142 -16402
rect 10382 -16402 10462 -16392
rect 10382 -16412 10392 -16402
rect 10132 -16462 10392 -16412
rect 10452 -16462 10462 -16402
rect 10062 -16472 10462 -16462
rect 10520 -16052 10920 -16042
rect 10520 -16112 10530 -16052
rect 10590 -16102 10850 -16052
rect 10590 -16112 10600 -16102
rect 10520 -16122 10600 -16112
rect 10840 -16112 10850 -16102
rect 10910 -16112 10920 -16052
rect 10840 -16122 10920 -16112
rect 10520 -16392 10580 -16122
rect 10850 -16132 10920 -16122
rect 10660 -16182 10690 -16162
rect 10640 -16222 10690 -16182
rect 10750 -16182 10780 -16162
rect 10750 -16222 10800 -16182
rect 10640 -16292 10800 -16222
rect 10640 -16332 10690 -16292
rect 10660 -16352 10690 -16332
rect 10750 -16332 10800 -16292
rect 10750 -16352 10780 -16332
rect 10860 -16392 10920 -16132
rect 10520 -16402 10600 -16392
rect 10520 -16462 10530 -16402
rect 10590 -16412 10600 -16402
rect 10840 -16402 10920 -16392
rect 10840 -16412 10850 -16402
rect 10590 -16462 10850 -16412
rect 10910 -16462 10920 -16402
rect 10520 -16472 10920 -16462
rect 10976 -16052 11376 -16042
rect 10976 -16112 10986 -16052
rect 11046 -16102 11306 -16052
rect 11046 -16112 11056 -16102
rect 10976 -16122 11056 -16112
rect 11296 -16112 11306 -16102
rect 11366 -16112 11376 -16052
rect 11296 -16122 11376 -16112
rect 10976 -16392 11036 -16122
rect 11306 -16132 11376 -16122
rect 11116 -16182 11146 -16162
rect 11096 -16222 11146 -16182
rect 11206 -16182 11236 -16162
rect 11206 -16222 11256 -16182
rect 11096 -16292 11256 -16222
rect 11096 -16332 11146 -16292
rect 11116 -16352 11146 -16332
rect 11206 -16332 11256 -16292
rect 11206 -16352 11236 -16332
rect 11316 -16392 11376 -16132
rect 10976 -16402 11056 -16392
rect 10976 -16462 10986 -16402
rect 11046 -16412 11056 -16402
rect 11296 -16402 11376 -16392
rect 11296 -16412 11306 -16402
rect 11046 -16462 11306 -16412
rect 11366 -16462 11376 -16402
rect 10976 -16472 11376 -16462
rect 11432 -16052 11832 -16042
rect 11432 -16112 11442 -16052
rect 11502 -16102 11762 -16052
rect 11502 -16112 11512 -16102
rect 11432 -16122 11512 -16112
rect 11752 -16112 11762 -16102
rect 11822 -16112 11832 -16052
rect 11752 -16122 11832 -16112
rect 11432 -16392 11492 -16122
rect 11762 -16132 11832 -16122
rect 11572 -16182 11602 -16162
rect 11552 -16222 11602 -16182
rect 11662 -16182 11692 -16162
rect 11662 -16222 11712 -16182
rect 11552 -16292 11712 -16222
rect 11552 -16332 11602 -16292
rect 11572 -16352 11602 -16332
rect 11662 -16332 11712 -16292
rect 11662 -16352 11692 -16332
rect 11772 -16392 11832 -16132
rect 11432 -16402 11512 -16392
rect 11432 -16462 11442 -16402
rect 11502 -16412 11512 -16402
rect 11752 -16402 11832 -16392
rect 11752 -16412 11762 -16402
rect 11502 -16462 11762 -16412
rect 11822 -16462 11832 -16402
rect 11432 -16472 11832 -16462
rect 11890 -16052 12290 -16042
rect 11890 -16112 11900 -16052
rect 11960 -16102 12220 -16052
rect 11960 -16112 11970 -16102
rect 11890 -16122 11970 -16112
rect 12210 -16112 12220 -16102
rect 12280 -16112 12290 -16052
rect 12210 -16122 12290 -16112
rect 11890 -16392 11950 -16122
rect 12220 -16132 12290 -16122
rect 12030 -16182 12060 -16162
rect 12010 -16222 12060 -16182
rect 12120 -16182 12150 -16162
rect 12120 -16222 12170 -16182
rect 12010 -16292 12170 -16222
rect 12010 -16332 12060 -16292
rect 12030 -16352 12060 -16332
rect 12120 -16332 12170 -16292
rect 12120 -16352 12150 -16332
rect 12230 -16392 12290 -16132
rect 11890 -16402 11970 -16392
rect 11890 -16462 11900 -16402
rect 11960 -16412 11970 -16402
rect 12210 -16402 12290 -16392
rect 12210 -16412 12220 -16402
rect 11960 -16462 12220 -16412
rect 12280 -16462 12290 -16402
rect 11890 -16472 12290 -16462
rect 12346 -16052 12746 -16042
rect 12346 -16112 12356 -16052
rect 12416 -16102 12676 -16052
rect 12416 -16112 12426 -16102
rect 12346 -16122 12426 -16112
rect 12666 -16112 12676 -16102
rect 12736 -16112 12746 -16052
rect 12666 -16122 12746 -16112
rect 12346 -16392 12406 -16122
rect 12676 -16132 12746 -16122
rect 12486 -16182 12516 -16162
rect 12466 -16222 12516 -16182
rect 12576 -16182 12606 -16162
rect 12576 -16222 12626 -16182
rect 12466 -16292 12626 -16222
rect 12466 -16332 12516 -16292
rect 12486 -16352 12516 -16332
rect 12576 -16332 12626 -16292
rect 12576 -16352 12606 -16332
rect 12686 -16392 12746 -16132
rect 12346 -16402 12426 -16392
rect 12346 -16462 12356 -16402
rect 12416 -16412 12426 -16402
rect 12666 -16402 12746 -16392
rect 12666 -16412 12676 -16402
rect 12416 -16462 12676 -16412
rect 12736 -16462 12746 -16402
rect 12346 -16472 12746 -16462
rect 12802 -16052 13202 -16042
rect 12802 -16112 12812 -16052
rect 12872 -16102 13132 -16052
rect 12872 -16112 12882 -16102
rect 12802 -16122 12882 -16112
rect 13122 -16112 13132 -16102
rect 13192 -16112 13202 -16052
rect 13122 -16122 13202 -16112
rect 12802 -16392 12862 -16122
rect 13132 -16132 13202 -16122
rect 12942 -16182 12972 -16162
rect 12922 -16222 12972 -16182
rect 13032 -16182 13062 -16162
rect 13032 -16222 13082 -16182
rect 12922 -16292 13082 -16222
rect 12922 -16332 12972 -16292
rect 12942 -16352 12972 -16332
rect 13032 -16332 13082 -16292
rect 13032 -16352 13062 -16332
rect 13142 -16392 13202 -16132
rect 12802 -16402 12882 -16392
rect 12802 -16462 12812 -16402
rect 12872 -16412 12882 -16402
rect 13122 -16402 13202 -16392
rect 13122 -16412 13132 -16402
rect 12872 -16462 13132 -16412
rect 13192 -16462 13202 -16402
rect 12802 -16472 13202 -16462
rect 13260 -16052 13660 -16042
rect 13260 -16112 13270 -16052
rect 13330 -16102 13590 -16052
rect 13330 -16112 13340 -16102
rect 13260 -16122 13340 -16112
rect 13580 -16112 13590 -16102
rect 13650 -16112 13660 -16052
rect 13580 -16122 13660 -16112
rect 13260 -16392 13320 -16122
rect 13590 -16132 13660 -16122
rect 13400 -16182 13430 -16162
rect 13380 -16222 13430 -16182
rect 13490 -16182 13520 -16162
rect 13490 -16222 13540 -16182
rect 13380 -16292 13540 -16222
rect 13380 -16332 13430 -16292
rect 13400 -16352 13430 -16332
rect 13490 -16332 13540 -16292
rect 13490 -16352 13520 -16332
rect 13600 -16392 13660 -16132
rect 13260 -16402 13340 -16392
rect 13260 -16462 13270 -16402
rect 13330 -16412 13340 -16402
rect 13580 -16402 13660 -16392
rect 13580 -16412 13590 -16402
rect 13330 -16462 13590 -16412
rect 13650 -16462 13660 -16402
rect 13260 -16472 13660 -16462
rect 13716 -16052 14116 -16042
rect 13716 -16112 13726 -16052
rect 13786 -16102 14046 -16052
rect 13786 -16112 13796 -16102
rect 13716 -16122 13796 -16112
rect 14036 -16112 14046 -16102
rect 14106 -16112 14116 -16052
rect 14036 -16122 14116 -16112
rect 13716 -16392 13776 -16122
rect 14046 -16132 14116 -16122
rect 13856 -16182 13886 -16162
rect 13836 -16222 13886 -16182
rect 13946 -16182 13976 -16162
rect 13946 -16222 13996 -16182
rect 13836 -16292 13996 -16222
rect 13836 -16332 13886 -16292
rect 13856 -16352 13886 -16332
rect 13946 -16332 13996 -16292
rect 13946 -16352 13976 -16332
rect 14056 -16392 14116 -16132
rect 13716 -16402 13796 -16392
rect 13716 -16462 13726 -16402
rect 13786 -16412 13796 -16402
rect 14036 -16402 14116 -16392
rect 14036 -16412 14046 -16402
rect 13786 -16462 14046 -16412
rect 14106 -16462 14116 -16402
rect 13716 -16472 14116 -16462
rect 14172 -16052 14572 -16042
rect 14172 -16112 14182 -16052
rect 14242 -16102 14502 -16052
rect 14242 -16112 14252 -16102
rect 14172 -16122 14252 -16112
rect 14492 -16112 14502 -16102
rect 14562 -16112 14572 -16052
rect 14492 -16122 14572 -16112
rect 14172 -16392 14232 -16122
rect 14502 -16132 14572 -16122
rect 14312 -16182 14342 -16162
rect 14292 -16222 14342 -16182
rect 14402 -16182 14432 -16162
rect 14402 -16222 14452 -16182
rect 14292 -16292 14452 -16222
rect 14292 -16332 14342 -16292
rect 14312 -16352 14342 -16332
rect 14402 -16332 14452 -16292
rect 14402 -16352 14432 -16332
rect 14512 -16392 14572 -16132
rect 14172 -16402 14252 -16392
rect 14172 -16462 14182 -16402
rect 14242 -16412 14252 -16402
rect 14492 -16402 14572 -16392
rect 14492 -16412 14502 -16402
rect 14242 -16462 14502 -16412
rect 14562 -16462 14572 -16402
rect 14172 -16472 14572 -16462
rect 14630 -16052 15030 -16042
rect 14630 -16112 14640 -16052
rect 14700 -16102 14960 -16052
rect 14700 -16112 14710 -16102
rect 14630 -16122 14710 -16112
rect 14950 -16112 14960 -16102
rect 15020 -16112 15030 -16052
rect 14950 -16122 15030 -16112
rect 14630 -16392 14690 -16122
rect 14960 -16132 15030 -16122
rect 14770 -16182 14800 -16162
rect 14750 -16222 14800 -16182
rect 14860 -16182 14890 -16162
rect 14860 -16222 14910 -16182
rect 14750 -16292 14910 -16222
rect 14750 -16332 14800 -16292
rect 14770 -16352 14800 -16332
rect 14860 -16332 14910 -16292
rect 14860 -16352 14890 -16332
rect 14970 -16392 15030 -16132
rect 14630 -16402 14710 -16392
rect 14630 -16462 14640 -16402
rect 14700 -16412 14710 -16402
rect 14950 -16402 15030 -16392
rect 14950 -16412 14960 -16402
rect 14700 -16462 14960 -16412
rect 15020 -16462 15030 -16402
rect 14630 -16472 15030 -16462
rect 15086 -16052 15486 -16042
rect 15086 -16112 15096 -16052
rect 15156 -16102 15416 -16052
rect 15156 -16112 15166 -16102
rect 15086 -16122 15166 -16112
rect 15406 -16112 15416 -16102
rect 15476 -16112 15486 -16052
rect 15406 -16122 15486 -16112
rect 15086 -16392 15146 -16122
rect 15416 -16132 15486 -16122
rect 15226 -16182 15256 -16162
rect 15206 -16222 15256 -16182
rect 15316 -16182 15346 -16162
rect 15316 -16222 15366 -16182
rect 15206 -16292 15366 -16222
rect 15206 -16332 15256 -16292
rect 15226 -16352 15256 -16332
rect 15316 -16332 15366 -16292
rect 15316 -16352 15346 -16332
rect 15426 -16392 15486 -16132
rect 15086 -16402 15166 -16392
rect 15086 -16462 15096 -16402
rect 15156 -16412 15166 -16402
rect 15406 -16402 15486 -16392
rect 15406 -16412 15416 -16402
rect 15156 -16462 15416 -16412
rect 15476 -16462 15486 -16402
rect 15086 -16472 15486 -16462
rect 0 -16544 400 -16534
rect 0 -16604 10 -16544
rect 70 -16594 330 -16544
rect 70 -16604 80 -16594
rect 0 -16614 80 -16604
rect 320 -16604 330 -16594
rect 390 -16604 400 -16544
rect 320 -16614 400 -16604
rect 0 -16884 60 -16614
rect 330 -16624 400 -16614
rect 140 -16674 170 -16654
rect 120 -16714 170 -16674
rect 230 -16674 260 -16654
rect 230 -16714 280 -16674
rect 120 -16784 280 -16714
rect 120 -16824 170 -16784
rect 140 -16844 170 -16824
rect 230 -16824 280 -16784
rect 230 -16844 260 -16824
rect 340 -16884 400 -16624
rect 0 -16894 80 -16884
rect 0 -16954 10 -16894
rect 70 -16904 80 -16894
rect 320 -16894 400 -16884
rect 320 -16904 330 -16894
rect 70 -16954 330 -16904
rect 390 -16954 400 -16894
rect 0 -16964 400 -16954
rect 456 -16544 856 -16534
rect 456 -16604 466 -16544
rect 526 -16594 786 -16544
rect 526 -16604 536 -16594
rect 456 -16614 536 -16604
rect 776 -16604 786 -16594
rect 846 -16604 856 -16544
rect 776 -16614 856 -16604
rect 456 -16884 516 -16614
rect 786 -16624 856 -16614
rect 596 -16674 626 -16654
rect 576 -16714 626 -16674
rect 686 -16674 716 -16654
rect 686 -16714 736 -16674
rect 576 -16784 736 -16714
rect 576 -16824 626 -16784
rect 596 -16844 626 -16824
rect 686 -16824 736 -16784
rect 686 -16844 716 -16824
rect 796 -16884 856 -16624
rect 456 -16894 536 -16884
rect 456 -16954 466 -16894
rect 526 -16904 536 -16894
rect 776 -16894 856 -16884
rect 776 -16904 786 -16894
rect 526 -16954 786 -16904
rect 846 -16954 856 -16894
rect 456 -16964 856 -16954
rect 912 -16544 1312 -16534
rect 912 -16604 922 -16544
rect 982 -16594 1242 -16544
rect 982 -16604 992 -16594
rect 912 -16614 992 -16604
rect 1232 -16604 1242 -16594
rect 1302 -16604 1312 -16544
rect 1232 -16614 1312 -16604
rect 912 -16884 972 -16614
rect 1242 -16624 1312 -16614
rect 1052 -16674 1082 -16654
rect 1032 -16714 1082 -16674
rect 1142 -16674 1172 -16654
rect 1142 -16714 1192 -16674
rect 1032 -16784 1192 -16714
rect 1032 -16824 1082 -16784
rect 1052 -16844 1082 -16824
rect 1142 -16824 1192 -16784
rect 1142 -16844 1172 -16824
rect 1252 -16884 1312 -16624
rect 912 -16894 992 -16884
rect 912 -16954 922 -16894
rect 982 -16904 992 -16894
rect 1232 -16894 1312 -16884
rect 1232 -16904 1242 -16894
rect 982 -16954 1242 -16904
rect 1302 -16954 1312 -16894
rect 912 -16964 1312 -16954
rect 1370 -16544 1770 -16534
rect 1370 -16604 1380 -16544
rect 1440 -16594 1700 -16544
rect 1440 -16604 1450 -16594
rect 1370 -16614 1450 -16604
rect 1690 -16604 1700 -16594
rect 1760 -16604 1770 -16544
rect 1690 -16614 1770 -16604
rect 1370 -16884 1430 -16614
rect 1700 -16624 1770 -16614
rect 1510 -16674 1540 -16654
rect 1490 -16714 1540 -16674
rect 1600 -16674 1630 -16654
rect 1600 -16714 1650 -16674
rect 1490 -16784 1650 -16714
rect 1490 -16824 1540 -16784
rect 1510 -16844 1540 -16824
rect 1600 -16824 1650 -16784
rect 1600 -16844 1630 -16824
rect 1710 -16884 1770 -16624
rect 1370 -16894 1450 -16884
rect 1370 -16954 1380 -16894
rect 1440 -16904 1450 -16894
rect 1690 -16894 1770 -16884
rect 1690 -16904 1700 -16894
rect 1440 -16954 1700 -16904
rect 1760 -16954 1770 -16894
rect 1370 -16964 1770 -16954
rect 1826 -16544 2226 -16534
rect 1826 -16604 1836 -16544
rect 1896 -16594 2156 -16544
rect 1896 -16604 1906 -16594
rect 1826 -16614 1906 -16604
rect 2146 -16604 2156 -16594
rect 2216 -16604 2226 -16544
rect 2146 -16614 2226 -16604
rect 1826 -16884 1886 -16614
rect 2156 -16624 2226 -16614
rect 1966 -16674 1996 -16654
rect 1946 -16714 1996 -16674
rect 2056 -16674 2086 -16654
rect 2056 -16714 2106 -16674
rect 1946 -16784 2106 -16714
rect 1946 -16824 1996 -16784
rect 1966 -16844 1996 -16824
rect 2056 -16824 2106 -16784
rect 2056 -16844 2086 -16824
rect 2166 -16884 2226 -16624
rect 1826 -16894 1906 -16884
rect 1826 -16954 1836 -16894
rect 1896 -16904 1906 -16894
rect 2146 -16894 2226 -16884
rect 2146 -16904 2156 -16894
rect 1896 -16954 2156 -16904
rect 2216 -16954 2226 -16894
rect 1826 -16964 2226 -16954
rect 2282 -16544 2682 -16534
rect 2282 -16604 2292 -16544
rect 2352 -16594 2612 -16544
rect 2352 -16604 2362 -16594
rect 2282 -16614 2362 -16604
rect 2602 -16604 2612 -16594
rect 2672 -16604 2682 -16544
rect 2602 -16614 2682 -16604
rect 2282 -16884 2342 -16614
rect 2612 -16624 2682 -16614
rect 2422 -16674 2452 -16654
rect 2402 -16714 2452 -16674
rect 2512 -16674 2542 -16654
rect 2512 -16714 2562 -16674
rect 2402 -16784 2562 -16714
rect 2402 -16824 2452 -16784
rect 2422 -16844 2452 -16824
rect 2512 -16824 2562 -16784
rect 2512 -16844 2542 -16824
rect 2622 -16884 2682 -16624
rect 2282 -16894 2362 -16884
rect 2282 -16954 2292 -16894
rect 2352 -16904 2362 -16894
rect 2602 -16894 2682 -16884
rect 2602 -16904 2612 -16894
rect 2352 -16954 2612 -16904
rect 2672 -16954 2682 -16894
rect 2282 -16964 2682 -16954
rect 2740 -16544 3140 -16534
rect 2740 -16604 2750 -16544
rect 2810 -16594 3070 -16544
rect 2810 -16604 2820 -16594
rect 2740 -16614 2820 -16604
rect 3060 -16604 3070 -16594
rect 3130 -16604 3140 -16544
rect 3060 -16614 3140 -16604
rect 2740 -16884 2800 -16614
rect 3070 -16624 3140 -16614
rect 2880 -16674 2910 -16654
rect 2860 -16714 2910 -16674
rect 2970 -16674 3000 -16654
rect 2970 -16714 3020 -16674
rect 2860 -16784 3020 -16714
rect 2860 -16824 2910 -16784
rect 2880 -16844 2910 -16824
rect 2970 -16824 3020 -16784
rect 2970 -16844 3000 -16824
rect 3080 -16884 3140 -16624
rect 2740 -16894 2820 -16884
rect 2740 -16954 2750 -16894
rect 2810 -16904 2820 -16894
rect 3060 -16894 3140 -16884
rect 3060 -16904 3070 -16894
rect 2810 -16954 3070 -16904
rect 3130 -16954 3140 -16894
rect 2740 -16964 3140 -16954
rect 3196 -16544 3596 -16534
rect 3196 -16604 3206 -16544
rect 3266 -16594 3526 -16544
rect 3266 -16604 3276 -16594
rect 3196 -16614 3276 -16604
rect 3516 -16604 3526 -16594
rect 3586 -16604 3596 -16544
rect 3516 -16614 3596 -16604
rect 3196 -16884 3256 -16614
rect 3526 -16624 3596 -16614
rect 3336 -16674 3366 -16654
rect 3316 -16714 3366 -16674
rect 3426 -16674 3456 -16654
rect 3426 -16714 3476 -16674
rect 3316 -16784 3476 -16714
rect 3316 -16824 3366 -16784
rect 3336 -16844 3366 -16824
rect 3426 -16824 3476 -16784
rect 3426 -16844 3456 -16824
rect 3536 -16884 3596 -16624
rect 3196 -16894 3276 -16884
rect 3196 -16954 3206 -16894
rect 3266 -16904 3276 -16894
rect 3516 -16894 3596 -16884
rect 3516 -16904 3526 -16894
rect 3266 -16954 3526 -16904
rect 3586 -16954 3596 -16894
rect 3196 -16964 3596 -16954
rect 3652 -16544 4052 -16534
rect 3652 -16604 3662 -16544
rect 3722 -16594 3982 -16544
rect 3722 -16604 3732 -16594
rect 3652 -16614 3732 -16604
rect 3972 -16604 3982 -16594
rect 4042 -16604 4052 -16544
rect 3972 -16614 4052 -16604
rect 3652 -16884 3712 -16614
rect 3982 -16624 4052 -16614
rect 3792 -16674 3822 -16654
rect 3772 -16714 3822 -16674
rect 3882 -16674 3912 -16654
rect 3882 -16714 3932 -16674
rect 3772 -16784 3932 -16714
rect 3772 -16824 3822 -16784
rect 3792 -16844 3822 -16824
rect 3882 -16824 3932 -16784
rect 3882 -16844 3912 -16824
rect 3992 -16884 4052 -16624
rect 3652 -16894 3732 -16884
rect 3652 -16954 3662 -16894
rect 3722 -16904 3732 -16894
rect 3972 -16894 4052 -16884
rect 3972 -16904 3982 -16894
rect 3722 -16954 3982 -16904
rect 4042 -16954 4052 -16894
rect 3652 -16964 4052 -16954
rect 4110 -16544 4510 -16534
rect 4110 -16604 4120 -16544
rect 4180 -16594 4440 -16544
rect 4180 -16604 4190 -16594
rect 4110 -16614 4190 -16604
rect 4430 -16604 4440 -16594
rect 4500 -16604 4510 -16544
rect 4430 -16614 4510 -16604
rect 4110 -16884 4170 -16614
rect 4440 -16624 4510 -16614
rect 4250 -16674 4280 -16654
rect 4230 -16714 4280 -16674
rect 4340 -16674 4370 -16654
rect 4340 -16714 4390 -16674
rect 4230 -16784 4390 -16714
rect 4230 -16824 4280 -16784
rect 4250 -16844 4280 -16824
rect 4340 -16824 4390 -16784
rect 4340 -16844 4370 -16824
rect 4450 -16884 4510 -16624
rect 4110 -16894 4190 -16884
rect 4110 -16954 4120 -16894
rect 4180 -16904 4190 -16894
rect 4430 -16894 4510 -16884
rect 4430 -16904 4440 -16894
rect 4180 -16954 4440 -16904
rect 4500 -16954 4510 -16894
rect 4110 -16964 4510 -16954
rect 4566 -16544 4966 -16534
rect 4566 -16604 4576 -16544
rect 4636 -16594 4896 -16544
rect 4636 -16604 4646 -16594
rect 4566 -16614 4646 -16604
rect 4886 -16604 4896 -16594
rect 4956 -16604 4966 -16544
rect 4886 -16614 4966 -16604
rect 4566 -16884 4626 -16614
rect 4896 -16624 4966 -16614
rect 4706 -16674 4736 -16654
rect 4686 -16714 4736 -16674
rect 4796 -16674 4826 -16654
rect 4796 -16714 4846 -16674
rect 4686 -16784 4846 -16714
rect 4686 -16824 4736 -16784
rect 4706 -16844 4736 -16824
rect 4796 -16824 4846 -16784
rect 4796 -16844 4826 -16824
rect 4906 -16884 4966 -16624
rect 4566 -16894 4646 -16884
rect 4566 -16954 4576 -16894
rect 4636 -16904 4646 -16894
rect 4886 -16894 4966 -16884
rect 4886 -16904 4896 -16894
rect 4636 -16954 4896 -16904
rect 4956 -16954 4966 -16894
rect 4566 -16964 4966 -16954
rect 5022 -16544 5422 -16534
rect 5022 -16604 5032 -16544
rect 5092 -16594 5352 -16544
rect 5092 -16604 5102 -16594
rect 5022 -16614 5102 -16604
rect 5342 -16604 5352 -16594
rect 5412 -16604 5422 -16544
rect 5342 -16614 5422 -16604
rect 5022 -16884 5082 -16614
rect 5352 -16624 5422 -16614
rect 5162 -16674 5192 -16654
rect 5142 -16714 5192 -16674
rect 5252 -16674 5282 -16654
rect 5252 -16714 5302 -16674
rect 5142 -16784 5302 -16714
rect 5142 -16824 5192 -16784
rect 5162 -16844 5192 -16824
rect 5252 -16824 5302 -16784
rect 5252 -16844 5282 -16824
rect 5362 -16884 5422 -16624
rect 5022 -16894 5102 -16884
rect 5022 -16954 5032 -16894
rect 5092 -16904 5102 -16894
rect 5342 -16894 5422 -16884
rect 5342 -16904 5352 -16894
rect 5092 -16954 5352 -16904
rect 5412 -16954 5422 -16894
rect 5022 -16964 5422 -16954
rect 5480 -16544 5880 -16534
rect 5480 -16604 5490 -16544
rect 5550 -16594 5810 -16544
rect 5550 -16604 5560 -16594
rect 5480 -16614 5560 -16604
rect 5800 -16604 5810 -16594
rect 5870 -16604 5880 -16544
rect 5800 -16614 5880 -16604
rect 5480 -16884 5540 -16614
rect 5810 -16624 5880 -16614
rect 5620 -16674 5650 -16654
rect 5600 -16714 5650 -16674
rect 5710 -16674 5740 -16654
rect 5710 -16714 5760 -16674
rect 5600 -16784 5760 -16714
rect 5600 -16824 5650 -16784
rect 5620 -16844 5650 -16824
rect 5710 -16824 5760 -16784
rect 5710 -16844 5740 -16824
rect 5820 -16884 5880 -16624
rect 5480 -16894 5560 -16884
rect 5480 -16954 5490 -16894
rect 5550 -16904 5560 -16894
rect 5800 -16894 5880 -16884
rect 5800 -16904 5810 -16894
rect 5550 -16954 5810 -16904
rect 5870 -16954 5880 -16894
rect 5480 -16964 5880 -16954
rect 5936 -16544 6336 -16534
rect 5936 -16604 5946 -16544
rect 6006 -16594 6266 -16544
rect 6006 -16604 6016 -16594
rect 5936 -16614 6016 -16604
rect 6256 -16604 6266 -16594
rect 6326 -16604 6336 -16544
rect 6256 -16614 6336 -16604
rect 5936 -16884 5996 -16614
rect 6266 -16624 6336 -16614
rect 6076 -16674 6106 -16654
rect 6056 -16714 6106 -16674
rect 6166 -16674 6196 -16654
rect 6166 -16714 6216 -16674
rect 6056 -16784 6216 -16714
rect 6056 -16824 6106 -16784
rect 6076 -16844 6106 -16824
rect 6166 -16824 6216 -16784
rect 6166 -16844 6196 -16824
rect 6276 -16884 6336 -16624
rect 5936 -16894 6016 -16884
rect 5936 -16954 5946 -16894
rect 6006 -16904 6016 -16894
rect 6256 -16894 6336 -16884
rect 6256 -16904 6266 -16894
rect 6006 -16954 6266 -16904
rect 6326 -16954 6336 -16894
rect 5936 -16964 6336 -16954
rect 6392 -16544 6792 -16534
rect 6392 -16604 6402 -16544
rect 6462 -16594 6722 -16544
rect 6462 -16604 6472 -16594
rect 6392 -16614 6472 -16604
rect 6712 -16604 6722 -16594
rect 6782 -16604 6792 -16544
rect 6712 -16614 6792 -16604
rect 6392 -16884 6452 -16614
rect 6722 -16624 6792 -16614
rect 6532 -16674 6562 -16654
rect 6512 -16714 6562 -16674
rect 6622 -16674 6652 -16654
rect 6622 -16714 6672 -16674
rect 6512 -16784 6672 -16714
rect 6512 -16824 6562 -16784
rect 6532 -16844 6562 -16824
rect 6622 -16824 6672 -16784
rect 6622 -16844 6652 -16824
rect 6732 -16884 6792 -16624
rect 6392 -16894 6472 -16884
rect 6392 -16954 6402 -16894
rect 6462 -16904 6472 -16894
rect 6712 -16894 6792 -16884
rect 6712 -16904 6722 -16894
rect 6462 -16954 6722 -16904
rect 6782 -16954 6792 -16894
rect 6392 -16964 6792 -16954
rect 6850 -16544 7250 -16534
rect 6850 -16604 6860 -16544
rect 6920 -16594 7180 -16544
rect 6920 -16604 6930 -16594
rect 6850 -16614 6930 -16604
rect 7170 -16604 7180 -16594
rect 7240 -16604 7250 -16544
rect 7170 -16614 7250 -16604
rect 6850 -16884 6910 -16614
rect 7180 -16624 7250 -16614
rect 6990 -16674 7020 -16654
rect 6970 -16714 7020 -16674
rect 7080 -16674 7110 -16654
rect 7080 -16714 7130 -16674
rect 6970 -16784 7130 -16714
rect 6970 -16824 7020 -16784
rect 6990 -16844 7020 -16824
rect 7080 -16824 7130 -16784
rect 7080 -16844 7110 -16824
rect 7190 -16884 7250 -16624
rect 6850 -16894 6930 -16884
rect 6850 -16954 6860 -16894
rect 6920 -16904 6930 -16894
rect 7170 -16894 7250 -16884
rect 7170 -16904 7180 -16894
rect 6920 -16954 7180 -16904
rect 7240 -16954 7250 -16894
rect 6850 -16964 7250 -16954
rect 7306 -16544 7706 -16534
rect 7306 -16604 7316 -16544
rect 7376 -16594 7636 -16544
rect 7376 -16604 7386 -16594
rect 7306 -16614 7386 -16604
rect 7626 -16604 7636 -16594
rect 7696 -16604 7706 -16544
rect 7626 -16614 7706 -16604
rect 7306 -16884 7366 -16614
rect 7636 -16624 7706 -16614
rect 7446 -16674 7476 -16654
rect 7426 -16714 7476 -16674
rect 7536 -16674 7566 -16654
rect 7536 -16714 7586 -16674
rect 7426 -16784 7586 -16714
rect 7426 -16824 7476 -16784
rect 7446 -16844 7476 -16824
rect 7536 -16824 7586 -16784
rect 7536 -16844 7566 -16824
rect 7646 -16884 7706 -16624
rect 7306 -16894 7386 -16884
rect 7306 -16954 7316 -16894
rect 7376 -16904 7386 -16894
rect 7626 -16894 7706 -16884
rect 7626 -16904 7636 -16894
rect 7376 -16954 7636 -16904
rect 7696 -16954 7706 -16894
rect 7306 -16964 7706 -16954
rect 7762 -16544 8162 -16534
rect 7762 -16604 7772 -16544
rect 7832 -16594 8092 -16544
rect 7832 -16604 7842 -16594
rect 7762 -16614 7842 -16604
rect 8082 -16604 8092 -16594
rect 8152 -16604 8162 -16544
rect 8082 -16614 8162 -16604
rect 7762 -16884 7822 -16614
rect 8092 -16624 8162 -16614
rect 7902 -16674 7932 -16654
rect 7882 -16714 7932 -16674
rect 7992 -16674 8022 -16654
rect 7992 -16714 8042 -16674
rect 7882 -16784 8042 -16714
rect 7882 -16824 7932 -16784
rect 7902 -16844 7932 -16824
rect 7992 -16824 8042 -16784
rect 7992 -16844 8022 -16824
rect 8102 -16884 8162 -16624
rect 7762 -16894 7842 -16884
rect 7762 -16954 7772 -16894
rect 7832 -16904 7842 -16894
rect 8082 -16894 8162 -16884
rect 8082 -16904 8092 -16894
rect 7832 -16954 8092 -16904
rect 8152 -16954 8162 -16894
rect 7762 -16964 8162 -16954
rect 8236 -16544 8636 -16534
rect 8236 -16604 8246 -16544
rect 8306 -16594 8566 -16544
rect 8306 -16604 8316 -16594
rect 8236 -16614 8316 -16604
rect 8556 -16604 8566 -16594
rect 8626 -16604 8636 -16544
rect 8556 -16614 8636 -16604
rect 8236 -16884 8296 -16614
rect 8566 -16624 8636 -16614
rect 8376 -16674 8406 -16654
rect 8356 -16714 8406 -16674
rect 8466 -16674 8496 -16654
rect 8466 -16714 8516 -16674
rect 8356 -16784 8516 -16714
rect 8356 -16824 8406 -16784
rect 8376 -16844 8406 -16824
rect 8466 -16824 8516 -16784
rect 8466 -16844 8496 -16824
rect 8576 -16884 8636 -16624
rect 8236 -16894 8316 -16884
rect 8236 -16954 8246 -16894
rect 8306 -16904 8316 -16894
rect 8556 -16894 8636 -16884
rect 8556 -16904 8566 -16894
rect 8306 -16954 8566 -16904
rect 8626 -16954 8636 -16894
rect 8236 -16964 8636 -16954
rect 8692 -16544 9092 -16534
rect 8692 -16604 8702 -16544
rect 8762 -16594 9022 -16544
rect 8762 -16604 8772 -16594
rect 8692 -16614 8772 -16604
rect 9012 -16604 9022 -16594
rect 9082 -16604 9092 -16544
rect 9012 -16614 9092 -16604
rect 8692 -16884 8752 -16614
rect 9022 -16624 9092 -16614
rect 8832 -16674 8862 -16654
rect 8812 -16714 8862 -16674
rect 8922 -16674 8952 -16654
rect 8922 -16714 8972 -16674
rect 8812 -16784 8972 -16714
rect 8812 -16824 8862 -16784
rect 8832 -16844 8862 -16824
rect 8922 -16824 8972 -16784
rect 8922 -16844 8952 -16824
rect 9032 -16884 9092 -16624
rect 8692 -16894 8772 -16884
rect 8692 -16954 8702 -16894
rect 8762 -16904 8772 -16894
rect 9012 -16894 9092 -16884
rect 9012 -16904 9022 -16894
rect 8762 -16954 9022 -16904
rect 9082 -16954 9092 -16894
rect 8692 -16964 9092 -16954
rect 9150 -16544 9550 -16534
rect 9150 -16604 9160 -16544
rect 9220 -16594 9480 -16544
rect 9220 -16604 9230 -16594
rect 9150 -16614 9230 -16604
rect 9470 -16604 9480 -16594
rect 9540 -16604 9550 -16544
rect 9470 -16614 9550 -16604
rect 9150 -16884 9210 -16614
rect 9480 -16624 9550 -16614
rect 9290 -16674 9320 -16654
rect 9270 -16714 9320 -16674
rect 9380 -16674 9410 -16654
rect 9380 -16714 9430 -16674
rect 9270 -16784 9430 -16714
rect 9270 -16824 9320 -16784
rect 9290 -16844 9320 -16824
rect 9380 -16824 9430 -16784
rect 9380 -16844 9410 -16824
rect 9490 -16884 9550 -16624
rect 9150 -16894 9230 -16884
rect 9150 -16954 9160 -16894
rect 9220 -16904 9230 -16894
rect 9470 -16894 9550 -16884
rect 9470 -16904 9480 -16894
rect 9220 -16954 9480 -16904
rect 9540 -16954 9550 -16894
rect 9150 -16964 9550 -16954
rect 9606 -16544 10006 -16534
rect 9606 -16604 9616 -16544
rect 9676 -16594 9936 -16544
rect 9676 -16604 9686 -16594
rect 9606 -16614 9686 -16604
rect 9926 -16604 9936 -16594
rect 9996 -16604 10006 -16544
rect 9926 -16614 10006 -16604
rect 9606 -16884 9666 -16614
rect 9936 -16624 10006 -16614
rect 9746 -16674 9776 -16654
rect 9726 -16714 9776 -16674
rect 9836 -16674 9866 -16654
rect 9836 -16714 9886 -16674
rect 9726 -16784 9886 -16714
rect 9726 -16824 9776 -16784
rect 9746 -16844 9776 -16824
rect 9836 -16824 9886 -16784
rect 9836 -16844 9866 -16824
rect 9946 -16884 10006 -16624
rect 9606 -16894 9686 -16884
rect 9606 -16954 9616 -16894
rect 9676 -16904 9686 -16894
rect 9926 -16894 10006 -16884
rect 9926 -16904 9936 -16894
rect 9676 -16954 9936 -16904
rect 9996 -16954 10006 -16894
rect 9606 -16964 10006 -16954
rect 10062 -16544 10462 -16534
rect 10062 -16604 10072 -16544
rect 10132 -16594 10392 -16544
rect 10132 -16604 10142 -16594
rect 10062 -16614 10142 -16604
rect 10382 -16604 10392 -16594
rect 10452 -16604 10462 -16544
rect 10382 -16614 10462 -16604
rect 10062 -16884 10122 -16614
rect 10392 -16624 10462 -16614
rect 10202 -16674 10232 -16654
rect 10182 -16714 10232 -16674
rect 10292 -16674 10322 -16654
rect 10292 -16714 10342 -16674
rect 10182 -16784 10342 -16714
rect 10182 -16824 10232 -16784
rect 10202 -16844 10232 -16824
rect 10292 -16824 10342 -16784
rect 10292 -16844 10322 -16824
rect 10402 -16884 10462 -16624
rect 10062 -16894 10142 -16884
rect 10062 -16954 10072 -16894
rect 10132 -16904 10142 -16894
rect 10382 -16894 10462 -16884
rect 10382 -16904 10392 -16894
rect 10132 -16954 10392 -16904
rect 10452 -16954 10462 -16894
rect 10062 -16964 10462 -16954
rect 10520 -16544 10920 -16534
rect 10520 -16604 10530 -16544
rect 10590 -16594 10850 -16544
rect 10590 -16604 10600 -16594
rect 10520 -16614 10600 -16604
rect 10840 -16604 10850 -16594
rect 10910 -16604 10920 -16544
rect 10840 -16614 10920 -16604
rect 10520 -16884 10580 -16614
rect 10850 -16624 10920 -16614
rect 10660 -16674 10690 -16654
rect 10640 -16714 10690 -16674
rect 10750 -16674 10780 -16654
rect 10750 -16714 10800 -16674
rect 10640 -16784 10800 -16714
rect 10640 -16824 10690 -16784
rect 10660 -16844 10690 -16824
rect 10750 -16824 10800 -16784
rect 10750 -16844 10780 -16824
rect 10860 -16884 10920 -16624
rect 10520 -16894 10600 -16884
rect 10520 -16954 10530 -16894
rect 10590 -16904 10600 -16894
rect 10840 -16894 10920 -16884
rect 10840 -16904 10850 -16894
rect 10590 -16954 10850 -16904
rect 10910 -16954 10920 -16894
rect 10520 -16964 10920 -16954
rect 10976 -16544 11376 -16534
rect 10976 -16604 10986 -16544
rect 11046 -16594 11306 -16544
rect 11046 -16604 11056 -16594
rect 10976 -16614 11056 -16604
rect 11296 -16604 11306 -16594
rect 11366 -16604 11376 -16544
rect 11296 -16614 11376 -16604
rect 10976 -16884 11036 -16614
rect 11306 -16624 11376 -16614
rect 11116 -16674 11146 -16654
rect 11096 -16714 11146 -16674
rect 11206 -16674 11236 -16654
rect 11206 -16714 11256 -16674
rect 11096 -16784 11256 -16714
rect 11096 -16824 11146 -16784
rect 11116 -16844 11146 -16824
rect 11206 -16824 11256 -16784
rect 11206 -16844 11236 -16824
rect 11316 -16884 11376 -16624
rect 10976 -16894 11056 -16884
rect 10976 -16954 10986 -16894
rect 11046 -16904 11056 -16894
rect 11296 -16894 11376 -16884
rect 11296 -16904 11306 -16894
rect 11046 -16954 11306 -16904
rect 11366 -16954 11376 -16894
rect 10976 -16964 11376 -16954
rect 11432 -16544 11832 -16534
rect 11432 -16604 11442 -16544
rect 11502 -16594 11762 -16544
rect 11502 -16604 11512 -16594
rect 11432 -16614 11512 -16604
rect 11752 -16604 11762 -16594
rect 11822 -16604 11832 -16544
rect 11752 -16614 11832 -16604
rect 11432 -16884 11492 -16614
rect 11762 -16624 11832 -16614
rect 11572 -16674 11602 -16654
rect 11552 -16714 11602 -16674
rect 11662 -16674 11692 -16654
rect 11662 -16714 11712 -16674
rect 11552 -16784 11712 -16714
rect 11552 -16824 11602 -16784
rect 11572 -16844 11602 -16824
rect 11662 -16824 11712 -16784
rect 11662 -16844 11692 -16824
rect 11772 -16884 11832 -16624
rect 11432 -16894 11512 -16884
rect 11432 -16954 11442 -16894
rect 11502 -16904 11512 -16894
rect 11752 -16894 11832 -16884
rect 11752 -16904 11762 -16894
rect 11502 -16954 11762 -16904
rect 11822 -16954 11832 -16894
rect 11432 -16964 11832 -16954
rect 11890 -16544 12290 -16534
rect 11890 -16604 11900 -16544
rect 11960 -16594 12220 -16544
rect 11960 -16604 11970 -16594
rect 11890 -16614 11970 -16604
rect 12210 -16604 12220 -16594
rect 12280 -16604 12290 -16544
rect 12210 -16614 12290 -16604
rect 11890 -16884 11950 -16614
rect 12220 -16624 12290 -16614
rect 12030 -16674 12060 -16654
rect 12010 -16714 12060 -16674
rect 12120 -16674 12150 -16654
rect 12120 -16714 12170 -16674
rect 12010 -16784 12170 -16714
rect 12010 -16824 12060 -16784
rect 12030 -16844 12060 -16824
rect 12120 -16824 12170 -16784
rect 12120 -16844 12150 -16824
rect 12230 -16884 12290 -16624
rect 11890 -16894 11970 -16884
rect 11890 -16954 11900 -16894
rect 11960 -16904 11970 -16894
rect 12210 -16894 12290 -16884
rect 12210 -16904 12220 -16894
rect 11960 -16954 12220 -16904
rect 12280 -16954 12290 -16894
rect 11890 -16964 12290 -16954
rect 12346 -16544 12746 -16534
rect 12346 -16604 12356 -16544
rect 12416 -16594 12676 -16544
rect 12416 -16604 12426 -16594
rect 12346 -16614 12426 -16604
rect 12666 -16604 12676 -16594
rect 12736 -16604 12746 -16544
rect 12666 -16614 12746 -16604
rect 12346 -16884 12406 -16614
rect 12676 -16624 12746 -16614
rect 12486 -16674 12516 -16654
rect 12466 -16714 12516 -16674
rect 12576 -16674 12606 -16654
rect 12576 -16714 12626 -16674
rect 12466 -16784 12626 -16714
rect 12466 -16824 12516 -16784
rect 12486 -16844 12516 -16824
rect 12576 -16824 12626 -16784
rect 12576 -16844 12606 -16824
rect 12686 -16884 12746 -16624
rect 12346 -16894 12426 -16884
rect 12346 -16954 12356 -16894
rect 12416 -16904 12426 -16894
rect 12666 -16894 12746 -16884
rect 12666 -16904 12676 -16894
rect 12416 -16954 12676 -16904
rect 12736 -16954 12746 -16894
rect 12346 -16964 12746 -16954
rect 12802 -16544 13202 -16534
rect 12802 -16604 12812 -16544
rect 12872 -16594 13132 -16544
rect 12872 -16604 12882 -16594
rect 12802 -16614 12882 -16604
rect 13122 -16604 13132 -16594
rect 13192 -16604 13202 -16544
rect 13122 -16614 13202 -16604
rect 12802 -16884 12862 -16614
rect 13132 -16624 13202 -16614
rect 12942 -16674 12972 -16654
rect 12922 -16714 12972 -16674
rect 13032 -16674 13062 -16654
rect 13032 -16714 13082 -16674
rect 12922 -16784 13082 -16714
rect 12922 -16824 12972 -16784
rect 12942 -16844 12972 -16824
rect 13032 -16824 13082 -16784
rect 13032 -16844 13062 -16824
rect 13142 -16884 13202 -16624
rect 12802 -16894 12882 -16884
rect 12802 -16954 12812 -16894
rect 12872 -16904 12882 -16894
rect 13122 -16894 13202 -16884
rect 13122 -16904 13132 -16894
rect 12872 -16954 13132 -16904
rect 13192 -16954 13202 -16894
rect 12802 -16964 13202 -16954
rect 13260 -16544 13660 -16534
rect 13260 -16604 13270 -16544
rect 13330 -16594 13590 -16544
rect 13330 -16604 13340 -16594
rect 13260 -16614 13340 -16604
rect 13580 -16604 13590 -16594
rect 13650 -16604 13660 -16544
rect 13580 -16614 13660 -16604
rect 13260 -16884 13320 -16614
rect 13590 -16624 13660 -16614
rect 13400 -16674 13430 -16654
rect 13380 -16714 13430 -16674
rect 13490 -16674 13520 -16654
rect 13490 -16714 13540 -16674
rect 13380 -16784 13540 -16714
rect 13380 -16824 13430 -16784
rect 13400 -16844 13430 -16824
rect 13490 -16824 13540 -16784
rect 13490 -16844 13520 -16824
rect 13600 -16884 13660 -16624
rect 13260 -16894 13340 -16884
rect 13260 -16954 13270 -16894
rect 13330 -16904 13340 -16894
rect 13580 -16894 13660 -16884
rect 13580 -16904 13590 -16894
rect 13330 -16954 13590 -16904
rect 13650 -16954 13660 -16894
rect 13260 -16964 13660 -16954
rect 13716 -16544 14116 -16534
rect 13716 -16604 13726 -16544
rect 13786 -16594 14046 -16544
rect 13786 -16604 13796 -16594
rect 13716 -16614 13796 -16604
rect 14036 -16604 14046 -16594
rect 14106 -16604 14116 -16544
rect 14036 -16614 14116 -16604
rect 13716 -16884 13776 -16614
rect 14046 -16624 14116 -16614
rect 13856 -16674 13886 -16654
rect 13836 -16714 13886 -16674
rect 13946 -16674 13976 -16654
rect 13946 -16714 13996 -16674
rect 13836 -16784 13996 -16714
rect 13836 -16824 13886 -16784
rect 13856 -16844 13886 -16824
rect 13946 -16824 13996 -16784
rect 13946 -16844 13976 -16824
rect 14056 -16884 14116 -16624
rect 13716 -16894 13796 -16884
rect 13716 -16954 13726 -16894
rect 13786 -16904 13796 -16894
rect 14036 -16894 14116 -16884
rect 14036 -16904 14046 -16894
rect 13786 -16954 14046 -16904
rect 14106 -16954 14116 -16894
rect 13716 -16964 14116 -16954
rect 14172 -16544 14572 -16534
rect 14172 -16604 14182 -16544
rect 14242 -16594 14502 -16544
rect 14242 -16604 14252 -16594
rect 14172 -16614 14252 -16604
rect 14492 -16604 14502 -16594
rect 14562 -16604 14572 -16544
rect 14492 -16614 14572 -16604
rect 14172 -16884 14232 -16614
rect 14502 -16624 14572 -16614
rect 14312 -16674 14342 -16654
rect 14292 -16714 14342 -16674
rect 14402 -16674 14432 -16654
rect 14402 -16714 14452 -16674
rect 14292 -16784 14452 -16714
rect 14292 -16824 14342 -16784
rect 14312 -16844 14342 -16824
rect 14402 -16824 14452 -16784
rect 14402 -16844 14432 -16824
rect 14512 -16884 14572 -16624
rect 14172 -16894 14252 -16884
rect 14172 -16954 14182 -16894
rect 14242 -16904 14252 -16894
rect 14492 -16894 14572 -16884
rect 14492 -16904 14502 -16894
rect 14242 -16954 14502 -16904
rect 14562 -16954 14572 -16894
rect 14172 -16964 14572 -16954
rect 14630 -16544 15030 -16534
rect 14630 -16604 14640 -16544
rect 14700 -16594 14960 -16544
rect 14700 -16604 14710 -16594
rect 14630 -16614 14710 -16604
rect 14950 -16604 14960 -16594
rect 15020 -16604 15030 -16544
rect 14950 -16614 15030 -16604
rect 14630 -16884 14690 -16614
rect 14960 -16624 15030 -16614
rect 14770 -16674 14800 -16654
rect 14750 -16714 14800 -16674
rect 14860 -16674 14890 -16654
rect 14860 -16714 14910 -16674
rect 14750 -16784 14910 -16714
rect 14750 -16824 14800 -16784
rect 14770 -16844 14800 -16824
rect 14860 -16824 14910 -16784
rect 14860 -16844 14890 -16824
rect 14970 -16884 15030 -16624
rect 14630 -16894 14710 -16884
rect 14630 -16954 14640 -16894
rect 14700 -16904 14710 -16894
rect 14950 -16894 15030 -16884
rect 14950 -16904 14960 -16894
rect 14700 -16954 14960 -16904
rect 15020 -16954 15030 -16894
rect 14630 -16964 15030 -16954
rect 15086 -16544 15486 -16534
rect 15086 -16604 15096 -16544
rect 15156 -16594 15416 -16544
rect 15156 -16604 15166 -16594
rect 15086 -16614 15166 -16604
rect 15406 -16604 15416 -16594
rect 15476 -16604 15486 -16544
rect 15406 -16614 15486 -16604
rect 15086 -16884 15146 -16614
rect 15416 -16624 15486 -16614
rect 15226 -16674 15256 -16654
rect 15206 -16714 15256 -16674
rect 15316 -16674 15346 -16654
rect 15316 -16714 15366 -16674
rect 15206 -16784 15366 -16714
rect 15206 -16824 15256 -16784
rect 15226 -16844 15256 -16824
rect 15316 -16824 15366 -16784
rect 15316 -16844 15346 -16824
rect 15426 -16884 15486 -16624
rect 15086 -16894 15166 -16884
rect 15086 -16954 15096 -16894
rect 15156 -16904 15166 -16894
rect 15406 -16894 15486 -16884
rect 15406 -16904 15416 -16894
rect 15156 -16954 15416 -16904
rect 15476 -16954 15486 -16894
rect 15086 -16964 15486 -16954
rect 1 -17041 401 -17031
rect 1 -17101 11 -17041
rect 71 -17091 331 -17041
rect 71 -17101 81 -17091
rect 1 -17111 81 -17101
rect 321 -17101 331 -17091
rect 391 -17101 401 -17041
rect 321 -17111 401 -17101
rect 1 -17381 61 -17111
rect 331 -17121 401 -17111
rect 141 -17171 171 -17151
rect 121 -17211 171 -17171
rect 231 -17171 261 -17151
rect 231 -17211 281 -17171
rect 121 -17281 281 -17211
rect 121 -17321 171 -17281
rect 141 -17341 171 -17321
rect 231 -17321 281 -17281
rect 231 -17341 261 -17321
rect 341 -17381 401 -17121
rect 1 -17391 81 -17381
rect 1 -17451 11 -17391
rect 71 -17401 81 -17391
rect 321 -17391 401 -17381
rect 321 -17401 331 -17391
rect 71 -17451 331 -17401
rect 391 -17451 401 -17391
rect 1 -17461 401 -17451
rect 457 -17041 857 -17031
rect 457 -17101 467 -17041
rect 527 -17091 787 -17041
rect 527 -17101 537 -17091
rect 457 -17111 537 -17101
rect 777 -17101 787 -17091
rect 847 -17101 857 -17041
rect 777 -17111 857 -17101
rect 457 -17381 517 -17111
rect 787 -17121 857 -17111
rect 597 -17171 627 -17151
rect 577 -17211 627 -17171
rect 687 -17171 717 -17151
rect 687 -17211 737 -17171
rect 577 -17281 737 -17211
rect 577 -17321 627 -17281
rect 597 -17341 627 -17321
rect 687 -17321 737 -17281
rect 687 -17341 717 -17321
rect 797 -17381 857 -17121
rect 457 -17391 537 -17381
rect 457 -17451 467 -17391
rect 527 -17401 537 -17391
rect 777 -17391 857 -17381
rect 777 -17401 787 -17391
rect 527 -17451 787 -17401
rect 847 -17451 857 -17391
rect 457 -17461 857 -17451
rect 913 -17041 1313 -17031
rect 913 -17101 923 -17041
rect 983 -17091 1243 -17041
rect 983 -17101 993 -17091
rect 913 -17111 993 -17101
rect 1233 -17101 1243 -17091
rect 1303 -17101 1313 -17041
rect 1233 -17111 1313 -17101
rect 913 -17381 973 -17111
rect 1243 -17121 1313 -17111
rect 1053 -17171 1083 -17151
rect 1033 -17211 1083 -17171
rect 1143 -17171 1173 -17151
rect 1143 -17211 1193 -17171
rect 1033 -17281 1193 -17211
rect 1033 -17321 1083 -17281
rect 1053 -17341 1083 -17321
rect 1143 -17321 1193 -17281
rect 1143 -17341 1173 -17321
rect 1253 -17381 1313 -17121
rect 913 -17391 993 -17381
rect 913 -17451 923 -17391
rect 983 -17401 993 -17391
rect 1233 -17391 1313 -17381
rect 1233 -17401 1243 -17391
rect 983 -17451 1243 -17401
rect 1303 -17451 1313 -17391
rect 913 -17461 1313 -17451
rect 1371 -17041 1771 -17031
rect 1371 -17101 1381 -17041
rect 1441 -17091 1701 -17041
rect 1441 -17101 1451 -17091
rect 1371 -17111 1451 -17101
rect 1691 -17101 1701 -17091
rect 1761 -17101 1771 -17041
rect 1691 -17111 1771 -17101
rect 1371 -17381 1431 -17111
rect 1701 -17121 1771 -17111
rect 1511 -17171 1541 -17151
rect 1491 -17211 1541 -17171
rect 1601 -17171 1631 -17151
rect 1601 -17211 1651 -17171
rect 1491 -17281 1651 -17211
rect 1491 -17321 1541 -17281
rect 1511 -17341 1541 -17321
rect 1601 -17321 1651 -17281
rect 1601 -17341 1631 -17321
rect 1711 -17381 1771 -17121
rect 1371 -17391 1451 -17381
rect 1371 -17451 1381 -17391
rect 1441 -17401 1451 -17391
rect 1691 -17391 1771 -17381
rect 1691 -17401 1701 -17391
rect 1441 -17451 1701 -17401
rect 1761 -17451 1771 -17391
rect 1371 -17461 1771 -17451
rect 1827 -17041 2227 -17031
rect 1827 -17101 1837 -17041
rect 1897 -17091 2157 -17041
rect 1897 -17101 1907 -17091
rect 1827 -17111 1907 -17101
rect 2147 -17101 2157 -17091
rect 2217 -17101 2227 -17041
rect 2147 -17111 2227 -17101
rect 1827 -17381 1887 -17111
rect 2157 -17121 2227 -17111
rect 1967 -17171 1997 -17151
rect 1947 -17211 1997 -17171
rect 2057 -17171 2087 -17151
rect 2057 -17211 2107 -17171
rect 1947 -17281 2107 -17211
rect 1947 -17321 1997 -17281
rect 1967 -17341 1997 -17321
rect 2057 -17321 2107 -17281
rect 2057 -17341 2087 -17321
rect 2167 -17381 2227 -17121
rect 1827 -17391 1907 -17381
rect 1827 -17451 1837 -17391
rect 1897 -17401 1907 -17391
rect 2147 -17391 2227 -17381
rect 2147 -17401 2157 -17391
rect 1897 -17451 2157 -17401
rect 2217 -17451 2227 -17391
rect 1827 -17461 2227 -17451
rect 2283 -17041 2683 -17031
rect 2283 -17101 2293 -17041
rect 2353 -17091 2613 -17041
rect 2353 -17101 2363 -17091
rect 2283 -17111 2363 -17101
rect 2603 -17101 2613 -17091
rect 2673 -17101 2683 -17041
rect 2603 -17111 2683 -17101
rect 2283 -17381 2343 -17111
rect 2613 -17121 2683 -17111
rect 2423 -17171 2453 -17151
rect 2403 -17211 2453 -17171
rect 2513 -17171 2543 -17151
rect 2513 -17211 2563 -17171
rect 2403 -17281 2563 -17211
rect 2403 -17321 2453 -17281
rect 2423 -17341 2453 -17321
rect 2513 -17321 2563 -17281
rect 2513 -17341 2543 -17321
rect 2623 -17381 2683 -17121
rect 2283 -17391 2363 -17381
rect 2283 -17451 2293 -17391
rect 2353 -17401 2363 -17391
rect 2603 -17391 2683 -17381
rect 2603 -17401 2613 -17391
rect 2353 -17451 2613 -17401
rect 2673 -17451 2683 -17391
rect 2283 -17461 2683 -17451
rect 2741 -17041 3141 -17031
rect 2741 -17101 2751 -17041
rect 2811 -17091 3071 -17041
rect 2811 -17101 2821 -17091
rect 2741 -17111 2821 -17101
rect 3061 -17101 3071 -17091
rect 3131 -17101 3141 -17041
rect 3061 -17111 3141 -17101
rect 2741 -17381 2801 -17111
rect 3071 -17121 3141 -17111
rect 2881 -17171 2911 -17151
rect 2861 -17211 2911 -17171
rect 2971 -17171 3001 -17151
rect 2971 -17211 3021 -17171
rect 2861 -17281 3021 -17211
rect 2861 -17321 2911 -17281
rect 2881 -17341 2911 -17321
rect 2971 -17321 3021 -17281
rect 2971 -17341 3001 -17321
rect 3081 -17381 3141 -17121
rect 2741 -17391 2821 -17381
rect 2741 -17451 2751 -17391
rect 2811 -17401 2821 -17391
rect 3061 -17391 3141 -17381
rect 3061 -17401 3071 -17391
rect 2811 -17451 3071 -17401
rect 3131 -17451 3141 -17391
rect 2741 -17461 3141 -17451
rect 3197 -17041 3597 -17031
rect 3197 -17101 3207 -17041
rect 3267 -17091 3527 -17041
rect 3267 -17101 3277 -17091
rect 3197 -17111 3277 -17101
rect 3517 -17101 3527 -17091
rect 3587 -17101 3597 -17041
rect 3517 -17111 3597 -17101
rect 3197 -17381 3257 -17111
rect 3527 -17121 3597 -17111
rect 3337 -17171 3367 -17151
rect 3317 -17211 3367 -17171
rect 3427 -17171 3457 -17151
rect 3427 -17211 3477 -17171
rect 3317 -17281 3477 -17211
rect 3317 -17321 3367 -17281
rect 3337 -17341 3367 -17321
rect 3427 -17321 3477 -17281
rect 3427 -17341 3457 -17321
rect 3537 -17381 3597 -17121
rect 3197 -17391 3277 -17381
rect 3197 -17451 3207 -17391
rect 3267 -17401 3277 -17391
rect 3517 -17391 3597 -17381
rect 3517 -17401 3527 -17391
rect 3267 -17451 3527 -17401
rect 3587 -17451 3597 -17391
rect 3197 -17461 3597 -17451
rect 3653 -17041 4053 -17031
rect 3653 -17101 3663 -17041
rect 3723 -17091 3983 -17041
rect 3723 -17101 3733 -17091
rect 3653 -17111 3733 -17101
rect 3973 -17101 3983 -17091
rect 4043 -17101 4053 -17041
rect 3973 -17111 4053 -17101
rect 3653 -17381 3713 -17111
rect 3983 -17121 4053 -17111
rect 3793 -17171 3823 -17151
rect 3773 -17211 3823 -17171
rect 3883 -17171 3913 -17151
rect 3883 -17211 3933 -17171
rect 3773 -17281 3933 -17211
rect 3773 -17321 3823 -17281
rect 3793 -17341 3823 -17321
rect 3883 -17321 3933 -17281
rect 3883 -17341 3913 -17321
rect 3993 -17381 4053 -17121
rect 3653 -17391 3733 -17381
rect 3653 -17451 3663 -17391
rect 3723 -17401 3733 -17391
rect 3973 -17391 4053 -17381
rect 3973 -17401 3983 -17391
rect 3723 -17451 3983 -17401
rect 4043 -17451 4053 -17391
rect 3653 -17461 4053 -17451
rect 4111 -17041 4511 -17031
rect 4111 -17101 4121 -17041
rect 4181 -17091 4441 -17041
rect 4181 -17101 4191 -17091
rect 4111 -17111 4191 -17101
rect 4431 -17101 4441 -17091
rect 4501 -17101 4511 -17041
rect 4431 -17111 4511 -17101
rect 4111 -17381 4171 -17111
rect 4441 -17121 4511 -17111
rect 4251 -17171 4281 -17151
rect 4231 -17211 4281 -17171
rect 4341 -17171 4371 -17151
rect 4341 -17211 4391 -17171
rect 4231 -17281 4391 -17211
rect 4231 -17321 4281 -17281
rect 4251 -17341 4281 -17321
rect 4341 -17321 4391 -17281
rect 4341 -17341 4371 -17321
rect 4451 -17381 4511 -17121
rect 4111 -17391 4191 -17381
rect 4111 -17451 4121 -17391
rect 4181 -17401 4191 -17391
rect 4431 -17391 4511 -17381
rect 4431 -17401 4441 -17391
rect 4181 -17451 4441 -17401
rect 4501 -17451 4511 -17391
rect 4111 -17461 4511 -17451
rect 4567 -17041 4967 -17031
rect 4567 -17101 4577 -17041
rect 4637 -17091 4897 -17041
rect 4637 -17101 4647 -17091
rect 4567 -17111 4647 -17101
rect 4887 -17101 4897 -17091
rect 4957 -17101 4967 -17041
rect 4887 -17111 4967 -17101
rect 4567 -17381 4627 -17111
rect 4897 -17121 4967 -17111
rect 4707 -17171 4737 -17151
rect 4687 -17211 4737 -17171
rect 4797 -17171 4827 -17151
rect 4797 -17211 4847 -17171
rect 4687 -17281 4847 -17211
rect 4687 -17321 4737 -17281
rect 4707 -17341 4737 -17321
rect 4797 -17321 4847 -17281
rect 4797 -17341 4827 -17321
rect 4907 -17381 4967 -17121
rect 4567 -17391 4647 -17381
rect 4567 -17451 4577 -17391
rect 4637 -17401 4647 -17391
rect 4887 -17391 4967 -17381
rect 4887 -17401 4897 -17391
rect 4637 -17451 4897 -17401
rect 4957 -17451 4967 -17391
rect 4567 -17461 4967 -17451
rect 5023 -17041 5423 -17031
rect 5023 -17101 5033 -17041
rect 5093 -17091 5353 -17041
rect 5093 -17101 5103 -17091
rect 5023 -17111 5103 -17101
rect 5343 -17101 5353 -17091
rect 5413 -17101 5423 -17041
rect 5343 -17111 5423 -17101
rect 5023 -17381 5083 -17111
rect 5353 -17121 5423 -17111
rect 5163 -17171 5193 -17151
rect 5143 -17211 5193 -17171
rect 5253 -17171 5283 -17151
rect 5253 -17211 5303 -17171
rect 5143 -17281 5303 -17211
rect 5143 -17321 5193 -17281
rect 5163 -17341 5193 -17321
rect 5253 -17321 5303 -17281
rect 5253 -17341 5283 -17321
rect 5363 -17381 5423 -17121
rect 5023 -17391 5103 -17381
rect 5023 -17451 5033 -17391
rect 5093 -17401 5103 -17391
rect 5343 -17391 5423 -17381
rect 5343 -17401 5353 -17391
rect 5093 -17451 5353 -17401
rect 5413 -17451 5423 -17391
rect 5023 -17461 5423 -17451
rect 5481 -17041 5881 -17031
rect 5481 -17101 5491 -17041
rect 5551 -17091 5811 -17041
rect 5551 -17101 5561 -17091
rect 5481 -17111 5561 -17101
rect 5801 -17101 5811 -17091
rect 5871 -17101 5881 -17041
rect 5801 -17111 5881 -17101
rect 5481 -17381 5541 -17111
rect 5811 -17121 5881 -17111
rect 5621 -17171 5651 -17151
rect 5601 -17211 5651 -17171
rect 5711 -17171 5741 -17151
rect 5711 -17211 5761 -17171
rect 5601 -17281 5761 -17211
rect 5601 -17321 5651 -17281
rect 5621 -17341 5651 -17321
rect 5711 -17321 5761 -17281
rect 5711 -17341 5741 -17321
rect 5821 -17381 5881 -17121
rect 5481 -17391 5561 -17381
rect 5481 -17451 5491 -17391
rect 5551 -17401 5561 -17391
rect 5801 -17391 5881 -17381
rect 5801 -17401 5811 -17391
rect 5551 -17451 5811 -17401
rect 5871 -17451 5881 -17391
rect 5481 -17461 5881 -17451
rect 5937 -17041 6337 -17031
rect 5937 -17101 5947 -17041
rect 6007 -17091 6267 -17041
rect 6007 -17101 6017 -17091
rect 5937 -17111 6017 -17101
rect 6257 -17101 6267 -17091
rect 6327 -17101 6337 -17041
rect 6257 -17111 6337 -17101
rect 5937 -17381 5997 -17111
rect 6267 -17121 6337 -17111
rect 6077 -17171 6107 -17151
rect 6057 -17211 6107 -17171
rect 6167 -17171 6197 -17151
rect 6167 -17211 6217 -17171
rect 6057 -17281 6217 -17211
rect 6057 -17321 6107 -17281
rect 6077 -17341 6107 -17321
rect 6167 -17321 6217 -17281
rect 6167 -17341 6197 -17321
rect 6277 -17381 6337 -17121
rect 5937 -17391 6017 -17381
rect 5937 -17451 5947 -17391
rect 6007 -17401 6017 -17391
rect 6257 -17391 6337 -17381
rect 6257 -17401 6267 -17391
rect 6007 -17451 6267 -17401
rect 6327 -17451 6337 -17391
rect 5937 -17461 6337 -17451
rect 6393 -17041 6793 -17031
rect 6393 -17101 6403 -17041
rect 6463 -17091 6723 -17041
rect 6463 -17101 6473 -17091
rect 6393 -17111 6473 -17101
rect 6713 -17101 6723 -17091
rect 6783 -17101 6793 -17041
rect 6713 -17111 6793 -17101
rect 6393 -17381 6453 -17111
rect 6723 -17121 6793 -17111
rect 6533 -17171 6563 -17151
rect 6513 -17211 6563 -17171
rect 6623 -17171 6653 -17151
rect 6623 -17211 6673 -17171
rect 6513 -17281 6673 -17211
rect 6513 -17321 6563 -17281
rect 6533 -17341 6563 -17321
rect 6623 -17321 6673 -17281
rect 6623 -17341 6653 -17321
rect 6733 -17381 6793 -17121
rect 6393 -17391 6473 -17381
rect 6393 -17451 6403 -17391
rect 6463 -17401 6473 -17391
rect 6713 -17391 6793 -17381
rect 6713 -17401 6723 -17391
rect 6463 -17451 6723 -17401
rect 6783 -17451 6793 -17391
rect 6393 -17461 6793 -17451
rect 6851 -17041 7251 -17031
rect 6851 -17101 6861 -17041
rect 6921 -17091 7181 -17041
rect 6921 -17101 6931 -17091
rect 6851 -17111 6931 -17101
rect 7171 -17101 7181 -17091
rect 7241 -17101 7251 -17041
rect 7171 -17111 7251 -17101
rect 6851 -17381 6911 -17111
rect 7181 -17121 7251 -17111
rect 6991 -17171 7021 -17151
rect 6971 -17211 7021 -17171
rect 7081 -17171 7111 -17151
rect 7081 -17211 7131 -17171
rect 6971 -17281 7131 -17211
rect 6971 -17321 7021 -17281
rect 6991 -17341 7021 -17321
rect 7081 -17321 7131 -17281
rect 7081 -17341 7111 -17321
rect 7191 -17381 7251 -17121
rect 6851 -17391 6931 -17381
rect 6851 -17451 6861 -17391
rect 6921 -17401 6931 -17391
rect 7171 -17391 7251 -17381
rect 7171 -17401 7181 -17391
rect 6921 -17451 7181 -17401
rect 7241 -17451 7251 -17391
rect 6851 -17461 7251 -17451
rect 7307 -17041 7707 -17031
rect 7307 -17101 7317 -17041
rect 7377 -17091 7637 -17041
rect 7377 -17101 7387 -17091
rect 7307 -17111 7387 -17101
rect 7627 -17101 7637 -17091
rect 7697 -17101 7707 -17041
rect 7627 -17111 7707 -17101
rect 7307 -17381 7367 -17111
rect 7637 -17121 7707 -17111
rect 7447 -17171 7477 -17151
rect 7427 -17211 7477 -17171
rect 7537 -17171 7567 -17151
rect 7537 -17211 7587 -17171
rect 7427 -17281 7587 -17211
rect 7427 -17321 7477 -17281
rect 7447 -17341 7477 -17321
rect 7537 -17321 7587 -17281
rect 7537 -17341 7567 -17321
rect 7647 -17381 7707 -17121
rect 7307 -17391 7387 -17381
rect 7307 -17451 7317 -17391
rect 7377 -17401 7387 -17391
rect 7627 -17391 7707 -17381
rect 7627 -17401 7637 -17391
rect 7377 -17451 7637 -17401
rect 7697 -17451 7707 -17391
rect 7307 -17461 7707 -17451
rect 7763 -17041 8163 -17031
rect 7763 -17101 7773 -17041
rect 7833 -17091 8093 -17041
rect 7833 -17101 7843 -17091
rect 7763 -17111 7843 -17101
rect 8083 -17101 8093 -17091
rect 8153 -17101 8163 -17041
rect 8083 -17111 8163 -17101
rect 7763 -17381 7823 -17111
rect 8093 -17121 8163 -17111
rect 7903 -17171 7933 -17151
rect 7883 -17211 7933 -17171
rect 7993 -17171 8023 -17151
rect 7993 -17211 8043 -17171
rect 7883 -17281 8043 -17211
rect 7883 -17321 7933 -17281
rect 7903 -17341 7933 -17321
rect 7993 -17321 8043 -17281
rect 7993 -17341 8023 -17321
rect 8103 -17381 8163 -17121
rect 7763 -17391 7843 -17381
rect 7763 -17451 7773 -17391
rect 7833 -17401 7843 -17391
rect 8083 -17391 8163 -17381
rect 8083 -17401 8093 -17391
rect 7833 -17451 8093 -17401
rect 8153 -17451 8163 -17391
rect 7763 -17461 8163 -17451
rect 8237 -17041 8637 -17031
rect 8237 -17101 8247 -17041
rect 8307 -17091 8567 -17041
rect 8307 -17101 8317 -17091
rect 8237 -17111 8317 -17101
rect 8557 -17101 8567 -17091
rect 8627 -17101 8637 -17041
rect 8557 -17111 8637 -17101
rect 8237 -17381 8297 -17111
rect 8567 -17121 8637 -17111
rect 8377 -17171 8407 -17151
rect 8357 -17211 8407 -17171
rect 8467 -17171 8497 -17151
rect 8467 -17211 8517 -17171
rect 8357 -17281 8517 -17211
rect 8357 -17321 8407 -17281
rect 8377 -17341 8407 -17321
rect 8467 -17321 8517 -17281
rect 8467 -17341 8497 -17321
rect 8577 -17381 8637 -17121
rect 8237 -17391 8317 -17381
rect 8237 -17451 8247 -17391
rect 8307 -17401 8317 -17391
rect 8557 -17391 8637 -17381
rect 8557 -17401 8567 -17391
rect 8307 -17451 8567 -17401
rect 8627 -17451 8637 -17391
rect 8237 -17461 8637 -17451
rect 8693 -17041 9093 -17031
rect 8693 -17101 8703 -17041
rect 8763 -17091 9023 -17041
rect 8763 -17101 8773 -17091
rect 8693 -17111 8773 -17101
rect 9013 -17101 9023 -17091
rect 9083 -17101 9093 -17041
rect 9013 -17111 9093 -17101
rect 8693 -17381 8753 -17111
rect 9023 -17121 9093 -17111
rect 8833 -17171 8863 -17151
rect 8813 -17211 8863 -17171
rect 8923 -17171 8953 -17151
rect 8923 -17211 8973 -17171
rect 8813 -17281 8973 -17211
rect 8813 -17321 8863 -17281
rect 8833 -17341 8863 -17321
rect 8923 -17321 8973 -17281
rect 8923 -17341 8953 -17321
rect 9033 -17381 9093 -17121
rect 8693 -17391 8773 -17381
rect 8693 -17451 8703 -17391
rect 8763 -17401 8773 -17391
rect 9013 -17391 9093 -17381
rect 9013 -17401 9023 -17391
rect 8763 -17451 9023 -17401
rect 9083 -17451 9093 -17391
rect 8693 -17461 9093 -17451
rect 9151 -17041 9551 -17031
rect 9151 -17101 9161 -17041
rect 9221 -17091 9481 -17041
rect 9221 -17101 9231 -17091
rect 9151 -17111 9231 -17101
rect 9471 -17101 9481 -17091
rect 9541 -17101 9551 -17041
rect 9471 -17111 9551 -17101
rect 9151 -17381 9211 -17111
rect 9481 -17121 9551 -17111
rect 9291 -17171 9321 -17151
rect 9271 -17211 9321 -17171
rect 9381 -17171 9411 -17151
rect 9381 -17211 9431 -17171
rect 9271 -17281 9431 -17211
rect 9271 -17321 9321 -17281
rect 9291 -17341 9321 -17321
rect 9381 -17321 9431 -17281
rect 9381 -17341 9411 -17321
rect 9491 -17381 9551 -17121
rect 9151 -17391 9231 -17381
rect 9151 -17451 9161 -17391
rect 9221 -17401 9231 -17391
rect 9471 -17391 9551 -17381
rect 9471 -17401 9481 -17391
rect 9221 -17451 9481 -17401
rect 9541 -17451 9551 -17391
rect 9151 -17461 9551 -17451
rect 9607 -17041 10007 -17031
rect 9607 -17101 9617 -17041
rect 9677 -17091 9937 -17041
rect 9677 -17101 9687 -17091
rect 9607 -17111 9687 -17101
rect 9927 -17101 9937 -17091
rect 9997 -17101 10007 -17041
rect 9927 -17111 10007 -17101
rect 9607 -17381 9667 -17111
rect 9937 -17121 10007 -17111
rect 9747 -17171 9777 -17151
rect 9727 -17211 9777 -17171
rect 9837 -17171 9867 -17151
rect 9837 -17211 9887 -17171
rect 9727 -17281 9887 -17211
rect 9727 -17321 9777 -17281
rect 9747 -17341 9777 -17321
rect 9837 -17321 9887 -17281
rect 9837 -17341 9867 -17321
rect 9947 -17381 10007 -17121
rect 9607 -17391 9687 -17381
rect 9607 -17451 9617 -17391
rect 9677 -17401 9687 -17391
rect 9927 -17391 10007 -17381
rect 9927 -17401 9937 -17391
rect 9677 -17451 9937 -17401
rect 9997 -17451 10007 -17391
rect 9607 -17461 10007 -17451
rect 10063 -17041 10463 -17031
rect 10063 -17101 10073 -17041
rect 10133 -17091 10393 -17041
rect 10133 -17101 10143 -17091
rect 10063 -17111 10143 -17101
rect 10383 -17101 10393 -17091
rect 10453 -17101 10463 -17041
rect 10383 -17111 10463 -17101
rect 10063 -17381 10123 -17111
rect 10393 -17121 10463 -17111
rect 10203 -17171 10233 -17151
rect 10183 -17211 10233 -17171
rect 10293 -17171 10323 -17151
rect 10293 -17211 10343 -17171
rect 10183 -17281 10343 -17211
rect 10183 -17321 10233 -17281
rect 10203 -17341 10233 -17321
rect 10293 -17321 10343 -17281
rect 10293 -17341 10323 -17321
rect 10403 -17381 10463 -17121
rect 10063 -17391 10143 -17381
rect 10063 -17451 10073 -17391
rect 10133 -17401 10143 -17391
rect 10383 -17391 10463 -17381
rect 10383 -17401 10393 -17391
rect 10133 -17451 10393 -17401
rect 10453 -17451 10463 -17391
rect 10063 -17461 10463 -17451
rect 10521 -17041 10921 -17031
rect 10521 -17101 10531 -17041
rect 10591 -17091 10851 -17041
rect 10591 -17101 10601 -17091
rect 10521 -17111 10601 -17101
rect 10841 -17101 10851 -17091
rect 10911 -17101 10921 -17041
rect 10841 -17111 10921 -17101
rect 10521 -17381 10581 -17111
rect 10851 -17121 10921 -17111
rect 10661 -17171 10691 -17151
rect 10641 -17211 10691 -17171
rect 10751 -17171 10781 -17151
rect 10751 -17211 10801 -17171
rect 10641 -17281 10801 -17211
rect 10641 -17321 10691 -17281
rect 10661 -17341 10691 -17321
rect 10751 -17321 10801 -17281
rect 10751 -17341 10781 -17321
rect 10861 -17381 10921 -17121
rect 10521 -17391 10601 -17381
rect 10521 -17451 10531 -17391
rect 10591 -17401 10601 -17391
rect 10841 -17391 10921 -17381
rect 10841 -17401 10851 -17391
rect 10591 -17451 10851 -17401
rect 10911 -17451 10921 -17391
rect 10521 -17461 10921 -17451
rect 10977 -17041 11377 -17031
rect 10977 -17101 10987 -17041
rect 11047 -17091 11307 -17041
rect 11047 -17101 11057 -17091
rect 10977 -17111 11057 -17101
rect 11297 -17101 11307 -17091
rect 11367 -17101 11377 -17041
rect 11297 -17111 11377 -17101
rect 10977 -17381 11037 -17111
rect 11307 -17121 11377 -17111
rect 11117 -17171 11147 -17151
rect 11097 -17211 11147 -17171
rect 11207 -17171 11237 -17151
rect 11207 -17211 11257 -17171
rect 11097 -17281 11257 -17211
rect 11097 -17321 11147 -17281
rect 11117 -17341 11147 -17321
rect 11207 -17321 11257 -17281
rect 11207 -17341 11237 -17321
rect 11317 -17381 11377 -17121
rect 10977 -17391 11057 -17381
rect 10977 -17451 10987 -17391
rect 11047 -17401 11057 -17391
rect 11297 -17391 11377 -17381
rect 11297 -17401 11307 -17391
rect 11047 -17451 11307 -17401
rect 11367 -17451 11377 -17391
rect 10977 -17461 11377 -17451
rect 11433 -17041 11833 -17031
rect 11433 -17101 11443 -17041
rect 11503 -17091 11763 -17041
rect 11503 -17101 11513 -17091
rect 11433 -17111 11513 -17101
rect 11753 -17101 11763 -17091
rect 11823 -17101 11833 -17041
rect 11753 -17111 11833 -17101
rect 11433 -17381 11493 -17111
rect 11763 -17121 11833 -17111
rect 11573 -17171 11603 -17151
rect 11553 -17211 11603 -17171
rect 11663 -17171 11693 -17151
rect 11663 -17211 11713 -17171
rect 11553 -17281 11713 -17211
rect 11553 -17321 11603 -17281
rect 11573 -17341 11603 -17321
rect 11663 -17321 11713 -17281
rect 11663 -17341 11693 -17321
rect 11773 -17381 11833 -17121
rect 11433 -17391 11513 -17381
rect 11433 -17451 11443 -17391
rect 11503 -17401 11513 -17391
rect 11753 -17391 11833 -17381
rect 11753 -17401 11763 -17391
rect 11503 -17451 11763 -17401
rect 11823 -17451 11833 -17391
rect 11433 -17461 11833 -17451
rect 11891 -17041 12291 -17031
rect 11891 -17101 11901 -17041
rect 11961 -17091 12221 -17041
rect 11961 -17101 11971 -17091
rect 11891 -17111 11971 -17101
rect 12211 -17101 12221 -17091
rect 12281 -17101 12291 -17041
rect 12211 -17111 12291 -17101
rect 11891 -17381 11951 -17111
rect 12221 -17121 12291 -17111
rect 12031 -17171 12061 -17151
rect 12011 -17211 12061 -17171
rect 12121 -17171 12151 -17151
rect 12121 -17211 12171 -17171
rect 12011 -17281 12171 -17211
rect 12011 -17321 12061 -17281
rect 12031 -17341 12061 -17321
rect 12121 -17321 12171 -17281
rect 12121 -17341 12151 -17321
rect 12231 -17381 12291 -17121
rect 11891 -17391 11971 -17381
rect 11891 -17451 11901 -17391
rect 11961 -17401 11971 -17391
rect 12211 -17391 12291 -17381
rect 12211 -17401 12221 -17391
rect 11961 -17451 12221 -17401
rect 12281 -17451 12291 -17391
rect 11891 -17461 12291 -17451
rect 12347 -17041 12747 -17031
rect 12347 -17101 12357 -17041
rect 12417 -17091 12677 -17041
rect 12417 -17101 12427 -17091
rect 12347 -17111 12427 -17101
rect 12667 -17101 12677 -17091
rect 12737 -17101 12747 -17041
rect 12667 -17111 12747 -17101
rect 12347 -17381 12407 -17111
rect 12677 -17121 12747 -17111
rect 12487 -17171 12517 -17151
rect 12467 -17211 12517 -17171
rect 12577 -17171 12607 -17151
rect 12577 -17211 12627 -17171
rect 12467 -17281 12627 -17211
rect 12467 -17321 12517 -17281
rect 12487 -17341 12517 -17321
rect 12577 -17321 12627 -17281
rect 12577 -17341 12607 -17321
rect 12687 -17381 12747 -17121
rect 12347 -17391 12427 -17381
rect 12347 -17451 12357 -17391
rect 12417 -17401 12427 -17391
rect 12667 -17391 12747 -17381
rect 12667 -17401 12677 -17391
rect 12417 -17451 12677 -17401
rect 12737 -17451 12747 -17391
rect 12347 -17461 12747 -17451
rect 12803 -17041 13203 -17031
rect 12803 -17101 12813 -17041
rect 12873 -17091 13133 -17041
rect 12873 -17101 12883 -17091
rect 12803 -17111 12883 -17101
rect 13123 -17101 13133 -17091
rect 13193 -17101 13203 -17041
rect 13123 -17111 13203 -17101
rect 12803 -17381 12863 -17111
rect 13133 -17121 13203 -17111
rect 12943 -17171 12973 -17151
rect 12923 -17211 12973 -17171
rect 13033 -17171 13063 -17151
rect 13033 -17211 13083 -17171
rect 12923 -17281 13083 -17211
rect 12923 -17321 12973 -17281
rect 12943 -17341 12973 -17321
rect 13033 -17321 13083 -17281
rect 13033 -17341 13063 -17321
rect 13143 -17381 13203 -17121
rect 12803 -17391 12883 -17381
rect 12803 -17451 12813 -17391
rect 12873 -17401 12883 -17391
rect 13123 -17391 13203 -17381
rect 13123 -17401 13133 -17391
rect 12873 -17451 13133 -17401
rect 13193 -17451 13203 -17391
rect 12803 -17461 13203 -17451
rect 13261 -17041 13661 -17031
rect 13261 -17101 13271 -17041
rect 13331 -17091 13591 -17041
rect 13331 -17101 13341 -17091
rect 13261 -17111 13341 -17101
rect 13581 -17101 13591 -17091
rect 13651 -17101 13661 -17041
rect 13581 -17111 13661 -17101
rect 13261 -17381 13321 -17111
rect 13591 -17121 13661 -17111
rect 13401 -17171 13431 -17151
rect 13381 -17211 13431 -17171
rect 13491 -17171 13521 -17151
rect 13491 -17211 13541 -17171
rect 13381 -17281 13541 -17211
rect 13381 -17321 13431 -17281
rect 13401 -17341 13431 -17321
rect 13491 -17321 13541 -17281
rect 13491 -17341 13521 -17321
rect 13601 -17381 13661 -17121
rect 13261 -17391 13341 -17381
rect 13261 -17451 13271 -17391
rect 13331 -17401 13341 -17391
rect 13581 -17391 13661 -17381
rect 13581 -17401 13591 -17391
rect 13331 -17451 13591 -17401
rect 13651 -17451 13661 -17391
rect 13261 -17461 13661 -17451
rect 13717 -17041 14117 -17031
rect 13717 -17101 13727 -17041
rect 13787 -17091 14047 -17041
rect 13787 -17101 13797 -17091
rect 13717 -17111 13797 -17101
rect 14037 -17101 14047 -17091
rect 14107 -17101 14117 -17041
rect 14037 -17111 14117 -17101
rect 13717 -17381 13777 -17111
rect 14047 -17121 14117 -17111
rect 13857 -17171 13887 -17151
rect 13837 -17211 13887 -17171
rect 13947 -17171 13977 -17151
rect 13947 -17211 13997 -17171
rect 13837 -17281 13997 -17211
rect 13837 -17321 13887 -17281
rect 13857 -17341 13887 -17321
rect 13947 -17321 13997 -17281
rect 13947 -17341 13977 -17321
rect 14057 -17381 14117 -17121
rect 13717 -17391 13797 -17381
rect 13717 -17451 13727 -17391
rect 13787 -17401 13797 -17391
rect 14037 -17391 14117 -17381
rect 14037 -17401 14047 -17391
rect 13787 -17451 14047 -17401
rect 14107 -17451 14117 -17391
rect 13717 -17461 14117 -17451
rect 14173 -17041 14573 -17031
rect 14173 -17101 14183 -17041
rect 14243 -17091 14503 -17041
rect 14243 -17101 14253 -17091
rect 14173 -17111 14253 -17101
rect 14493 -17101 14503 -17091
rect 14563 -17101 14573 -17041
rect 14493 -17111 14573 -17101
rect 14173 -17381 14233 -17111
rect 14503 -17121 14573 -17111
rect 14313 -17171 14343 -17151
rect 14293 -17211 14343 -17171
rect 14403 -17171 14433 -17151
rect 14403 -17211 14453 -17171
rect 14293 -17281 14453 -17211
rect 14293 -17321 14343 -17281
rect 14313 -17341 14343 -17321
rect 14403 -17321 14453 -17281
rect 14403 -17341 14433 -17321
rect 14513 -17381 14573 -17121
rect 14173 -17391 14253 -17381
rect 14173 -17451 14183 -17391
rect 14243 -17401 14253 -17391
rect 14493 -17391 14573 -17381
rect 14493 -17401 14503 -17391
rect 14243 -17451 14503 -17401
rect 14563 -17451 14573 -17391
rect 14173 -17461 14573 -17451
rect 14631 -17041 15031 -17031
rect 14631 -17101 14641 -17041
rect 14701 -17091 14961 -17041
rect 14701 -17101 14711 -17091
rect 14631 -17111 14711 -17101
rect 14951 -17101 14961 -17091
rect 15021 -17101 15031 -17041
rect 14951 -17111 15031 -17101
rect 14631 -17381 14691 -17111
rect 14961 -17121 15031 -17111
rect 14771 -17171 14801 -17151
rect 14751 -17211 14801 -17171
rect 14861 -17171 14891 -17151
rect 14861 -17211 14911 -17171
rect 14751 -17281 14911 -17211
rect 14751 -17321 14801 -17281
rect 14771 -17341 14801 -17321
rect 14861 -17321 14911 -17281
rect 14861 -17341 14891 -17321
rect 14971 -17381 15031 -17121
rect 14631 -17391 14711 -17381
rect 14631 -17451 14641 -17391
rect 14701 -17401 14711 -17391
rect 14951 -17391 15031 -17381
rect 14951 -17401 14961 -17391
rect 14701 -17451 14961 -17401
rect 15021 -17451 15031 -17391
rect 14631 -17461 15031 -17451
rect 15087 -17041 15487 -17031
rect 15087 -17101 15097 -17041
rect 15157 -17091 15417 -17041
rect 15157 -17101 15167 -17091
rect 15087 -17111 15167 -17101
rect 15407 -17101 15417 -17091
rect 15477 -17101 15487 -17041
rect 15407 -17111 15487 -17101
rect 15087 -17381 15147 -17111
rect 15417 -17121 15487 -17111
rect 15227 -17171 15257 -17151
rect 15207 -17211 15257 -17171
rect 15317 -17171 15347 -17151
rect 15317 -17211 15367 -17171
rect 15207 -17281 15367 -17211
rect 15207 -17321 15257 -17281
rect 15227 -17341 15257 -17321
rect 15317 -17321 15367 -17281
rect 15317 -17341 15347 -17321
rect 15427 -17381 15487 -17121
rect 15087 -17391 15167 -17381
rect 15087 -17451 15097 -17391
rect 15157 -17401 15167 -17391
rect 15407 -17391 15487 -17381
rect 15407 -17401 15417 -17391
rect 15157 -17451 15417 -17401
rect 15477 -17451 15487 -17391
rect 15087 -17461 15487 -17451
rect 1 -17533 401 -17523
rect 1 -17593 11 -17533
rect 71 -17583 331 -17533
rect 71 -17593 81 -17583
rect 1 -17603 81 -17593
rect 321 -17593 331 -17583
rect 391 -17593 401 -17533
rect 321 -17603 401 -17593
rect 1 -17873 61 -17603
rect 331 -17613 401 -17603
rect 141 -17663 171 -17643
rect 121 -17703 171 -17663
rect 231 -17663 261 -17643
rect 231 -17703 281 -17663
rect 121 -17773 281 -17703
rect 121 -17813 171 -17773
rect 141 -17833 171 -17813
rect 231 -17813 281 -17773
rect 231 -17833 261 -17813
rect 341 -17873 401 -17613
rect 1 -17883 81 -17873
rect 1 -17943 11 -17883
rect 71 -17893 81 -17883
rect 321 -17883 401 -17873
rect 321 -17893 331 -17883
rect 71 -17943 331 -17893
rect 391 -17943 401 -17883
rect 1 -17953 401 -17943
rect 457 -17533 857 -17523
rect 457 -17593 467 -17533
rect 527 -17583 787 -17533
rect 527 -17593 537 -17583
rect 457 -17603 537 -17593
rect 777 -17593 787 -17583
rect 847 -17593 857 -17533
rect 777 -17603 857 -17593
rect 457 -17873 517 -17603
rect 787 -17613 857 -17603
rect 597 -17663 627 -17643
rect 577 -17703 627 -17663
rect 687 -17663 717 -17643
rect 687 -17703 737 -17663
rect 577 -17773 737 -17703
rect 577 -17813 627 -17773
rect 597 -17833 627 -17813
rect 687 -17813 737 -17773
rect 687 -17833 717 -17813
rect 797 -17873 857 -17613
rect 457 -17883 537 -17873
rect 457 -17943 467 -17883
rect 527 -17893 537 -17883
rect 777 -17883 857 -17873
rect 777 -17893 787 -17883
rect 527 -17943 787 -17893
rect 847 -17943 857 -17883
rect 457 -17953 857 -17943
rect 913 -17533 1313 -17523
rect 913 -17593 923 -17533
rect 983 -17583 1243 -17533
rect 983 -17593 993 -17583
rect 913 -17603 993 -17593
rect 1233 -17593 1243 -17583
rect 1303 -17593 1313 -17533
rect 1233 -17603 1313 -17593
rect 913 -17873 973 -17603
rect 1243 -17613 1313 -17603
rect 1053 -17663 1083 -17643
rect 1033 -17703 1083 -17663
rect 1143 -17663 1173 -17643
rect 1143 -17703 1193 -17663
rect 1033 -17773 1193 -17703
rect 1033 -17813 1083 -17773
rect 1053 -17833 1083 -17813
rect 1143 -17813 1193 -17773
rect 1143 -17833 1173 -17813
rect 1253 -17873 1313 -17613
rect 913 -17883 993 -17873
rect 913 -17943 923 -17883
rect 983 -17893 993 -17883
rect 1233 -17883 1313 -17873
rect 1233 -17893 1243 -17883
rect 983 -17943 1243 -17893
rect 1303 -17943 1313 -17883
rect 913 -17953 1313 -17943
rect 1371 -17533 1771 -17523
rect 1371 -17593 1381 -17533
rect 1441 -17583 1701 -17533
rect 1441 -17593 1451 -17583
rect 1371 -17603 1451 -17593
rect 1691 -17593 1701 -17583
rect 1761 -17593 1771 -17533
rect 1691 -17603 1771 -17593
rect 1371 -17873 1431 -17603
rect 1701 -17613 1771 -17603
rect 1511 -17663 1541 -17643
rect 1491 -17703 1541 -17663
rect 1601 -17663 1631 -17643
rect 1601 -17703 1651 -17663
rect 1491 -17773 1651 -17703
rect 1491 -17813 1541 -17773
rect 1511 -17833 1541 -17813
rect 1601 -17813 1651 -17773
rect 1601 -17833 1631 -17813
rect 1711 -17873 1771 -17613
rect 1371 -17883 1451 -17873
rect 1371 -17943 1381 -17883
rect 1441 -17893 1451 -17883
rect 1691 -17883 1771 -17873
rect 1691 -17893 1701 -17883
rect 1441 -17943 1701 -17893
rect 1761 -17943 1771 -17883
rect 1371 -17953 1771 -17943
rect 1827 -17533 2227 -17523
rect 1827 -17593 1837 -17533
rect 1897 -17583 2157 -17533
rect 1897 -17593 1907 -17583
rect 1827 -17603 1907 -17593
rect 2147 -17593 2157 -17583
rect 2217 -17593 2227 -17533
rect 2147 -17603 2227 -17593
rect 1827 -17873 1887 -17603
rect 2157 -17613 2227 -17603
rect 1967 -17663 1997 -17643
rect 1947 -17703 1997 -17663
rect 2057 -17663 2087 -17643
rect 2057 -17703 2107 -17663
rect 1947 -17773 2107 -17703
rect 1947 -17813 1997 -17773
rect 1967 -17833 1997 -17813
rect 2057 -17813 2107 -17773
rect 2057 -17833 2087 -17813
rect 2167 -17873 2227 -17613
rect 1827 -17883 1907 -17873
rect 1827 -17943 1837 -17883
rect 1897 -17893 1907 -17883
rect 2147 -17883 2227 -17873
rect 2147 -17893 2157 -17883
rect 1897 -17943 2157 -17893
rect 2217 -17943 2227 -17883
rect 1827 -17953 2227 -17943
rect 2283 -17533 2683 -17523
rect 2283 -17593 2293 -17533
rect 2353 -17583 2613 -17533
rect 2353 -17593 2363 -17583
rect 2283 -17603 2363 -17593
rect 2603 -17593 2613 -17583
rect 2673 -17593 2683 -17533
rect 2603 -17603 2683 -17593
rect 2283 -17873 2343 -17603
rect 2613 -17613 2683 -17603
rect 2423 -17663 2453 -17643
rect 2403 -17703 2453 -17663
rect 2513 -17663 2543 -17643
rect 2513 -17703 2563 -17663
rect 2403 -17773 2563 -17703
rect 2403 -17813 2453 -17773
rect 2423 -17833 2453 -17813
rect 2513 -17813 2563 -17773
rect 2513 -17833 2543 -17813
rect 2623 -17873 2683 -17613
rect 2283 -17883 2363 -17873
rect 2283 -17943 2293 -17883
rect 2353 -17893 2363 -17883
rect 2603 -17883 2683 -17873
rect 2603 -17893 2613 -17883
rect 2353 -17943 2613 -17893
rect 2673 -17943 2683 -17883
rect 2283 -17953 2683 -17943
rect 2741 -17533 3141 -17523
rect 2741 -17593 2751 -17533
rect 2811 -17583 3071 -17533
rect 2811 -17593 2821 -17583
rect 2741 -17603 2821 -17593
rect 3061 -17593 3071 -17583
rect 3131 -17593 3141 -17533
rect 3061 -17603 3141 -17593
rect 2741 -17873 2801 -17603
rect 3071 -17613 3141 -17603
rect 2881 -17663 2911 -17643
rect 2861 -17703 2911 -17663
rect 2971 -17663 3001 -17643
rect 2971 -17703 3021 -17663
rect 2861 -17773 3021 -17703
rect 2861 -17813 2911 -17773
rect 2881 -17833 2911 -17813
rect 2971 -17813 3021 -17773
rect 2971 -17833 3001 -17813
rect 3081 -17873 3141 -17613
rect 2741 -17883 2821 -17873
rect 2741 -17943 2751 -17883
rect 2811 -17893 2821 -17883
rect 3061 -17883 3141 -17873
rect 3061 -17893 3071 -17883
rect 2811 -17943 3071 -17893
rect 3131 -17943 3141 -17883
rect 2741 -17953 3141 -17943
rect 3197 -17533 3597 -17523
rect 3197 -17593 3207 -17533
rect 3267 -17583 3527 -17533
rect 3267 -17593 3277 -17583
rect 3197 -17603 3277 -17593
rect 3517 -17593 3527 -17583
rect 3587 -17593 3597 -17533
rect 3517 -17603 3597 -17593
rect 3197 -17873 3257 -17603
rect 3527 -17613 3597 -17603
rect 3337 -17663 3367 -17643
rect 3317 -17703 3367 -17663
rect 3427 -17663 3457 -17643
rect 3427 -17703 3477 -17663
rect 3317 -17773 3477 -17703
rect 3317 -17813 3367 -17773
rect 3337 -17833 3367 -17813
rect 3427 -17813 3477 -17773
rect 3427 -17833 3457 -17813
rect 3537 -17873 3597 -17613
rect 3197 -17883 3277 -17873
rect 3197 -17943 3207 -17883
rect 3267 -17893 3277 -17883
rect 3517 -17883 3597 -17873
rect 3517 -17893 3527 -17883
rect 3267 -17943 3527 -17893
rect 3587 -17943 3597 -17883
rect 3197 -17953 3597 -17943
rect 3653 -17533 4053 -17523
rect 3653 -17593 3663 -17533
rect 3723 -17583 3983 -17533
rect 3723 -17593 3733 -17583
rect 3653 -17603 3733 -17593
rect 3973 -17593 3983 -17583
rect 4043 -17593 4053 -17533
rect 3973 -17603 4053 -17593
rect 3653 -17873 3713 -17603
rect 3983 -17613 4053 -17603
rect 3793 -17663 3823 -17643
rect 3773 -17703 3823 -17663
rect 3883 -17663 3913 -17643
rect 3883 -17703 3933 -17663
rect 3773 -17773 3933 -17703
rect 3773 -17813 3823 -17773
rect 3793 -17833 3823 -17813
rect 3883 -17813 3933 -17773
rect 3883 -17833 3913 -17813
rect 3993 -17873 4053 -17613
rect 3653 -17883 3733 -17873
rect 3653 -17943 3663 -17883
rect 3723 -17893 3733 -17883
rect 3973 -17883 4053 -17873
rect 3973 -17893 3983 -17883
rect 3723 -17943 3983 -17893
rect 4043 -17943 4053 -17883
rect 3653 -17953 4053 -17943
rect 4111 -17533 4511 -17523
rect 4111 -17593 4121 -17533
rect 4181 -17583 4441 -17533
rect 4181 -17593 4191 -17583
rect 4111 -17603 4191 -17593
rect 4431 -17593 4441 -17583
rect 4501 -17593 4511 -17533
rect 4431 -17603 4511 -17593
rect 4111 -17873 4171 -17603
rect 4441 -17613 4511 -17603
rect 4251 -17663 4281 -17643
rect 4231 -17703 4281 -17663
rect 4341 -17663 4371 -17643
rect 4341 -17703 4391 -17663
rect 4231 -17773 4391 -17703
rect 4231 -17813 4281 -17773
rect 4251 -17833 4281 -17813
rect 4341 -17813 4391 -17773
rect 4341 -17833 4371 -17813
rect 4451 -17873 4511 -17613
rect 4111 -17883 4191 -17873
rect 4111 -17943 4121 -17883
rect 4181 -17893 4191 -17883
rect 4431 -17883 4511 -17873
rect 4431 -17893 4441 -17883
rect 4181 -17943 4441 -17893
rect 4501 -17943 4511 -17883
rect 4111 -17953 4511 -17943
rect 4567 -17533 4967 -17523
rect 4567 -17593 4577 -17533
rect 4637 -17583 4897 -17533
rect 4637 -17593 4647 -17583
rect 4567 -17603 4647 -17593
rect 4887 -17593 4897 -17583
rect 4957 -17593 4967 -17533
rect 4887 -17603 4967 -17593
rect 4567 -17873 4627 -17603
rect 4897 -17613 4967 -17603
rect 4707 -17663 4737 -17643
rect 4687 -17703 4737 -17663
rect 4797 -17663 4827 -17643
rect 4797 -17703 4847 -17663
rect 4687 -17773 4847 -17703
rect 4687 -17813 4737 -17773
rect 4707 -17833 4737 -17813
rect 4797 -17813 4847 -17773
rect 4797 -17833 4827 -17813
rect 4907 -17873 4967 -17613
rect 4567 -17883 4647 -17873
rect 4567 -17943 4577 -17883
rect 4637 -17893 4647 -17883
rect 4887 -17883 4967 -17873
rect 4887 -17893 4897 -17883
rect 4637 -17943 4897 -17893
rect 4957 -17943 4967 -17883
rect 4567 -17953 4967 -17943
rect 5023 -17533 5423 -17523
rect 5023 -17593 5033 -17533
rect 5093 -17583 5353 -17533
rect 5093 -17593 5103 -17583
rect 5023 -17603 5103 -17593
rect 5343 -17593 5353 -17583
rect 5413 -17593 5423 -17533
rect 5343 -17603 5423 -17593
rect 5023 -17873 5083 -17603
rect 5353 -17613 5423 -17603
rect 5163 -17663 5193 -17643
rect 5143 -17703 5193 -17663
rect 5253 -17663 5283 -17643
rect 5253 -17703 5303 -17663
rect 5143 -17773 5303 -17703
rect 5143 -17813 5193 -17773
rect 5163 -17833 5193 -17813
rect 5253 -17813 5303 -17773
rect 5253 -17833 5283 -17813
rect 5363 -17873 5423 -17613
rect 5023 -17883 5103 -17873
rect 5023 -17943 5033 -17883
rect 5093 -17893 5103 -17883
rect 5343 -17883 5423 -17873
rect 5343 -17893 5353 -17883
rect 5093 -17943 5353 -17893
rect 5413 -17943 5423 -17883
rect 5023 -17953 5423 -17943
rect 5481 -17533 5881 -17523
rect 5481 -17593 5491 -17533
rect 5551 -17583 5811 -17533
rect 5551 -17593 5561 -17583
rect 5481 -17603 5561 -17593
rect 5801 -17593 5811 -17583
rect 5871 -17593 5881 -17533
rect 5801 -17603 5881 -17593
rect 5481 -17873 5541 -17603
rect 5811 -17613 5881 -17603
rect 5621 -17663 5651 -17643
rect 5601 -17703 5651 -17663
rect 5711 -17663 5741 -17643
rect 5711 -17703 5761 -17663
rect 5601 -17773 5761 -17703
rect 5601 -17813 5651 -17773
rect 5621 -17833 5651 -17813
rect 5711 -17813 5761 -17773
rect 5711 -17833 5741 -17813
rect 5821 -17873 5881 -17613
rect 5481 -17883 5561 -17873
rect 5481 -17943 5491 -17883
rect 5551 -17893 5561 -17883
rect 5801 -17883 5881 -17873
rect 5801 -17893 5811 -17883
rect 5551 -17943 5811 -17893
rect 5871 -17943 5881 -17883
rect 5481 -17953 5881 -17943
rect 5937 -17533 6337 -17523
rect 5937 -17593 5947 -17533
rect 6007 -17583 6267 -17533
rect 6007 -17593 6017 -17583
rect 5937 -17603 6017 -17593
rect 6257 -17593 6267 -17583
rect 6327 -17593 6337 -17533
rect 6257 -17603 6337 -17593
rect 5937 -17873 5997 -17603
rect 6267 -17613 6337 -17603
rect 6077 -17663 6107 -17643
rect 6057 -17703 6107 -17663
rect 6167 -17663 6197 -17643
rect 6167 -17703 6217 -17663
rect 6057 -17773 6217 -17703
rect 6057 -17813 6107 -17773
rect 6077 -17833 6107 -17813
rect 6167 -17813 6217 -17773
rect 6167 -17833 6197 -17813
rect 6277 -17873 6337 -17613
rect 5937 -17883 6017 -17873
rect 5937 -17943 5947 -17883
rect 6007 -17893 6017 -17883
rect 6257 -17883 6337 -17873
rect 6257 -17893 6267 -17883
rect 6007 -17943 6267 -17893
rect 6327 -17943 6337 -17883
rect 5937 -17953 6337 -17943
rect 6393 -17533 6793 -17523
rect 6393 -17593 6403 -17533
rect 6463 -17583 6723 -17533
rect 6463 -17593 6473 -17583
rect 6393 -17603 6473 -17593
rect 6713 -17593 6723 -17583
rect 6783 -17593 6793 -17533
rect 6713 -17603 6793 -17593
rect 6393 -17873 6453 -17603
rect 6723 -17613 6793 -17603
rect 6533 -17663 6563 -17643
rect 6513 -17703 6563 -17663
rect 6623 -17663 6653 -17643
rect 6623 -17703 6673 -17663
rect 6513 -17773 6673 -17703
rect 6513 -17813 6563 -17773
rect 6533 -17833 6563 -17813
rect 6623 -17813 6673 -17773
rect 6623 -17833 6653 -17813
rect 6733 -17873 6793 -17613
rect 6393 -17883 6473 -17873
rect 6393 -17943 6403 -17883
rect 6463 -17893 6473 -17883
rect 6713 -17883 6793 -17873
rect 6713 -17893 6723 -17883
rect 6463 -17943 6723 -17893
rect 6783 -17943 6793 -17883
rect 6393 -17953 6793 -17943
rect 6851 -17533 7251 -17523
rect 6851 -17593 6861 -17533
rect 6921 -17583 7181 -17533
rect 6921 -17593 6931 -17583
rect 6851 -17603 6931 -17593
rect 7171 -17593 7181 -17583
rect 7241 -17593 7251 -17533
rect 7171 -17603 7251 -17593
rect 6851 -17873 6911 -17603
rect 7181 -17613 7251 -17603
rect 6991 -17663 7021 -17643
rect 6971 -17703 7021 -17663
rect 7081 -17663 7111 -17643
rect 7081 -17703 7131 -17663
rect 6971 -17773 7131 -17703
rect 6971 -17813 7021 -17773
rect 6991 -17833 7021 -17813
rect 7081 -17813 7131 -17773
rect 7081 -17833 7111 -17813
rect 7191 -17873 7251 -17613
rect 6851 -17883 6931 -17873
rect 6851 -17943 6861 -17883
rect 6921 -17893 6931 -17883
rect 7171 -17883 7251 -17873
rect 7171 -17893 7181 -17883
rect 6921 -17943 7181 -17893
rect 7241 -17943 7251 -17883
rect 6851 -17953 7251 -17943
rect 7307 -17533 7707 -17523
rect 7307 -17593 7317 -17533
rect 7377 -17583 7637 -17533
rect 7377 -17593 7387 -17583
rect 7307 -17603 7387 -17593
rect 7627 -17593 7637 -17583
rect 7697 -17593 7707 -17533
rect 7627 -17603 7707 -17593
rect 7307 -17873 7367 -17603
rect 7637 -17613 7707 -17603
rect 7447 -17663 7477 -17643
rect 7427 -17703 7477 -17663
rect 7537 -17663 7567 -17643
rect 7537 -17703 7587 -17663
rect 7427 -17773 7587 -17703
rect 7427 -17813 7477 -17773
rect 7447 -17833 7477 -17813
rect 7537 -17813 7587 -17773
rect 7537 -17833 7567 -17813
rect 7647 -17873 7707 -17613
rect 7307 -17883 7387 -17873
rect 7307 -17943 7317 -17883
rect 7377 -17893 7387 -17883
rect 7627 -17883 7707 -17873
rect 7627 -17893 7637 -17883
rect 7377 -17943 7637 -17893
rect 7697 -17943 7707 -17883
rect 7307 -17953 7707 -17943
rect 7763 -17533 8163 -17523
rect 7763 -17593 7773 -17533
rect 7833 -17583 8093 -17533
rect 7833 -17593 7843 -17583
rect 7763 -17603 7843 -17593
rect 8083 -17593 8093 -17583
rect 8153 -17593 8163 -17533
rect 8083 -17603 8163 -17593
rect 7763 -17873 7823 -17603
rect 8093 -17613 8163 -17603
rect 7903 -17663 7933 -17643
rect 7883 -17703 7933 -17663
rect 7993 -17663 8023 -17643
rect 7993 -17703 8043 -17663
rect 7883 -17773 8043 -17703
rect 7883 -17813 7933 -17773
rect 7903 -17833 7933 -17813
rect 7993 -17813 8043 -17773
rect 7993 -17833 8023 -17813
rect 8103 -17873 8163 -17613
rect 7763 -17883 7843 -17873
rect 7763 -17943 7773 -17883
rect 7833 -17893 7843 -17883
rect 8083 -17883 8163 -17873
rect 8083 -17893 8093 -17883
rect 7833 -17943 8093 -17893
rect 8153 -17943 8163 -17883
rect 7763 -17953 8163 -17943
rect 8237 -17533 8637 -17523
rect 8237 -17593 8247 -17533
rect 8307 -17583 8567 -17533
rect 8307 -17593 8317 -17583
rect 8237 -17603 8317 -17593
rect 8557 -17593 8567 -17583
rect 8627 -17593 8637 -17533
rect 8557 -17603 8637 -17593
rect 8237 -17873 8297 -17603
rect 8567 -17613 8637 -17603
rect 8377 -17663 8407 -17643
rect 8357 -17703 8407 -17663
rect 8467 -17663 8497 -17643
rect 8467 -17703 8517 -17663
rect 8357 -17773 8517 -17703
rect 8357 -17813 8407 -17773
rect 8377 -17833 8407 -17813
rect 8467 -17813 8517 -17773
rect 8467 -17833 8497 -17813
rect 8577 -17873 8637 -17613
rect 8237 -17883 8317 -17873
rect 8237 -17943 8247 -17883
rect 8307 -17893 8317 -17883
rect 8557 -17883 8637 -17873
rect 8557 -17893 8567 -17883
rect 8307 -17943 8567 -17893
rect 8627 -17943 8637 -17883
rect 8237 -17953 8637 -17943
rect 8693 -17533 9093 -17523
rect 8693 -17593 8703 -17533
rect 8763 -17583 9023 -17533
rect 8763 -17593 8773 -17583
rect 8693 -17603 8773 -17593
rect 9013 -17593 9023 -17583
rect 9083 -17593 9093 -17533
rect 9013 -17603 9093 -17593
rect 8693 -17873 8753 -17603
rect 9023 -17613 9093 -17603
rect 8833 -17663 8863 -17643
rect 8813 -17703 8863 -17663
rect 8923 -17663 8953 -17643
rect 8923 -17703 8973 -17663
rect 8813 -17773 8973 -17703
rect 8813 -17813 8863 -17773
rect 8833 -17833 8863 -17813
rect 8923 -17813 8973 -17773
rect 8923 -17833 8953 -17813
rect 9033 -17873 9093 -17613
rect 8693 -17883 8773 -17873
rect 8693 -17943 8703 -17883
rect 8763 -17893 8773 -17883
rect 9013 -17883 9093 -17873
rect 9013 -17893 9023 -17883
rect 8763 -17943 9023 -17893
rect 9083 -17943 9093 -17883
rect 8693 -17953 9093 -17943
rect 9151 -17533 9551 -17523
rect 9151 -17593 9161 -17533
rect 9221 -17583 9481 -17533
rect 9221 -17593 9231 -17583
rect 9151 -17603 9231 -17593
rect 9471 -17593 9481 -17583
rect 9541 -17593 9551 -17533
rect 9471 -17603 9551 -17593
rect 9151 -17873 9211 -17603
rect 9481 -17613 9551 -17603
rect 9291 -17663 9321 -17643
rect 9271 -17703 9321 -17663
rect 9381 -17663 9411 -17643
rect 9381 -17703 9431 -17663
rect 9271 -17773 9431 -17703
rect 9271 -17813 9321 -17773
rect 9291 -17833 9321 -17813
rect 9381 -17813 9431 -17773
rect 9381 -17833 9411 -17813
rect 9491 -17873 9551 -17613
rect 9151 -17883 9231 -17873
rect 9151 -17943 9161 -17883
rect 9221 -17893 9231 -17883
rect 9471 -17883 9551 -17873
rect 9471 -17893 9481 -17883
rect 9221 -17943 9481 -17893
rect 9541 -17943 9551 -17883
rect 9151 -17953 9551 -17943
rect 9607 -17533 10007 -17523
rect 9607 -17593 9617 -17533
rect 9677 -17583 9937 -17533
rect 9677 -17593 9687 -17583
rect 9607 -17603 9687 -17593
rect 9927 -17593 9937 -17583
rect 9997 -17593 10007 -17533
rect 9927 -17603 10007 -17593
rect 9607 -17873 9667 -17603
rect 9937 -17613 10007 -17603
rect 9747 -17663 9777 -17643
rect 9727 -17703 9777 -17663
rect 9837 -17663 9867 -17643
rect 9837 -17703 9887 -17663
rect 9727 -17773 9887 -17703
rect 9727 -17813 9777 -17773
rect 9747 -17833 9777 -17813
rect 9837 -17813 9887 -17773
rect 9837 -17833 9867 -17813
rect 9947 -17873 10007 -17613
rect 9607 -17883 9687 -17873
rect 9607 -17943 9617 -17883
rect 9677 -17893 9687 -17883
rect 9927 -17883 10007 -17873
rect 9927 -17893 9937 -17883
rect 9677 -17943 9937 -17893
rect 9997 -17943 10007 -17883
rect 9607 -17953 10007 -17943
rect 10063 -17533 10463 -17523
rect 10063 -17593 10073 -17533
rect 10133 -17583 10393 -17533
rect 10133 -17593 10143 -17583
rect 10063 -17603 10143 -17593
rect 10383 -17593 10393 -17583
rect 10453 -17593 10463 -17533
rect 10383 -17603 10463 -17593
rect 10063 -17873 10123 -17603
rect 10393 -17613 10463 -17603
rect 10203 -17663 10233 -17643
rect 10183 -17703 10233 -17663
rect 10293 -17663 10323 -17643
rect 10293 -17703 10343 -17663
rect 10183 -17773 10343 -17703
rect 10183 -17813 10233 -17773
rect 10203 -17833 10233 -17813
rect 10293 -17813 10343 -17773
rect 10293 -17833 10323 -17813
rect 10403 -17873 10463 -17613
rect 10063 -17883 10143 -17873
rect 10063 -17943 10073 -17883
rect 10133 -17893 10143 -17883
rect 10383 -17883 10463 -17873
rect 10383 -17893 10393 -17883
rect 10133 -17943 10393 -17893
rect 10453 -17943 10463 -17883
rect 10063 -17953 10463 -17943
rect 10521 -17533 10921 -17523
rect 10521 -17593 10531 -17533
rect 10591 -17583 10851 -17533
rect 10591 -17593 10601 -17583
rect 10521 -17603 10601 -17593
rect 10841 -17593 10851 -17583
rect 10911 -17593 10921 -17533
rect 10841 -17603 10921 -17593
rect 10521 -17873 10581 -17603
rect 10851 -17613 10921 -17603
rect 10661 -17663 10691 -17643
rect 10641 -17703 10691 -17663
rect 10751 -17663 10781 -17643
rect 10751 -17703 10801 -17663
rect 10641 -17773 10801 -17703
rect 10641 -17813 10691 -17773
rect 10661 -17833 10691 -17813
rect 10751 -17813 10801 -17773
rect 10751 -17833 10781 -17813
rect 10861 -17873 10921 -17613
rect 10521 -17883 10601 -17873
rect 10521 -17943 10531 -17883
rect 10591 -17893 10601 -17883
rect 10841 -17883 10921 -17873
rect 10841 -17893 10851 -17883
rect 10591 -17943 10851 -17893
rect 10911 -17943 10921 -17883
rect 10521 -17953 10921 -17943
rect 10977 -17533 11377 -17523
rect 10977 -17593 10987 -17533
rect 11047 -17583 11307 -17533
rect 11047 -17593 11057 -17583
rect 10977 -17603 11057 -17593
rect 11297 -17593 11307 -17583
rect 11367 -17593 11377 -17533
rect 11297 -17603 11377 -17593
rect 10977 -17873 11037 -17603
rect 11307 -17613 11377 -17603
rect 11117 -17663 11147 -17643
rect 11097 -17703 11147 -17663
rect 11207 -17663 11237 -17643
rect 11207 -17703 11257 -17663
rect 11097 -17773 11257 -17703
rect 11097 -17813 11147 -17773
rect 11117 -17833 11147 -17813
rect 11207 -17813 11257 -17773
rect 11207 -17833 11237 -17813
rect 11317 -17873 11377 -17613
rect 10977 -17883 11057 -17873
rect 10977 -17943 10987 -17883
rect 11047 -17893 11057 -17883
rect 11297 -17883 11377 -17873
rect 11297 -17893 11307 -17883
rect 11047 -17943 11307 -17893
rect 11367 -17943 11377 -17883
rect 10977 -17953 11377 -17943
rect 11433 -17533 11833 -17523
rect 11433 -17593 11443 -17533
rect 11503 -17583 11763 -17533
rect 11503 -17593 11513 -17583
rect 11433 -17603 11513 -17593
rect 11753 -17593 11763 -17583
rect 11823 -17593 11833 -17533
rect 11753 -17603 11833 -17593
rect 11433 -17873 11493 -17603
rect 11763 -17613 11833 -17603
rect 11573 -17663 11603 -17643
rect 11553 -17703 11603 -17663
rect 11663 -17663 11693 -17643
rect 11663 -17703 11713 -17663
rect 11553 -17773 11713 -17703
rect 11553 -17813 11603 -17773
rect 11573 -17833 11603 -17813
rect 11663 -17813 11713 -17773
rect 11663 -17833 11693 -17813
rect 11773 -17873 11833 -17613
rect 11433 -17883 11513 -17873
rect 11433 -17943 11443 -17883
rect 11503 -17893 11513 -17883
rect 11753 -17883 11833 -17873
rect 11753 -17893 11763 -17883
rect 11503 -17943 11763 -17893
rect 11823 -17943 11833 -17883
rect 11433 -17953 11833 -17943
rect 11891 -17533 12291 -17523
rect 11891 -17593 11901 -17533
rect 11961 -17583 12221 -17533
rect 11961 -17593 11971 -17583
rect 11891 -17603 11971 -17593
rect 12211 -17593 12221 -17583
rect 12281 -17593 12291 -17533
rect 12211 -17603 12291 -17593
rect 11891 -17873 11951 -17603
rect 12221 -17613 12291 -17603
rect 12031 -17663 12061 -17643
rect 12011 -17703 12061 -17663
rect 12121 -17663 12151 -17643
rect 12121 -17703 12171 -17663
rect 12011 -17773 12171 -17703
rect 12011 -17813 12061 -17773
rect 12031 -17833 12061 -17813
rect 12121 -17813 12171 -17773
rect 12121 -17833 12151 -17813
rect 12231 -17873 12291 -17613
rect 11891 -17883 11971 -17873
rect 11891 -17943 11901 -17883
rect 11961 -17893 11971 -17883
rect 12211 -17883 12291 -17873
rect 12211 -17893 12221 -17883
rect 11961 -17943 12221 -17893
rect 12281 -17943 12291 -17883
rect 11891 -17953 12291 -17943
rect 12347 -17533 12747 -17523
rect 12347 -17593 12357 -17533
rect 12417 -17583 12677 -17533
rect 12417 -17593 12427 -17583
rect 12347 -17603 12427 -17593
rect 12667 -17593 12677 -17583
rect 12737 -17593 12747 -17533
rect 12667 -17603 12747 -17593
rect 12347 -17873 12407 -17603
rect 12677 -17613 12747 -17603
rect 12487 -17663 12517 -17643
rect 12467 -17703 12517 -17663
rect 12577 -17663 12607 -17643
rect 12577 -17703 12627 -17663
rect 12467 -17773 12627 -17703
rect 12467 -17813 12517 -17773
rect 12487 -17833 12517 -17813
rect 12577 -17813 12627 -17773
rect 12577 -17833 12607 -17813
rect 12687 -17873 12747 -17613
rect 12347 -17883 12427 -17873
rect 12347 -17943 12357 -17883
rect 12417 -17893 12427 -17883
rect 12667 -17883 12747 -17873
rect 12667 -17893 12677 -17883
rect 12417 -17943 12677 -17893
rect 12737 -17943 12747 -17883
rect 12347 -17953 12747 -17943
rect 12803 -17533 13203 -17523
rect 12803 -17593 12813 -17533
rect 12873 -17583 13133 -17533
rect 12873 -17593 12883 -17583
rect 12803 -17603 12883 -17593
rect 13123 -17593 13133 -17583
rect 13193 -17593 13203 -17533
rect 13123 -17603 13203 -17593
rect 12803 -17873 12863 -17603
rect 13133 -17613 13203 -17603
rect 12943 -17663 12973 -17643
rect 12923 -17703 12973 -17663
rect 13033 -17663 13063 -17643
rect 13033 -17703 13083 -17663
rect 12923 -17773 13083 -17703
rect 12923 -17813 12973 -17773
rect 12943 -17833 12973 -17813
rect 13033 -17813 13083 -17773
rect 13033 -17833 13063 -17813
rect 13143 -17873 13203 -17613
rect 12803 -17883 12883 -17873
rect 12803 -17943 12813 -17883
rect 12873 -17893 12883 -17883
rect 13123 -17883 13203 -17873
rect 13123 -17893 13133 -17883
rect 12873 -17943 13133 -17893
rect 13193 -17943 13203 -17883
rect 12803 -17953 13203 -17943
rect 13261 -17533 13661 -17523
rect 13261 -17593 13271 -17533
rect 13331 -17583 13591 -17533
rect 13331 -17593 13341 -17583
rect 13261 -17603 13341 -17593
rect 13581 -17593 13591 -17583
rect 13651 -17593 13661 -17533
rect 13581 -17603 13661 -17593
rect 13261 -17873 13321 -17603
rect 13591 -17613 13661 -17603
rect 13401 -17663 13431 -17643
rect 13381 -17703 13431 -17663
rect 13491 -17663 13521 -17643
rect 13491 -17703 13541 -17663
rect 13381 -17773 13541 -17703
rect 13381 -17813 13431 -17773
rect 13401 -17833 13431 -17813
rect 13491 -17813 13541 -17773
rect 13491 -17833 13521 -17813
rect 13601 -17873 13661 -17613
rect 13261 -17883 13341 -17873
rect 13261 -17943 13271 -17883
rect 13331 -17893 13341 -17883
rect 13581 -17883 13661 -17873
rect 13581 -17893 13591 -17883
rect 13331 -17943 13591 -17893
rect 13651 -17943 13661 -17883
rect 13261 -17953 13661 -17943
rect 13717 -17533 14117 -17523
rect 13717 -17593 13727 -17533
rect 13787 -17583 14047 -17533
rect 13787 -17593 13797 -17583
rect 13717 -17603 13797 -17593
rect 14037 -17593 14047 -17583
rect 14107 -17593 14117 -17533
rect 14037 -17603 14117 -17593
rect 13717 -17873 13777 -17603
rect 14047 -17613 14117 -17603
rect 13857 -17663 13887 -17643
rect 13837 -17703 13887 -17663
rect 13947 -17663 13977 -17643
rect 13947 -17703 13997 -17663
rect 13837 -17773 13997 -17703
rect 13837 -17813 13887 -17773
rect 13857 -17833 13887 -17813
rect 13947 -17813 13997 -17773
rect 13947 -17833 13977 -17813
rect 14057 -17873 14117 -17613
rect 13717 -17883 13797 -17873
rect 13717 -17943 13727 -17883
rect 13787 -17893 13797 -17883
rect 14037 -17883 14117 -17873
rect 14037 -17893 14047 -17883
rect 13787 -17943 14047 -17893
rect 14107 -17943 14117 -17883
rect 13717 -17953 14117 -17943
rect 14173 -17533 14573 -17523
rect 14173 -17593 14183 -17533
rect 14243 -17583 14503 -17533
rect 14243 -17593 14253 -17583
rect 14173 -17603 14253 -17593
rect 14493 -17593 14503 -17583
rect 14563 -17593 14573 -17533
rect 14493 -17603 14573 -17593
rect 14173 -17873 14233 -17603
rect 14503 -17613 14573 -17603
rect 14313 -17663 14343 -17643
rect 14293 -17703 14343 -17663
rect 14403 -17663 14433 -17643
rect 14403 -17703 14453 -17663
rect 14293 -17773 14453 -17703
rect 14293 -17813 14343 -17773
rect 14313 -17833 14343 -17813
rect 14403 -17813 14453 -17773
rect 14403 -17833 14433 -17813
rect 14513 -17873 14573 -17613
rect 14173 -17883 14253 -17873
rect 14173 -17943 14183 -17883
rect 14243 -17893 14253 -17883
rect 14493 -17883 14573 -17873
rect 14493 -17893 14503 -17883
rect 14243 -17943 14503 -17893
rect 14563 -17943 14573 -17883
rect 14173 -17953 14573 -17943
rect 14631 -17533 15031 -17523
rect 14631 -17593 14641 -17533
rect 14701 -17583 14961 -17533
rect 14701 -17593 14711 -17583
rect 14631 -17603 14711 -17593
rect 14951 -17593 14961 -17583
rect 15021 -17593 15031 -17533
rect 14951 -17603 15031 -17593
rect 14631 -17873 14691 -17603
rect 14961 -17613 15031 -17603
rect 14771 -17663 14801 -17643
rect 14751 -17703 14801 -17663
rect 14861 -17663 14891 -17643
rect 14861 -17703 14911 -17663
rect 14751 -17773 14911 -17703
rect 14751 -17813 14801 -17773
rect 14771 -17833 14801 -17813
rect 14861 -17813 14911 -17773
rect 14861 -17833 14891 -17813
rect 14971 -17873 15031 -17613
rect 14631 -17883 14711 -17873
rect 14631 -17943 14641 -17883
rect 14701 -17893 14711 -17883
rect 14951 -17883 15031 -17873
rect 14951 -17893 14961 -17883
rect 14701 -17943 14961 -17893
rect 15021 -17943 15031 -17883
rect 14631 -17953 15031 -17943
rect 15087 -17533 15487 -17523
rect 15087 -17593 15097 -17533
rect 15157 -17583 15417 -17533
rect 15157 -17593 15167 -17583
rect 15087 -17603 15167 -17593
rect 15407 -17593 15417 -17583
rect 15477 -17593 15487 -17533
rect 15407 -17603 15487 -17593
rect 15087 -17873 15147 -17603
rect 15417 -17613 15487 -17603
rect 15227 -17663 15257 -17643
rect 15207 -17703 15257 -17663
rect 15317 -17663 15347 -17643
rect 15317 -17703 15367 -17663
rect 15207 -17773 15367 -17703
rect 15207 -17813 15257 -17773
rect 15227 -17833 15257 -17813
rect 15317 -17813 15367 -17773
rect 15317 -17833 15347 -17813
rect 15427 -17873 15487 -17613
rect 15087 -17883 15167 -17873
rect 15087 -17943 15097 -17883
rect 15157 -17893 15167 -17883
rect 15407 -17883 15487 -17873
rect 15407 -17893 15417 -17883
rect 15157 -17943 15417 -17893
rect 15477 -17943 15487 -17883
rect 15087 -17953 15487 -17943
rect 1 -18049 401 -18039
rect 1 -18109 11 -18049
rect 71 -18099 331 -18049
rect 71 -18109 81 -18099
rect 1 -18119 81 -18109
rect 321 -18109 331 -18099
rect 391 -18109 401 -18049
rect 321 -18119 401 -18109
rect 1 -18389 61 -18119
rect 331 -18129 401 -18119
rect 141 -18179 171 -18159
rect 121 -18219 171 -18179
rect 231 -18179 261 -18159
rect 231 -18219 281 -18179
rect 121 -18289 281 -18219
rect 121 -18329 171 -18289
rect 141 -18349 171 -18329
rect 231 -18329 281 -18289
rect 231 -18349 261 -18329
rect 341 -18389 401 -18129
rect 1 -18399 81 -18389
rect 1 -18459 11 -18399
rect 71 -18409 81 -18399
rect 321 -18399 401 -18389
rect 321 -18409 331 -18399
rect 71 -18459 331 -18409
rect 391 -18459 401 -18399
rect 1 -18469 401 -18459
rect 457 -18049 857 -18039
rect 457 -18109 467 -18049
rect 527 -18099 787 -18049
rect 527 -18109 537 -18099
rect 457 -18119 537 -18109
rect 777 -18109 787 -18099
rect 847 -18109 857 -18049
rect 777 -18119 857 -18109
rect 457 -18389 517 -18119
rect 787 -18129 857 -18119
rect 597 -18179 627 -18159
rect 577 -18219 627 -18179
rect 687 -18179 717 -18159
rect 687 -18219 737 -18179
rect 577 -18289 737 -18219
rect 577 -18329 627 -18289
rect 597 -18349 627 -18329
rect 687 -18329 737 -18289
rect 687 -18349 717 -18329
rect 797 -18389 857 -18129
rect 457 -18399 537 -18389
rect 457 -18459 467 -18399
rect 527 -18409 537 -18399
rect 777 -18399 857 -18389
rect 777 -18409 787 -18399
rect 527 -18459 787 -18409
rect 847 -18459 857 -18399
rect 457 -18469 857 -18459
rect 913 -18049 1313 -18039
rect 913 -18109 923 -18049
rect 983 -18099 1243 -18049
rect 983 -18109 993 -18099
rect 913 -18119 993 -18109
rect 1233 -18109 1243 -18099
rect 1303 -18109 1313 -18049
rect 1233 -18119 1313 -18109
rect 913 -18389 973 -18119
rect 1243 -18129 1313 -18119
rect 1053 -18179 1083 -18159
rect 1033 -18219 1083 -18179
rect 1143 -18179 1173 -18159
rect 1143 -18219 1193 -18179
rect 1033 -18289 1193 -18219
rect 1033 -18329 1083 -18289
rect 1053 -18349 1083 -18329
rect 1143 -18329 1193 -18289
rect 1143 -18349 1173 -18329
rect 1253 -18389 1313 -18129
rect 913 -18399 993 -18389
rect 913 -18459 923 -18399
rect 983 -18409 993 -18399
rect 1233 -18399 1313 -18389
rect 1233 -18409 1243 -18399
rect 983 -18459 1243 -18409
rect 1303 -18459 1313 -18399
rect 913 -18469 1313 -18459
rect 1371 -18049 1771 -18039
rect 1371 -18109 1381 -18049
rect 1441 -18099 1701 -18049
rect 1441 -18109 1451 -18099
rect 1371 -18119 1451 -18109
rect 1691 -18109 1701 -18099
rect 1761 -18109 1771 -18049
rect 1691 -18119 1771 -18109
rect 1371 -18389 1431 -18119
rect 1701 -18129 1771 -18119
rect 1511 -18179 1541 -18159
rect 1491 -18219 1541 -18179
rect 1601 -18179 1631 -18159
rect 1601 -18219 1651 -18179
rect 1491 -18289 1651 -18219
rect 1491 -18329 1541 -18289
rect 1511 -18349 1541 -18329
rect 1601 -18329 1651 -18289
rect 1601 -18349 1631 -18329
rect 1711 -18389 1771 -18129
rect 1371 -18399 1451 -18389
rect 1371 -18459 1381 -18399
rect 1441 -18409 1451 -18399
rect 1691 -18399 1771 -18389
rect 1691 -18409 1701 -18399
rect 1441 -18459 1701 -18409
rect 1761 -18459 1771 -18399
rect 1371 -18469 1771 -18459
rect 1827 -18049 2227 -18039
rect 1827 -18109 1837 -18049
rect 1897 -18099 2157 -18049
rect 1897 -18109 1907 -18099
rect 1827 -18119 1907 -18109
rect 2147 -18109 2157 -18099
rect 2217 -18109 2227 -18049
rect 2147 -18119 2227 -18109
rect 1827 -18389 1887 -18119
rect 2157 -18129 2227 -18119
rect 1967 -18179 1997 -18159
rect 1947 -18219 1997 -18179
rect 2057 -18179 2087 -18159
rect 2057 -18219 2107 -18179
rect 1947 -18289 2107 -18219
rect 1947 -18329 1997 -18289
rect 1967 -18349 1997 -18329
rect 2057 -18329 2107 -18289
rect 2057 -18349 2087 -18329
rect 2167 -18389 2227 -18129
rect 1827 -18399 1907 -18389
rect 1827 -18459 1837 -18399
rect 1897 -18409 1907 -18399
rect 2147 -18399 2227 -18389
rect 2147 -18409 2157 -18399
rect 1897 -18459 2157 -18409
rect 2217 -18459 2227 -18399
rect 1827 -18469 2227 -18459
rect 2283 -18049 2683 -18039
rect 2283 -18109 2293 -18049
rect 2353 -18099 2613 -18049
rect 2353 -18109 2363 -18099
rect 2283 -18119 2363 -18109
rect 2603 -18109 2613 -18099
rect 2673 -18109 2683 -18049
rect 2603 -18119 2683 -18109
rect 2283 -18389 2343 -18119
rect 2613 -18129 2683 -18119
rect 2423 -18179 2453 -18159
rect 2403 -18219 2453 -18179
rect 2513 -18179 2543 -18159
rect 2513 -18219 2563 -18179
rect 2403 -18289 2563 -18219
rect 2403 -18329 2453 -18289
rect 2423 -18349 2453 -18329
rect 2513 -18329 2563 -18289
rect 2513 -18349 2543 -18329
rect 2623 -18389 2683 -18129
rect 2283 -18399 2363 -18389
rect 2283 -18459 2293 -18399
rect 2353 -18409 2363 -18399
rect 2603 -18399 2683 -18389
rect 2603 -18409 2613 -18399
rect 2353 -18459 2613 -18409
rect 2673 -18459 2683 -18399
rect 2283 -18469 2683 -18459
rect 2741 -18049 3141 -18039
rect 2741 -18109 2751 -18049
rect 2811 -18099 3071 -18049
rect 2811 -18109 2821 -18099
rect 2741 -18119 2821 -18109
rect 3061 -18109 3071 -18099
rect 3131 -18109 3141 -18049
rect 3061 -18119 3141 -18109
rect 2741 -18389 2801 -18119
rect 3071 -18129 3141 -18119
rect 2881 -18179 2911 -18159
rect 2861 -18219 2911 -18179
rect 2971 -18179 3001 -18159
rect 2971 -18219 3021 -18179
rect 2861 -18289 3021 -18219
rect 2861 -18329 2911 -18289
rect 2881 -18349 2911 -18329
rect 2971 -18329 3021 -18289
rect 2971 -18349 3001 -18329
rect 3081 -18389 3141 -18129
rect 2741 -18399 2821 -18389
rect 2741 -18459 2751 -18399
rect 2811 -18409 2821 -18399
rect 3061 -18399 3141 -18389
rect 3061 -18409 3071 -18399
rect 2811 -18459 3071 -18409
rect 3131 -18459 3141 -18399
rect 2741 -18469 3141 -18459
rect 3197 -18049 3597 -18039
rect 3197 -18109 3207 -18049
rect 3267 -18099 3527 -18049
rect 3267 -18109 3277 -18099
rect 3197 -18119 3277 -18109
rect 3517 -18109 3527 -18099
rect 3587 -18109 3597 -18049
rect 3517 -18119 3597 -18109
rect 3197 -18389 3257 -18119
rect 3527 -18129 3597 -18119
rect 3337 -18179 3367 -18159
rect 3317 -18219 3367 -18179
rect 3427 -18179 3457 -18159
rect 3427 -18219 3477 -18179
rect 3317 -18289 3477 -18219
rect 3317 -18329 3367 -18289
rect 3337 -18349 3367 -18329
rect 3427 -18329 3477 -18289
rect 3427 -18349 3457 -18329
rect 3537 -18389 3597 -18129
rect 3197 -18399 3277 -18389
rect 3197 -18459 3207 -18399
rect 3267 -18409 3277 -18399
rect 3517 -18399 3597 -18389
rect 3517 -18409 3527 -18399
rect 3267 -18459 3527 -18409
rect 3587 -18459 3597 -18399
rect 3197 -18469 3597 -18459
rect 3653 -18049 4053 -18039
rect 3653 -18109 3663 -18049
rect 3723 -18099 3983 -18049
rect 3723 -18109 3733 -18099
rect 3653 -18119 3733 -18109
rect 3973 -18109 3983 -18099
rect 4043 -18109 4053 -18049
rect 3973 -18119 4053 -18109
rect 3653 -18389 3713 -18119
rect 3983 -18129 4053 -18119
rect 3793 -18179 3823 -18159
rect 3773 -18219 3823 -18179
rect 3883 -18179 3913 -18159
rect 3883 -18219 3933 -18179
rect 3773 -18289 3933 -18219
rect 3773 -18329 3823 -18289
rect 3793 -18349 3823 -18329
rect 3883 -18329 3933 -18289
rect 3883 -18349 3913 -18329
rect 3993 -18389 4053 -18129
rect 3653 -18399 3733 -18389
rect 3653 -18459 3663 -18399
rect 3723 -18409 3733 -18399
rect 3973 -18399 4053 -18389
rect 3973 -18409 3983 -18399
rect 3723 -18459 3983 -18409
rect 4043 -18459 4053 -18399
rect 3653 -18469 4053 -18459
rect 4111 -18049 4511 -18039
rect 4111 -18109 4121 -18049
rect 4181 -18099 4441 -18049
rect 4181 -18109 4191 -18099
rect 4111 -18119 4191 -18109
rect 4431 -18109 4441 -18099
rect 4501 -18109 4511 -18049
rect 4431 -18119 4511 -18109
rect 4111 -18389 4171 -18119
rect 4441 -18129 4511 -18119
rect 4251 -18179 4281 -18159
rect 4231 -18219 4281 -18179
rect 4341 -18179 4371 -18159
rect 4341 -18219 4391 -18179
rect 4231 -18289 4391 -18219
rect 4231 -18329 4281 -18289
rect 4251 -18349 4281 -18329
rect 4341 -18329 4391 -18289
rect 4341 -18349 4371 -18329
rect 4451 -18389 4511 -18129
rect 4111 -18399 4191 -18389
rect 4111 -18459 4121 -18399
rect 4181 -18409 4191 -18399
rect 4431 -18399 4511 -18389
rect 4431 -18409 4441 -18399
rect 4181 -18459 4441 -18409
rect 4501 -18459 4511 -18399
rect 4111 -18469 4511 -18459
rect 4567 -18049 4967 -18039
rect 4567 -18109 4577 -18049
rect 4637 -18099 4897 -18049
rect 4637 -18109 4647 -18099
rect 4567 -18119 4647 -18109
rect 4887 -18109 4897 -18099
rect 4957 -18109 4967 -18049
rect 4887 -18119 4967 -18109
rect 4567 -18389 4627 -18119
rect 4897 -18129 4967 -18119
rect 4707 -18179 4737 -18159
rect 4687 -18219 4737 -18179
rect 4797 -18179 4827 -18159
rect 4797 -18219 4847 -18179
rect 4687 -18289 4847 -18219
rect 4687 -18329 4737 -18289
rect 4707 -18349 4737 -18329
rect 4797 -18329 4847 -18289
rect 4797 -18349 4827 -18329
rect 4907 -18389 4967 -18129
rect 4567 -18399 4647 -18389
rect 4567 -18459 4577 -18399
rect 4637 -18409 4647 -18399
rect 4887 -18399 4967 -18389
rect 4887 -18409 4897 -18399
rect 4637 -18459 4897 -18409
rect 4957 -18459 4967 -18399
rect 4567 -18469 4967 -18459
rect 5023 -18049 5423 -18039
rect 5023 -18109 5033 -18049
rect 5093 -18099 5353 -18049
rect 5093 -18109 5103 -18099
rect 5023 -18119 5103 -18109
rect 5343 -18109 5353 -18099
rect 5413 -18109 5423 -18049
rect 5343 -18119 5423 -18109
rect 5023 -18389 5083 -18119
rect 5353 -18129 5423 -18119
rect 5163 -18179 5193 -18159
rect 5143 -18219 5193 -18179
rect 5253 -18179 5283 -18159
rect 5253 -18219 5303 -18179
rect 5143 -18289 5303 -18219
rect 5143 -18329 5193 -18289
rect 5163 -18349 5193 -18329
rect 5253 -18329 5303 -18289
rect 5253 -18349 5283 -18329
rect 5363 -18389 5423 -18129
rect 5023 -18399 5103 -18389
rect 5023 -18459 5033 -18399
rect 5093 -18409 5103 -18399
rect 5343 -18399 5423 -18389
rect 5343 -18409 5353 -18399
rect 5093 -18459 5353 -18409
rect 5413 -18459 5423 -18399
rect 5023 -18469 5423 -18459
rect 5481 -18049 5881 -18039
rect 5481 -18109 5491 -18049
rect 5551 -18099 5811 -18049
rect 5551 -18109 5561 -18099
rect 5481 -18119 5561 -18109
rect 5801 -18109 5811 -18099
rect 5871 -18109 5881 -18049
rect 5801 -18119 5881 -18109
rect 5481 -18389 5541 -18119
rect 5811 -18129 5881 -18119
rect 5621 -18179 5651 -18159
rect 5601 -18219 5651 -18179
rect 5711 -18179 5741 -18159
rect 5711 -18219 5761 -18179
rect 5601 -18289 5761 -18219
rect 5601 -18329 5651 -18289
rect 5621 -18349 5651 -18329
rect 5711 -18329 5761 -18289
rect 5711 -18349 5741 -18329
rect 5821 -18389 5881 -18129
rect 5481 -18399 5561 -18389
rect 5481 -18459 5491 -18399
rect 5551 -18409 5561 -18399
rect 5801 -18399 5881 -18389
rect 5801 -18409 5811 -18399
rect 5551 -18459 5811 -18409
rect 5871 -18459 5881 -18399
rect 5481 -18469 5881 -18459
rect 5937 -18049 6337 -18039
rect 5937 -18109 5947 -18049
rect 6007 -18099 6267 -18049
rect 6007 -18109 6017 -18099
rect 5937 -18119 6017 -18109
rect 6257 -18109 6267 -18099
rect 6327 -18109 6337 -18049
rect 6257 -18119 6337 -18109
rect 5937 -18389 5997 -18119
rect 6267 -18129 6337 -18119
rect 6077 -18179 6107 -18159
rect 6057 -18219 6107 -18179
rect 6167 -18179 6197 -18159
rect 6167 -18219 6217 -18179
rect 6057 -18289 6217 -18219
rect 6057 -18329 6107 -18289
rect 6077 -18349 6107 -18329
rect 6167 -18329 6217 -18289
rect 6167 -18349 6197 -18329
rect 6277 -18389 6337 -18129
rect 5937 -18399 6017 -18389
rect 5937 -18459 5947 -18399
rect 6007 -18409 6017 -18399
rect 6257 -18399 6337 -18389
rect 6257 -18409 6267 -18399
rect 6007 -18459 6267 -18409
rect 6327 -18459 6337 -18399
rect 5937 -18469 6337 -18459
rect 6393 -18049 6793 -18039
rect 6393 -18109 6403 -18049
rect 6463 -18099 6723 -18049
rect 6463 -18109 6473 -18099
rect 6393 -18119 6473 -18109
rect 6713 -18109 6723 -18099
rect 6783 -18109 6793 -18049
rect 6713 -18119 6793 -18109
rect 6393 -18389 6453 -18119
rect 6723 -18129 6793 -18119
rect 6533 -18179 6563 -18159
rect 6513 -18219 6563 -18179
rect 6623 -18179 6653 -18159
rect 6623 -18219 6673 -18179
rect 6513 -18289 6673 -18219
rect 6513 -18329 6563 -18289
rect 6533 -18349 6563 -18329
rect 6623 -18329 6673 -18289
rect 6623 -18349 6653 -18329
rect 6733 -18389 6793 -18129
rect 6393 -18399 6473 -18389
rect 6393 -18459 6403 -18399
rect 6463 -18409 6473 -18399
rect 6713 -18399 6793 -18389
rect 6713 -18409 6723 -18399
rect 6463 -18459 6723 -18409
rect 6783 -18459 6793 -18399
rect 6393 -18469 6793 -18459
rect 6851 -18049 7251 -18039
rect 6851 -18109 6861 -18049
rect 6921 -18099 7181 -18049
rect 6921 -18109 6931 -18099
rect 6851 -18119 6931 -18109
rect 7171 -18109 7181 -18099
rect 7241 -18109 7251 -18049
rect 7171 -18119 7251 -18109
rect 6851 -18389 6911 -18119
rect 7181 -18129 7251 -18119
rect 6991 -18179 7021 -18159
rect 6971 -18219 7021 -18179
rect 7081 -18179 7111 -18159
rect 7081 -18219 7131 -18179
rect 6971 -18289 7131 -18219
rect 6971 -18329 7021 -18289
rect 6991 -18349 7021 -18329
rect 7081 -18329 7131 -18289
rect 7081 -18349 7111 -18329
rect 7191 -18389 7251 -18129
rect 6851 -18399 6931 -18389
rect 6851 -18459 6861 -18399
rect 6921 -18409 6931 -18399
rect 7171 -18399 7251 -18389
rect 7171 -18409 7181 -18399
rect 6921 -18459 7181 -18409
rect 7241 -18459 7251 -18399
rect 6851 -18469 7251 -18459
rect 7307 -18049 7707 -18039
rect 7307 -18109 7317 -18049
rect 7377 -18099 7637 -18049
rect 7377 -18109 7387 -18099
rect 7307 -18119 7387 -18109
rect 7627 -18109 7637 -18099
rect 7697 -18109 7707 -18049
rect 7627 -18119 7707 -18109
rect 7307 -18389 7367 -18119
rect 7637 -18129 7707 -18119
rect 7447 -18179 7477 -18159
rect 7427 -18219 7477 -18179
rect 7537 -18179 7567 -18159
rect 7537 -18219 7587 -18179
rect 7427 -18289 7587 -18219
rect 7427 -18329 7477 -18289
rect 7447 -18349 7477 -18329
rect 7537 -18329 7587 -18289
rect 7537 -18349 7567 -18329
rect 7647 -18389 7707 -18129
rect 7307 -18399 7387 -18389
rect 7307 -18459 7317 -18399
rect 7377 -18409 7387 -18399
rect 7627 -18399 7707 -18389
rect 7627 -18409 7637 -18399
rect 7377 -18459 7637 -18409
rect 7697 -18459 7707 -18399
rect 7307 -18469 7707 -18459
rect 7763 -18049 8163 -18039
rect 7763 -18109 7773 -18049
rect 7833 -18099 8093 -18049
rect 7833 -18109 7843 -18099
rect 7763 -18119 7843 -18109
rect 8083 -18109 8093 -18099
rect 8153 -18109 8163 -18049
rect 8083 -18119 8163 -18109
rect 7763 -18389 7823 -18119
rect 8093 -18129 8163 -18119
rect 7903 -18179 7933 -18159
rect 7883 -18219 7933 -18179
rect 7993 -18179 8023 -18159
rect 7993 -18219 8043 -18179
rect 7883 -18289 8043 -18219
rect 7883 -18329 7933 -18289
rect 7903 -18349 7933 -18329
rect 7993 -18329 8043 -18289
rect 7993 -18349 8023 -18329
rect 8103 -18389 8163 -18129
rect 7763 -18399 7843 -18389
rect 7763 -18459 7773 -18399
rect 7833 -18409 7843 -18399
rect 8083 -18399 8163 -18389
rect 8083 -18409 8093 -18399
rect 7833 -18459 8093 -18409
rect 8153 -18459 8163 -18399
rect 7763 -18469 8163 -18459
rect 8237 -18049 8637 -18039
rect 8237 -18109 8247 -18049
rect 8307 -18099 8567 -18049
rect 8307 -18109 8317 -18099
rect 8237 -18119 8317 -18109
rect 8557 -18109 8567 -18099
rect 8627 -18109 8637 -18049
rect 8557 -18119 8637 -18109
rect 8237 -18389 8297 -18119
rect 8567 -18129 8637 -18119
rect 8377 -18179 8407 -18159
rect 8357 -18219 8407 -18179
rect 8467 -18179 8497 -18159
rect 8467 -18219 8517 -18179
rect 8357 -18289 8517 -18219
rect 8357 -18329 8407 -18289
rect 8377 -18349 8407 -18329
rect 8467 -18329 8517 -18289
rect 8467 -18349 8497 -18329
rect 8577 -18389 8637 -18129
rect 8237 -18399 8317 -18389
rect 8237 -18459 8247 -18399
rect 8307 -18409 8317 -18399
rect 8557 -18399 8637 -18389
rect 8557 -18409 8567 -18399
rect 8307 -18459 8567 -18409
rect 8627 -18459 8637 -18399
rect 8237 -18469 8637 -18459
rect 8693 -18049 9093 -18039
rect 8693 -18109 8703 -18049
rect 8763 -18099 9023 -18049
rect 8763 -18109 8773 -18099
rect 8693 -18119 8773 -18109
rect 9013 -18109 9023 -18099
rect 9083 -18109 9093 -18049
rect 9013 -18119 9093 -18109
rect 8693 -18389 8753 -18119
rect 9023 -18129 9093 -18119
rect 8833 -18179 8863 -18159
rect 8813 -18219 8863 -18179
rect 8923 -18179 8953 -18159
rect 8923 -18219 8973 -18179
rect 8813 -18289 8973 -18219
rect 8813 -18329 8863 -18289
rect 8833 -18349 8863 -18329
rect 8923 -18329 8973 -18289
rect 8923 -18349 8953 -18329
rect 9033 -18389 9093 -18129
rect 8693 -18399 8773 -18389
rect 8693 -18459 8703 -18399
rect 8763 -18409 8773 -18399
rect 9013 -18399 9093 -18389
rect 9013 -18409 9023 -18399
rect 8763 -18459 9023 -18409
rect 9083 -18459 9093 -18399
rect 8693 -18469 9093 -18459
rect 9151 -18049 9551 -18039
rect 9151 -18109 9161 -18049
rect 9221 -18099 9481 -18049
rect 9221 -18109 9231 -18099
rect 9151 -18119 9231 -18109
rect 9471 -18109 9481 -18099
rect 9541 -18109 9551 -18049
rect 9471 -18119 9551 -18109
rect 9151 -18389 9211 -18119
rect 9481 -18129 9551 -18119
rect 9291 -18179 9321 -18159
rect 9271 -18219 9321 -18179
rect 9381 -18179 9411 -18159
rect 9381 -18219 9431 -18179
rect 9271 -18289 9431 -18219
rect 9271 -18329 9321 -18289
rect 9291 -18349 9321 -18329
rect 9381 -18329 9431 -18289
rect 9381 -18349 9411 -18329
rect 9491 -18389 9551 -18129
rect 9151 -18399 9231 -18389
rect 9151 -18459 9161 -18399
rect 9221 -18409 9231 -18399
rect 9471 -18399 9551 -18389
rect 9471 -18409 9481 -18399
rect 9221 -18459 9481 -18409
rect 9541 -18459 9551 -18399
rect 9151 -18469 9551 -18459
rect 9607 -18049 10007 -18039
rect 9607 -18109 9617 -18049
rect 9677 -18099 9937 -18049
rect 9677 -18109 9687 -18099
rect 9607 -18119 9687 -18109
rect 9927 -18109 9937 -18099
rect 9997 -18109 10007 -18049
rect 9927 -18119 10007 -18109
rect 9607 -18389 9667 -18119
rect 9937 -18129 10007 -18119
rect 9747 -18179 9777 -18159
rect 9727 -18219 9777 -18179
rect 9837 -18179 9867 -18159
rect 9837 -18219 9887 -18179
rect 9727 -18289 9887 -18219
rect 9727 -18329 9777 -18289
rect 9747 -18349 9777 -18329
rect 9837 -18329 9887 -18289
rect 9837 -18349 9867 -18329
rect 9947 -18389 10007 -18129
rect 9607 -18399 9687 -18389
rect 9607 -18459 9617 -18399
rect 9677 -18409 9687 -18399
rect 9927 -18399 10007 -18389
rect 9927 -18409 9937 -18399
rect 9677 -18459 9937 -18409
rect 9997 -18459 10007 -18399
rect 9607 -18469 10007 -18459
rect 10063 -18049 10463 -18039
rect 10063 -18109 10073 -18049
rect 10133 -18099 10393 -18049
rect 10133 -18109 10143 -18099
rect 10063 -18119 10143 -18109
rect 10383 -18109 10393 -18099
rect 10453 -18109 10463 -18049
rect 10383 -18119 10463 -18109
rect 10063 -18389 10123 -18119
rect 10393 -18129 10463 -18119
rect 10203 -18179 10233 -18159
rect 10183 -18219 10233 -18179
rect 10293 -18179 10323 -18159
rect 10293 -18219 10343 -18179
rect 10183 -18289 10343 -18219
rect 10183 -18329 10233 -18289
rect 10203 -18349 10233 -18329
rect 10293 -18329 10343 -18289
rect 10293 -18349 10323 -18329
rect 10403 -18389 10463 -18129
rect 10063 -18399 10143 -18389
rect 10063 -18459 10073 -18399
rect 10133 -18409 10143 -18399
rect 10383 -18399 10463 -18389
rect 10383 -18409 10393 -18399
rect 10133 -18459 10393 -18409
rect 10453 -18459 10463 -18399
rect 10063 -18469 10463 -18459
rect 10521 -18049 10921 -18039
rect 10521 -18109 10531 -18049
rect 10591 -18099 10851 -18049
rect 10591 -18109 10601 -18099
rect 10521 -18119 10601 -18109
rect 10841 -18109 10851 -18099
rect 10911 -18109 10921 -18049
rect 10841 -18119 10921 -18109
rect 10521 -18389 10581 -18119
rect 10851 -18129 10921 -18119
rect 10661 -18179 10691 -18159
rect 10641 -18219 10691 -18179
rect 10751 -18179 10781 -18159
rect 10751 -18219 10801 -18179
rect 10641 -18289 10801 -18219
rect 10641 -18329 10691 -18289
rect 10661 -18349 10691 -18329
rect 10751 -18329 10801 -18289
rect 10751 -18349 10781 -18329
rect 10861 -18389 10921 -18129
rect 10521 -18399 10601 -18389
rect 10521 -18459 10531 -18399
rect 10591 -18409 10601 -18399
rect 10841 -18399 10921 -18389
rect 10841 -18409 10851 -18399
rect 10591 -18459 10851 -18409
rect 10911 -18459 10921 -18399
rect 10521 -18469 10921 -18459
rect 10977 -18049 11377 -18039
rect 10977 -18109 10987 -18049
rect 11047 -18099 11307 -18049
rect 11047 -18109 11057 -18099
rect 10977 -18119 11057 -18109
rect 11297 -18109 11307 -18099
rect 11367 -18109 11377 -18049
rect 11297 -18119 11377 -18109
rect 10977 -18389 11037 -18119
rect 11307 -18129 11377 -18119
rect 11117 -18179 11147 -18159
rect 11097 -18219 11147 -18179
rect 11207 -18179 11237 -18159
rect 11207 -18219 11257 -18179
rect 11097 -18289 11257 -18219
rect 11097 -18329 11147 -18289
rect 11117 -18349 11147 -18329
rect 11207 -18329 11257 -18289
rect 11207 -18349 11237 -18329
rect 11317 -18389 11377 -18129
rect 10977 -18399 11057 -18389
rect 10977 -18459 10987 -18399
rect 11047 -18409 11057 -18399
rect 11297 -18399 11377 -18389
rect 11297 -18409 11307 -18399
rect 11047 -18459 11307 -18409
rect 11367 -18459 11377 -18399
rect 10977 -18469 11377 -18459
rect 11433 -18049 11833 -18039
rect 11433 -18109 11443 -18049
rect 11503 -18099 11763 -18049
rect 11503 -18109 11513 -18099
rect 11433 -18119 11513 -18109
rect 11753 -18109 11763 -18099
rect 11823 -18109 11833 -18049
rect 11753 -18119 11833 -18109
rect 11433 -18389 11493 -18119
rect 11763 -18129 11833 -18119
rect 11573 -18179 11603 -18159
rect 11553 -18219 11603 -18179
rect 11663 -18179 11693 -18159
rect 11663 -18219 11713 -18179
rect 11553 -18289 11713 -18219
rect 11553 -18329 11603 -18289
rect 11573 -18349 11603 -18329
rect 11663 -18329 11713 -18289
rect 11663 -18349 11693 -18329
rect 11773 -18389 11833 -18129
rect 11433 -18399 11513 -18389
rect 11433 -18459 11443 -18399
rect 11503 -18409 11513 -18399
rect 11753 -18399 11833 -18389
rect 11753 -18409 11763 -18399
rect 11503 -18459 11763 -18409
rect 11823 -18459 11833 -18399
rect 11433 -18469 11833 -18459
rect 11891 -18049 12291 -18039
rect 11891 -18109 11901 -18049
rect 11961 -18099 12221 -18049
rect 11961 -18109 11971 -18099
rect 11891 -18119 11971 -18109
rect 12211 -18109 12221 -18099
rect 12281 -18109 12291 -18049
rect 12211 -18119 12291 -18109
rect 11891 -18389 11951 -18119
rect 12221 -18129 12291 -18119
rect 12031 -18179 12061 -18159
rect 12011 -18219 12061 -18179
rect 12121 -18179 12151 -18159
rect 12121 -18219 12171 -18179
rect 12011 -18289 12171 -18219
rect 12011 -18329 12061 -18289
rect 12031 -18349 12061 -18329
rect 12121 -18329 12171 -18289
rect 12121 -18349 12151 -18329
rect 12231 -18389 12291 -18129
rect 11891 -18399 11971 -18389
rect 11891 -18459 11901 -18399
rect 11961 -18409 11971 -18399
rect 12211 -18399 12291 -18389
rect 12211 -18409 12221 -18399
rect 11961 -18459 12221 -18409
rect 12281 -18459 12291 -18399
rect 11891 -18469 12291 -18459
rect 12347 -18049 12747 -18039
rect 12347 -18109 12357 -18049
rect 12417 -18099 12677 -18049
rect 12417 -18109 12427 -18099
rect 12347 -18119 12427 -18109
rect 12667 -18109 12677 -18099
rect 12737 -18109 12747 -18049
rect 12667 -18119 12747 -18109
rect 12347 -18389 12407 -18119
rect 12677 -18129 12747 -18119
rect 12487 -18179 12517 -18159
rect 12467 -18219 12517 -18179
rect 12577 -18179 12607 -18159
rect 12577 -18219 12627 -18179
rect 12467 -18289 12627 -18219
rect 12467 -18329 12517 -18289
rect 12487 -18349 12517 -18329
rect 12577 -18329 12627 -18289
rect 12577 -18349 12607 -18329
rect 12687 -18389 12747 -18129
rect 12347 -18399 12427 -18389
rect 12347 -18459 12357 -18399
rect 12417 -18409 12427 -18399
rect 12667 -18399 12747 -18389
rect 12667 -18409 12677 -18399
rect 12417 -18459 12677 -18409
rect 12737 -18459 12747 -18399
rect 12347 -18469 12747 -18459
rect 12803 -18049 13203 -18039
rect 12803 -18109 12813 -18049
rect 12873 -18099 13133 -18049
rect 12873 -18109 12883 -18099
rect 12803 -18119 12883 -18109
rect 13123 -18109 13133 -18099
rect 13193 -18109 13203 -18049
rect 13123 -18119 13203 -18109
rect 12803 -18389 12863 -18119
rect 13133 -18129 13203 -18119
rect 12943 -18179 12973 -18159
rect 12923 -18219 12973 -18179
rect 13033 -18179 13063 -18159
rect 13033 -18219 13083 -18179
rect 12923 -18289 13083 -18219
rect 12923 -18329 12973 -18289
rect 12943 -18349 12973 -18329
rect 13033 -18329 13083 -18289
rect 13033 -18349 13063 -18329
rect 13143 -18389 13203 -18129
rect 12803 -18399 12883 -18389
rect 12803 -18459 12813 -18399
rect 12873 -18409 12883 -18399
rect 13123 -18399 13203 -18389
rect 13123 -18409 13133 -18399
rect 12873 -18459 13133 -18409
rect 13193 -18459 13203 -18399
rect 12803 -18469 13203 -18459
rect 13261 -18049 13661 -18039
rect 13261 -18109 13271 -18049
rect 13331 -18099 13591 -18049
rect 13331 -18109 13341 -18099
rect 13261 -18119 13341 -18109
rect 13581 -18109 13591 -18099
rect 13651 -18109 13661 -18049
rect 13581 -18119 13661 -18109
rect 13261 -18389 13321 -18119
rect 13591 -18129 13661 -18119
rect 13401 -18179 13431 -18159
rect 13381 -18219 13431 -18179
rect 13491 -18179 13521 -18159
rect 13491 -18219 13541 -18179
rect 13381 -18289 13541 -18219
rect 13381 -18329 13431 -18289
rect 13401 -18349 13431 -18329
rect 13491 -18329 13541 -18289
rect 13491 -18349 13521 -18329
rect 13601 -18389 13661 -18129
rect 13261 -18399 13341 -18389
rect 13261 -18459 13271 -18399
rect 13331 -18409 13341 -18399
rect 13581 -18399 13661 -18389
rect 13581 -18409 13591 -18399
rect 13331 -18459 13591 -18409
rect 13651 -18459 13661 -18399
rect 13261 -18469 13661 -18459
rect 13717 -18049 14117 -18039
rect 13717 -18109 13727 -18049
rect 13787 -18099 14047 -18049
rect 13787 -18109 13797 -18099
rect 13717 -18119 13797 -18109
rect 14037 -18109 14047 -18099
rect 14107 -18109 14117 -18049
rect 14037 -18119 14117 -18109
rect 13717 -18389 13777 -18119
rect 14047 -18129 14117 -18119
rect 13857 -18179 13887 -18159
rect 13837 -18219 13887 -18179
rect 13947 -18179 13977 -18159
rect 13947 -18219 13997 -18179
rect 13837 -18289 13997 -18219
rect 13837 -18329 13887 -18289
rect 13857 -18349 13887 -18329
rect 13947 -18329 13997 -18289
rect 13947 -18349 13977 -18329
rect 14057 -18389 14117 -18129
rect 13717 -18399 13797 -18389
rect 13717 -18459 13727 -18399
rect 13787 -18409 13797 -18399
rect 14037 -18399 14117 -18389
rect 14037 -18409 14047 -18399
rect 13787 -18459 14047 -18409
rect 14107 -18459 14117 -18399
rect 13717 -18469 14117 -18459
rect 14173 -18049 14573 -18039
rect 14173 -18109 14183 -18049
rect 14243 -18099 14503 -18049
rect 14243 -18109 14253 -18099
rect 14173 -18119 14253 -18109
rect 14493 -18109 14503 -18099
rect 14563 -18109 14573 -18049
rect 14493 -18119 14573 -18109
rect 14173 -18389 14233 -18119
rect 14503 -18129 14573 -18119
rect 14313 -18179 14343 -18159
rect 14293 -18219 14343 -18179
rect 14403 -18179 14433 -18159
rect 14403 -18219 14453 -18179
rect 14293 -18289 14453 -18219
rect 14293 -18329 14343 -18289
rect 14313 -18349 14343 -18329
rect 14403 -18329 14453 -18289
rect 14403 -18349 14433 -18329
rect 14513 -18389 14573 -18129
rect 14173 -18399 14253 -18389
rect 14173 -18459 14183 -18399
rect 14243 -18409 14253 -18399
rect 14493 -18399 14573 -18389
rect 14493 -18409 14503 -18399
rect 14243 -18459 14503 -18409
rect 14563 -18459 14573 -18399
rect 14173 -18469 14573 -18459
rect 14631 -18049 15031 -18039
rect 14631 -18109 14641 -18049
rect 14701 -18099 14961 -18049
rect 14701 -18109 14711 -18099
rect 14631 -18119 14711 -18109
rect 14951 -18109 14961 -18099
rect 15021 -18109 15031 -18049
rect 14951 -18119 15031 -18109
rect 14631 -18389 14691 -18119
rect 14961 -18129 15031 -18119
rect 14771 -18179 14801 -18159
rect 14751 -18219 14801 -18179
rect 14861 -18179 14891 -18159
rect 14861 -18219 14911 -18179
rect 14751 -18289 14911 -18219
rect 14751 -18329 14801 -18289
rect 14771 -18349 14801 -18329
rect 14861 -18329 14911 -18289
rect 14861 -18349 14891 -18329
rect 14971 -18389 15031 -18129
rect 14631 -18399 14711 -18389
rect 14631 -18459 14641 -18399
rect 14701 -18409 14711 -18399
rect 14951 -18399 15031 -18389
rect 14951 -18409 14961 -18399
rect 14701 -18459 14961 -18409
rect 15021 -18459 15031 -18399
rect 14631 -18469 15031 -18459
rect 15087 -18049 15487 -18039
rect 15087 -18109 15097 -18049
rect 15157 -18099 15417 -18049
rect 15157 -18109 15167 -18099
rect 15087 -18119 15167 -18109
rect 15407 -18109 15417 -18099
rect 15477 -18109 15487 -18049
rect 15407 -18119 15487 -18109
rect 15087 -18389 15147 -18119
rect 15417 -18129 15487 -18119
rect 15227 -18179 15257 -18159
rect 15207 -18219 15257 -18179
rect 15317 -18179 15347 -18159
rect 15317 -18219 15367 -18179
rect 15207 -18289 15367 -18219
rect 15207 -18329 15257 -18289
rect 15227 -18349 15257 -18329
rect 15317 -18329 15367 -18289
rect 15317 -18349 15347 -18329
rect 15427 -18389 15487 -18129
rect 15087 -18399 15167 -18389
rect 15087 -18459 15097 -18399
rect 15157 -18409 15167 -18399
rect 15407 -18399 15487 -18389
rect 15407 -18409 15417 -18399
rect 15157 -18459 15417 -18409
rect 15477 -18459 15487 -18399
rect 15087 -18469 15487 -18459
rect 1 -18551 401 -18541
rect 1 -18611 11 -18551
rect 71 -18601 331 -18551
rect 71 -18611 81 -18601
rect 1 -18621 81 -18611
rect 321 -18611 331 -18601
rect 391 -18611 401 -18551
rect 321 -18621 401 -18611
rect 1 -18891 61 -18621
rect 331 -18631 401 -18621
rect 141 -18681 171 -18661
rect 121 -18721 171 -18681
rect 231 -18681 261 -18661
rect 231 -18721 281 -18681
rect 121 -18791 281 -18721
rect 121 -18831 171 -18791
rect 141 -18851 171 -18831
rect 231 -18831 281 -18791
rect 231 -18851 261 -18831
rect 341 -18891 401 -18631
rect 1 -18901 81 -18891
rect 1 -18961 11 -18901
rect 71 -18911 81 -18901
rect 321 -18901 401 -18891
rect 321 -18911 331 -18901
rect 71 -18961 331 -18911
rect 391 -18961 401 -18901
rect 1 -18971 401 -18961
rect 457 -18551 857 -18541
rect 457 -18611 467 -18551
rect 527 -18601 787 -18551
rect 527 -18611 537 -18601
rect 457 -18621 537 -18611
rect 777 -18611 787 -18601
rect 847 -18611 857 -18551
rect 777 -18621 857 -18611
rect 457 -18891 517 -18621
rect 787 -18631 857 -18621
rect 597 -18681 627 -18661
rect 577 -18721 627 -18681
rect 687 -18681 717 -18661
rect 687 -18721 737 -18681
rect 577 -18791 737 -18721
rect 577 -18831 627 -18791
rect 597 -18851 627 -18831
rect 687 -18831 737 -18791
rect 687 -18851 717 -18831
rect 797 -18891 857 -18631
rect 457 -18901 537 -18891
rect 457 -18961 467 -18901
rect 527 -18911 537 -18901
rect 777 -18901 857 -18891
rect 777 -18911 787 -18901
rect 527 -18961 787 -18911
rect 847 -18961 857 -18901
rect 457 -18971 857 -18961
rect 913 -18551 1313 -18541
rect 913 -18611 923 -18551
rect 983 -18601 1243 -18551
rect 983 -18611 993 -18601
rect 913 -18621 993 -18611
rect 1233 -18611 1243 -18601
rect 1303 -18611 1313 -18551
rect 1233 -18621 1313 -18611
rect 913 -18891 973 -18621
rect 1243 -18631 1313 -18621
rect 1053 -18681 1083 -18661
rect 1033 -18721 1083 -18681
rect 1143 -18681 1173 -18661
rect 1143 -18721 1193 -18681
rect 1033 -18791 1193 -18721
rect 1033 -18831 1083 -18791
rect 1053 -18851 1083 -18831
rect 1143 -18831 1193 -18791
rect 1143 -18851 1173 -18831
rect 1253 -18891 1313 -18631
rect 913 -18901 993 -18891
rect 913 -18961 923 -18901
rect 983 -18911 993 -18901
rect 1233 -18901 1313 -18891
rect 1233 -18911 1243 -18901
rect 983 -18961 1243 -18911
rect 1303 -18961 1313 -18901
rect 913 -18971 1313 -18961
rect 1371 -18551 1771 -18541
rect 1371 -18611 1381 -18551
rect 1441 -18601 1701 -18551
rect 1441 -18611 1451 -18601
rect 1371 -18621 1451 -18611
rect 1691 -18611 1701 -18601
rect 1761 -18611 1771 -18551
rect 1691 -18621 1771 -18611
rect 1371 -18891 1431 -18621
rect 1701 -18631 1771 -18621
rect 1511 -18681 1541 -18661
rect 1491 -18721 1541 -18681
rect 1601 -18681 1631 -18661
rect 1601 -18721 1651 -18681
rect 1491 -18791 1651 -18721
rect 1491 -18831 1541 -18791
rect 1511 -18851 1541 -18831
rect 1601 -18831 1651 -18791
rect 1601 -18851 1631 -18831
rect 1711 -18891 1771 -18631
rect 1371 -18901 1451 -18891
rect 1371 -18961 1381 -18901
rect 1441 -18911 1451 -18901
rect 1691 -18901 1771 -18891
rect 1691 -18911 1701 -18901
rect 1441 -18961 1701 -18911
rect 1761 -18961 1771 -18901
rect 1371 -18971 1771 -18961
rect 1827 -18551 2227 -18541
rect 1827 -18611 1837 -18551
rect 1897 -18601 2157 -18551
rect 1897 -18611 1907 -18601
rect 1827 -18621 1907 -18611
rect 2147 -18611 2157 -18601
rect 2217 -18611 2227 -18551
rect 2147 -18621 2227 -18611
rect 1827 -18891 1887 -18621
rect 2157 -18631 2227 -18621
rect 1967 -18681 1997 -18661
rect 1947 -18721 1997 -18681
rect 2057 -18681 2087 -18661
rect 2057 -18721 2107 -18681
rect 1947 -18791 2107 -18721
rect 1947 -18831 1997 -18791
rect 1967 -18851 1997 -18831
rect 2057 -18831 2107 -18791
rect 2057 -18851 2087 -18831
rect 2167 -18891 2227 -18631
rect 1827 -18901 1907 -18891
rect 1827 -18961 1837 -18901
rect 1897 -18911 1907 -18901
rect 2147 -18901 2227 -18891
rect 2147 -18911 2157 -18901
rect 1897 -18961 2157 -18911
rect 2217 -18961 2227 -18901
rect 1827 -18971 2227 -18961
rect 2283 -18551 2683 -18541
rect 2283 -18611 2293 -18551
rect 2353 -18601 2613 -18551
rect 2353 -18611 2363 -18601
rect 2283 -18621 2363 -18611
rect 2603 -18611 2613 -18601
rect 2673 -18611 2683 -18551
rect 2603 -18621 2683 -18611
rect 2283 -18891 2343 -18621
rect 2613 -18631 2683 -18621
rect 2423 -18681 2453 -18661
rect 2403 -18721 2453 -18681
rect 2513 -18681 2543 -18661
rect 2513 -18721 2563 -18681
rect 2403 -18791 2563 -18721
rect 2403 -18831 2453 -18791
rect 2423 -18851 2453 -18831
rect 2513 -18831 2563 -18791
rect 2513 -18851 2543 -18831
rect 2623 -18891 2683 -18631
rect 2283 -18901 2363 -18891
rect 2283 -18961 2293 -18901
rect 2353 -18911 2363 -18901
rect 2603 -18901 2683 -18891
rect 2603 -18911 2613 -18901
rect 2353 -18961 2613 -18911
rect 2673 -18961 2683 -18901
rect 2283 -18971 2683 -18961
rect 2741 -18551 3141 -18541
rect 2741 -18611 2751 -18551
rect 2811 -18601 3071 -18551
rect 2811 -18611 2821 -18601
rect 2741 -18621 2821 -18611
rect 3061 -18611 3071 -18601
rect 3131 -18611 3141 -18551
rect 3061 -18621 3141 -18611
rect 2741 -18891 2801 -18621
rect 3071 -18631 3141 -18621
rect 2881 -18681 2911 -18661
rect 2861 -18721 2911 -18681
rect 2971 -18681 3001 -18661
rect 2971 -18721 3021 -18681
rect 2861 -18791 3021 -18721
rect 2861 -18831 2911 -18791
rect 2881 -18851 2911 -18831
rect 2971 -18831 3021 -18791
rect 2971 -18851 3001 -18831
rect 3081 -18891 3141 -18631
rect 2741 -18901 2821 -18891
rect 2741 -18961 2751 -18901
rect 2811 -18911 2821 -18901
rect 3061 -18901 3141 -18891
rect 3061 -18911 3071 -18901
rect 2811 -18961 3071 -18911
rect 3131 -18961 3141 -18901
rect 2741 -18971 3141 -18961
rect 3197 -18551 3597 -18541
rect 3197 -18611 3207 -18551
rect 3267 -18601 3527 -18551
rect 3267 -18611 3277 -18601
rect 3197 -18621 3277 -18611
rect 3517 -18611 3527 -18601
rect 3587 -18611 3597 -18551
rect 3517 -18621 3597 -18611
rect 3197 -18891 3257 -18621
rect 3527 -18631 3597 -18621
rect 3337 -18681 3367 -18661
rect 3317 -18721 3367 -18681
rect 3427 -18681 3457 -18661
rect 3427 -18721 3477 -18681
rect 3317 -18791 3477 -18721
rect 3317 -18831 3367 -18791
rect 3337 -18851 3367 -18831
rect 3427 -18831 3477 -18791
rect 3427 -18851 3457 -18831
rect 3537 -18891 3597 -18631
rect 3197 -18901 3277 -18891
rect 3197 -18961 3207 -18901
rect 3267 -18911 3277 -18901
rect 3517 -18901 3597 -18891
rect 3517 -18911 3527 -18901
rect 3267 -18961 3527 -18911
rect 3587 -18961 3597 -18901
rect 3197 -18971 3597 -18961
rect 3653 -18551 4053 -18541
rect 3653 -18611 3663 -18551
rect 3723 -18601 3983 -18551
rect 3723 -18611 3733 -18601
rect 3653 -18621 3733 -18611
rect 3973 -18611 3983 -18601
rect 4043 -18611 4053 -18551
rect 3973 -18621 4053 -18611
rect 3653 -18891 3713 -18621
rect 3983 -18631 4053 -18621
rect 3793 -18681 3823 -18661
rect 3773 -18721 3823 -18681
rect 3883 -18681 3913 -18661
rect 3883 -18721 3933 -18681
rect 3773 -18791 3933 -18721
rect 3773 -18831 3823 -18791
rect 3793 -18851 3823 -18831
rect 3883 -18831 3933 -18791
rect 3883 -18851 3913 -18831
rect 3993 -18891 4053 -18631
rect 3653 -18901 3733 -18891
rect 3653 -18961 3663 -18901
rect 3723 -18911 3733 -18901
rect 3973 -18901 4053 -18891
rect 3973 -18911 3983 -18901
rect 3723 -18961 3983 -18911
rect 4043 -18961 4053 -18901
rect 3653 -18971 4053 -18961
rect 4111 -18551 4511 -18541
rect 4111 -18611 4121 -18551
rect 4181 -18601 4441 -18551
rect 4181 -18611 4191 -18601
rect 4111 -18621 4191 -18611
rect 4431 -18611 4441 -18601
rect 4501 -18611 4511 -18551
rect 4431 -18621 4511 -18611
rect 4111 -18891 4171 -18621
rect 4441 -18631 4511 -18621
rect 4251 -18681 4281 -18661
rect 4231 -18721 4281 -18681
rect 4341 -18681 4371 -18661
rect 4341 -18721 4391 -18681
rect 4231 -18791 4391 -18721
rect 4231 -18831 4281 -18791
rect 4251 -18851 4281 -18831
rect 4341 -18831 4391 -18791
rect 4341 -18851 4371 -18831
rect 4451 -18891 4511 -18631
rect 4111 -18901 4191 -18891
rect 4111 -18961 4121 -18901
rect 4181 -18911 4191 -18901
rect 4431 -18901 4511 -18891
rect 4431 -18911 4441 -18901
rect 4181 -18961 4441 -18911
rect 4501 -18961 4511 -18901
rect 4111 -18971 4511 -18961
rect 4567 -18551 4967 -18541
rect 4567 -18611 4577 -18551
rect 4637 -18601 4897 -18551
rect 4637 -18611 4647 -18601
rect 4567 -18621 4647 -18611
rect 4887 -18611 4897 -18601
rect 4957 -18611 4967 -18551
rect 4887 -18621 4967 -18611
rect 4567 -18891 4627 -18621
rect 4897 -18631 4967 -18621
rect 4707 -18681 4737 -18661
rect 4687 -18721 4737 -18681
rect 4797 -18681 4827 -18661
rect 4797 -18721 4847 -18681
rect 4687 -18791 4847 -18721
rect 4687 -18831 4737 -18791
rect 4707 -18851 4737 -18831
rect 4797 -18831 4847 -18791
rect 4797 -18851 4827 -18831
rect 4907 -18891 4967 -18631
rect 4567 -18901 4647 -18891
rect 4567 -18961 4577 -18901
rect 4637 -18911 4647 -18901
rect 4887 -18901 4967 -18891
rect 4887 -18911 4897 -18901
rect 4637 -18961 4897 -18911
rect 4957 -18961 4967 -18901
rect 4567 -18971 4967 -18961
rect 5023 -18551 5423 -18541
rect 5023 -18611 5033 -18551
rect 5093 -18601 5353 -18551
rect 5093 -18611 5103 -18601
rect 5023 -18621 5103 -18611
rect 5343 -18611 5353 -18601
rect 5413 -18611 5423 -18551
rect 5343 -18621 5423 -18611
rect 5023 -18891 5083 -18621
rect 5353 -18631 5423 -18621
rect 5163 -18681 5193 -18661
rect 5143 -18721 5193 -18681
rect 5253 -18681 5283 -18661
rect 5253 -18721 5303 -18681
rect 5143 -18791 5303 -18721
rect 5143 -18831 5193 -18791
rect 5163 -18851 5193 -18831
rect 5253 -18831 5303 -18791
rect 5253 -18851 5283 -18831
rect 5363 -18891 5423 -18631
rect 5023 -18901 5103 -18891
rect 5023 -18961 5033 -18901
rect 5093 -18911 5103 -18901
rect 5343 -18901 5423 -18891
rect 5343 -18911 5353 -18901
rect 5093 -18961 5353 -18911
rect 5413 -18961 5423 -18901
rect 5023 -18971 5423 -18961
rect 5481 -18551 5881 -18541
rect 5481 -18611 5491 -18551
rect 5551 -18601 5811 -18551
rect 5551 -18611 5561 -18601
rect 5481 -18621 5561 -18611
rect 5801 -18611 5811 -18601
rect 5871 -18611 5881 -18551
rect 5801 -18621 5881 -18611
rect 5481 -18891 5541 -18621
rect 5811 -18631 5881 -18621
rect 5621 -18681 5651 -18661
rect 5601 -18721 5651 -18681
rect 5711 -18681 5741 -18661
rect 5711 -18721 5761 -18681
rect 5601 -18791 5761 -18721
rect 5601 -18831 5651 -18791
rect 5621 -18851 5651 -18831
rect 5711 -18831 5761 -18791
rect 5711 -18851 5741 -18831
rect 5821 -18891 5881 -18631
rect 5481 -18901 5561 -18891
rect 5481 -18961 5491 -18901
rect 5551 -18911 5561 -18901
rect 5801 -18901 5881 -18891
rect 5801 -18911 5811 -18901
rect 5551 -18961 5811 -18911
rect 5871 -18961 5881 -18901
rect 5481 -18971 5881 -18961
rect 5937 -18551 6337 -18541
rect 5937 -18611 5947 -18551
rect 6007 -18601 6267 -18551
rect 6007 -18611 6017 -18601
rect 5937 -18621 6017 -18611
rect 6257 -18611 6267 -18601
rect 6327 -18611 6337 -18551
rect 6257 -18621 6337 -18611
rect 5937 -18891 5997 -18621
rect 6267 -18631 6337 -18621
rect 6077 -18681 6107 -18661
rect 6057 -18721 6107 -18681
rect 6167 -18681 6197 -18661
rect 6167 -18721 6217 -18681
rect 6057 -18791 6217 -18721
rect 6057 -18831 6107 -18791
rect 6077 -18851 6107 -18831
rect 6167 -18831 6217 -18791
rect 6167 -18851 6197 -18831
rect 6277 -18891 6337 -18631
rect 5937 -18901 6017 -18891
rect 5937 -18961 5947 -18901
rect 6007 -18911 6017 -18901
rect 6257 -18901 6337 -18891
rect 6257 -18911 6267 -18901
rect 6007 -18961 6267 -18911
rect 6327 -18961 6337 -18901
rect 5937 -18971 6337 -18961
rect 6393 -18551 6793 -18541
rect 6393 -18611 6403 -18551
rect 6463 -18601 6723 -18551
rect 6463 -18611 6473 -18601
rect 6393 -18621 6473 -18611
rect 6713 -18611 6723 -18601
rect 6783 -18611 6793 -18551
rect 6713 -18621 6793 -18611
rect 6393 -18891 6453 -18621
rect 6723 -18631 6793 -18621
rect 6533 -18681 6563 -18661
rect 6513 -18721 6563 -18681
rect 6623 -18681 6653 -18661
rect 6623 -18721 6673 -18681
rect 6513 -18791 6673 -18721
rect 6513 -18831 6563 -18791
rect 6533 -18851 6563 -18831
rect 6623 -18831 6673 -18791
rect 6623 -18851 6653 -18831
rect 6733 -18891 6793 -18631
rect 6393 -18901 6473 -18891
rect 6393 -18961 6403 -18901
rect 6463 -18911 6473 -18901
rect 6713 -18901 6793 -18891
rect 6713 -18911 6723 -18901
rect 6463 -18961 6723 -18911
rect 6783 -18961 6793 -18901
rect 6393 -18971 6793 -18961
rect 6851 -18551 7251 -18541
rect 6851 -18611 6861 -18551
rect 6921 -18601 7181 -18551
rect 6921 -18611 6931 -18601
rect 6851 -18621 6931 -18611
rect 7171 -18611 7181 -18601
rect 7241 -18611 7251 -18551
rect 7171 -18621 7251 -18611
rect 6851 -18891 6911 -18621
rect 7181 -18631 7251 -18621
rect 6991 -18681 7021 -18661
rect 6971 -18721 7021 -18681
rect 7081 -18681 7111 -18661
rect 7081 -18721 7131 -18681
rect 6971 -18791 7131 -18721
rect 6971 -18831 7021 -18791
rect 6991 -18851 7021 -18831
rect 7081 -18831 7131 -18791
rect 7081 -18851 7111 -18831
rect 7191 -18891 7251 -18631
rect 6851 -18901 6931 -18891
rect 6851 -18961 6861 -18901
rect 6921 -18911 6931 -18901
rect 7171 -18901 7251 -18891
rect 7171 -18911 7181 -18901
rect 6921 -18961 7181 -18911
rect 7241 -18961 7251 -18901
rect 6851 -18971 7251 -18961
rect 7307 -18551 7707 -18541
rect 7307 -18611 7317 -18551
rect 7377 -18601 7637 -18551
rect 7377 -18611 7387 -18601
rect 7307 -18621 7387 -18611
rect 7627 -18611 7637 -18601
rect 7697 -18611 7707 -18551
rect 7627 -18621 7707 -18611
rect 7307 -18891 7367 -18621
rect 7637 -18631 7707 -18621
rect 7447 -18681 7477 -18661
rect 7427 -18721 7477 -18681
rect 7537 -18681 7567 -18661
rect 7537 -18721 7587 -18681
rect 7427 -18791 7587 -18721
rect 7427 -18831 7477 -18791
rect 7447 -18851 7477 -18831
rect 7537 -18831 7587 -18791
rect 7537 -18851 7567 -18831
rect 7647 -18891 7707 -18631
rect 7307 -18901 7387 -18891
rect 7307 -18961 7317 -18901
rect 7377 -18911 7387 -18901
rect 7627 -18901 7707 -18891
rect 7627 -18911 7637 -18901
rect 7377 -18961 7637 -18911
rect 7697 -18961 7707 -18901
rect 7307 -18971 7707 -18961
rect 7763 -18551 8163 -18541
rect 7763 -18611 7773 -18551
rect 7833 -18601 8093 -18551
rect 7833 -18611 7843 -18601
rect 7763 -18621 7843 -18611
rect 8083 -18611 8093 -18601
rect 8153 -18611 8163 -18551
rect 8083 -18621 8163 -18611
rect 7763 -18891 7823 -18621
rect 8093 -18631 8163 -18621
rect 7903 -18681 7933 -18661
rect 7883 -18721 7933 -18681
rect 7993 -18681 8023 -18661
rect 7993 -18721 8043 -18681
rect 7883 -18791 8043 -18721
rect 7883 -18831 7933 -18791
rect 7903 -18851 7933 -18831
rect 7993 -18831 8043 -18791
rect 7993 -18851 8023 -18831
rect 8103 -18891 8163 -18631
rect 7763 -18901 7843 -18891
rect 7763 -18961 7773 -18901
rect 7833 -18911 7843 -18901
rect 8083 -18901 8163 -18891
rect 8083 -18911 8093 -18901
rect 7833 -18961 8093 -18911
rect 8153 -18961 8163 -18901
rect 7763 -18971 8163 -18961
rect 8237 -18551 8637 -18541
rect 8237 -18611 8247 -18551
rect 8307 -18601 8567 -18551
rect 8307 -18611 8317 -18601
rect 8237 -18621 8317 -18611
rect 8557 -18611 8567 -18601
rect 8627 -18611 8637 -18551
rect 8557 -18621 8637 -18611
rect 8237 -18891 8297 -18621
rect 8567 -18631 8637 -18621
rect 8377 -18681 8407 -18661
rect 8357 -18721 8407 -18681
rect 8467 -18681 8497 -18661
rect 8467 -18721 8517 -18681
rect 8357 -18791 8517 -18721
rect 8357 -18831 8407 -18791
rect 8377 -18851 8407 -18831
rect 8467 -18831 8517 -18791
rect 8467 -18851 8497 -18831
rect 8577 -18891 8637 -18631
rect 8237 -18901 8317 -18891
rect 8237 -18961 8247 -18901
rect 8307 -18911 8317 -18901
rect 8557 -18901 8637 -18891
rect 8557 -18911 8567 -18901
rect 8307 -18961 8567 -18911
rect 8627 -18961 8637 -18901
rect 8237 -18971 8637 -18961
rect 8693 -18551 9093 -18541
rect 8693 -18611 8703 -18551
rect 8763 -18601 9023 -18551
rect 8763 -18611 8773 -18601
rect 8693 -18621 8773 -18611
rect 9013 -18611 9023 -18601
rect 9083 -18611 9093 -18551
rect 9013 -18621 9093 -18611
rect 8693 -18891 8753 -18621
rect 9023 -18631 9093 -18621
rect 8833 -18681 8863 -18661
rect 8813 -18721 8863 -18681
rect 8923 -18681 8953 -18661
rect 8923 -18721 8973 -18681
rect 8813 -18791 8973 -18721
rect 8813 -18831 8863 -18791
rect 8833 -18851 8863 -18831
rect 8923 -18831 8973 -18791
rect 8923 -18851 8953 -18831
rect 9033 -18891 9093 -18631
rect 8693 -18901 8773 -18891
rect 8693 -18961 8703 -18901
rect 8763 -18911 8773 -18901
rect 9013 -18901 9093 -18891
rect 9013 -18911 9023 -18901
rect 8763 -18961 9023 -18911
rect 9083 -18961 9093 -18901
rect 8693 -18971 9093 -18961
rect 9151 -18551 9551 -18541
rect 9151 -18611 9161 -18551
rect 9221 -18601 9481 -18551
rect 9221 -18611 9231 -18601
rect 9151 -18621 9231 -18611
rect 9471 -18611 9481 -18601
rect 9541 -18611 9551 -18551
rect 9471 -18621 9551 -18611
rect 9151 -18891 9211 -18621
rect 9481 -18631 9551 -18621
rect 9291 -18681 9321 -18661
rect 9271 -18721 9321 -18681
rect 9381 -18681 9411 -18661
rect 9381 -18721 9431 -18681
rect 9271 -18791 9431 -18721
rect 9271 -18831 9321 -18791
rect 9291 -18851 9321 -18831
rect 9381 -18831 9431 -18791
rect 9381 -18851 9411 -18831
rect 9491 -18891 9551 -18631
rect 9151 -18901 9231 -18891
rect 9151 -18961 9161 -18901
rect 9221 -18911 9231 -18901
rect 9471 -18901 9551 -18891
rect 9471 -18911 9481 -18901
rect 9221 -18961 9481 -18911
rect 9541 -18961 9551 -18901
rect 9151 -18971 9551 -18961
rect 9607 -18551 10007 -18541
rect 9607 -18611 9617 -18551
rect 9677 -18601 9937 -18551
rect 9677 -18611 9687 -18601
rect 9607 -18621 9687 -18611
rect 9927 -18611 9937 -18601
rect 9997 -18611 10007 -18551
rect 9927 -18621 10007 -18611
rect 9607 -18891 9667 -18621
rect 9937 -18631 10007 -18621
rect 9747 -18681 9777 -18661
rect 9727 -18721 9777 -18681
rect 9837 -18681 9867 -18661
rect 9837 -18721 9887 -18681
rect 9727 -18791 9887 -18721
rect 9727 -18831 9777 -18791
rect 9747 -18851 9777 -18831
rect 9837 -18831 9887 -18791
rect 9837 -18851 9867 -18831
rect 9947 -18891 10007 -18631
rect 9607 -18901 9687 -18891
rect 9607 -18961 9617 -18901
rect 9677 -18911 9687 -18901
rect 9927 -18901 10007 -18891
rect 9927 -18911 9937 -18901
rect 9677 -18961 9937 -18911
rect 9997 -18961 10007 -18901
rect 9607 -18971 10007 -18961
rect 10063 -18551 10463 -18541
rect 10063 -18611 10073 -18551
rect 10133 -18601 10393 -18551
rect 10133 -18611 10143 -18601
rect 10063 -18621 10143 -18611
rect 10383 -18611 10393 -18601
rect 10453 -18611 10463 -18551
rect 10383 -18621 10463 -18611
rect 10063 -18891 10123 -18621
rect 10393 -18631 10463 -18621
rect 10203 -18681 10233 -18661
rect 10183 -18721 10233 -18681
rect 10293 -18681 10323 -18661
rect 10293 -18721 10343 -18681
rect 10183 -18791 10343 -18721
rect 10183 -18831 10233 -18791
rect 10203 -18851 10233 -18831
rect 10293 -18831 10343 -18791
rect 10293 -18851 10323 -18831
rect 10403 -18891 10463 -18631
rect 10063 -18901 10143 -18891
rect 10063 -18961 10073 -18901
rect 10133 -18911 10143 -18901
rect 10383 -18901 10463 -18891
rect 10383 -18911 10393 -18901
rect 10133 -18961 10393 -18911
rect 10453 -18961 10463 -18901
rect 10063 -18971 10463 -18961
rect 10521 -18551 10921 -18541
rect 10521 -18611 10531 -18551
rect 10591 -18601 10851 -18551
rect 10591 -18611 10601 -18601
rect 10521 -18621 10601 -18611
rect 10841 -18611 10851 -18601
rect 10911 -18611 10921 -18551
rect 10841 -18621 10921 -18611
rect 10521 -18891 10581 -18621
rect 10851 -18631 10921 -18621
rect 10661 -18681 10691 -18661
rect 10641 -18721 10691 -18681
rect 10751 -18681 10781 -18661
rect 10751 -18721 10801 -18681
rect 10641 -18791 10801 -18721
rect 10641 -18831 10691 -18791
rect 10661 -18851 10691 -18831
rect 10751 -18831 10801 -18791
rect 10751 -18851 10781 -18831
rect 10861 -18891 10921 -18631
rect 10521 -18901 10601 -18891
rect 10521 -18961 10531 -18901
rect 10591 -18911 10601 -18901
rect 10841 -18901 10921 -18891
rect 10841 -18911 10851 -18901
rect 10591 -18961 10851 -18911
rect 10911 -18961 10921 -18901
rect 10521 -18971 10921 -18961
rect 10977 -18551 11377 -18541
rect 10977 -18611 10987 -18551
rect 11047 -18601 11307 -18551
rect 11047 -18611 11057 -18601
rect 10977 -18621 11057 -18611
rect 11297 -18611 11307 -18601
rect 11367 -18611 11377 -18551
rect 11297 -18621 11377 -18611
rect 10977 -18891 11037 -18621
rect 11307 -18631 11377 -18621
rect 11117 -18681 11147 -18661
rect 11097 -18721 11147 -18681
rect 11207 -18681 11237 -18661
rect 11207 -18721 11257 -18681
rect 11097 -18791 11257 -18721
rect 11097 -18831 11147 -18791
rect 11117 -18851 11147 -18831
rect 11207 -18831 11257 -18791
rect 11207 -18851 11237 -18831
rect 11317 -18891 11377 -18631
rect 10977 -18901 11057 -18891
rect 10977 -18961 10987 -18901
rect 11047 -18911 11057 -18901
rect 11297 -18901 11377 -18891
rect 11297 -18911 11307 -18901
rect 11047 -18961 11307 -18911
rect 11367 -18961 11377 -18901
rect 10977 -18971 11377 -18961
rect 11433 -18551 11833 -18541
rect 11433 -18611 11443 -18551
rect 11503 -18601 11763 -18551
rect 11503 -18611 11513 -18601
rect 11433 -18621 11513 -18611
rect 11753 -18611 11763 -18601
rect 11823 -18611 11833 -18551
rect 11753 -18621 11833 -18611
rect 11433 -18891 11493 -18621
rect 11763 -18631 11833 -18621
rect 11573 -18681 11603 -18661
rect 11553 -18721 11603 -18681
rect 11663 -18681 11693 -18661
rect 11663 -18721 11713 -18681
rect 11553 -18791 11713 -18721
rect 11553 -18831 11603 -18791
rect 11573 -18851 11603 -18831
rect 11663 -18831 11713 -18791
rect 11663 -18851 11693 -18831
rect 11773 -18891 11833 -18631
rect 11433 -18901 11513 -18891
rect 11433 -18961 11443 -18901
rect 11503 -18911 11513 -18901
rect 11753 -18901 11833 -18891
rect 11753 -18911 11763 -18901
rect 11503 -18961 11763 -18911
rect 11823 -18961 11833 -18901
rect 11433 -18971 11833 -18961
rect 11891 -18551 12291 -18541
rect 11891 -18611 11901 -18551
rect 11961 -18601 12221 -18551
rect 11961 -18611 11971 -18601
rect 11891 -18621 11971 -18611
rect 12211 -18611 12221 -18601
rect 12281 -18611 12291 -18551
rect 12211 -18621 12291 -18611
rect 11891 -18891 11951 -18621
rect 12221 -18631 12291 -18621
rect 12031 -18681 12061 -18661
rect 12011 -18721 12061 -18681
rect 12121 -18681 12151 -18661
rect 12121 -18721 12171 -18681
rect 12011 -18791 12171 -18721
rect 12011 -18831 12061 -18791
rect 12031 -18851 12061 -18831
rect 12121 -18831 12171 -18791
rect 12121 -18851 12151 -18831
rect 12231 -18891 12291 -18631
rect 11891 -18901 11971 -18891
rect 11891 -18961 11901 -18901
rect 11961 -18911 11971 -18901
rect 12211 -18901 12291 -18891
rect 12211 -18911 12221 -18901
rect 11961 -18961 12221 -18911
rect 12281 -18961 12291 -18901
rect 11891 -18971 12291 -18961
rect 12347 -18551 12747 -18541
rect 12347 -18611 12357 -18551
rect 12417 -18601 12677 -18551
rect 12417 -18611 12427 -18601
rect 12347 -18621 12427 -18611
rect 12667 -18611 12677 -18601
rect 12737 -18611 12747 -18551
rect 12667 -18621 12747 -18611
rect 12347 -18891 12407 -18621
rect 12677 -18631 12747 -18621
rect 12487 -18681 12517 -18661
rect 12467 -18721 12517 -18681
rect 12577 -18681 12607 -18661
rect 12577 -18721 12627 -18681
rect 12467 -18791 12627 -18721
rect 12467 -18831 12517 -18791
rect 12487 -18851 12517 -18831
rect 12577 -18831 12627 -18791
rect 12577 -18851 12607 -18831
rect 12687 -18891 12747 -18631
rect 12347 -18901 12427 -18891
rect 12347 -18961 12357 -18901
rect 12417 -18911 12427 -18901
rect 12667 -18901 12747 -18891
rect 12667 -18911 12677 -18901
rect 12417 -18961 12677 -18911
rect 12737 -18961 12747 -18901
rect 12347 -18971 12747 -18961
rect 12803 -18551 13203 -18541
rect 12803 -18611 12813 -18551
rect 12873 -18601 13133 -18551
rect 12873 -18611 12883 -18601
rect 12803 -18621 12883 -18611
rect 13123 -18611 13133 -18601
rect 13193 -18611 13203 -18551
rect 13123 -18621 13203 -18611
rect 12803 -18891 12863 -18621
rect 13133 -18631 13203 -18621
rect 12943 -18681 12973 -18661
rect 12923 -18721 12973 -18681
rect 13033 -18681 13063 -18661
rect 13033 -18721 13083 -18681
rect 12923 -18791 13083 -18721
rect 12923 -18831 12973 -18791
rect 12943 -18851 12973 -18831
rect 13033 -18831 13083 -18791
rect 13033 -18851 13063 -18831
rect 13143 -18891 13203 -18631
rect 12803 -18901 12883 -18891
rect 12803 -18961 12813 -18901
rect 12873 -18911 12883 -18901
rect 13123 -18901 13203 -18891
rect 13123 -18911 13133 -18901
rect 12873 -18961 13133 -18911
rect 13193 -18961 13203 -18901
rect 12803 -18971 13203 -18961
rect 13261 -18551 13661 -18541
rect 13261 -18611 13271 -18551
rect 13331 -18601 13591 -18551
rect 13331 -18611 13341 -18601
rect 13261 -18621 13341 -18611
rect 13581 -18611 13591 -18601
rect 13651 -18611 13661 -18551
rect 13581 -18621 13661 -18611
rect 13261 -18891 13321 -18621
rect 13591 -18631 13661 -18621
rect 13401 -18681 13431 -18661
rect 13381 -18721 13431 -18681
rect 13491 -18681 13521 -18661
rect 13491 -18721 13541 -18681
rect 13381 -18791 13541 -18721
rect 13381 -18831 13431 -18791
rect 13401 -18851 13431 -18831
rect 13491 -18831 13541 -18791
rect 13491 -18851 13521 -18831
rect 13601 -18891 13661 -18631
rect 13261 -18901 13341 -18891
rect 13261 -18961 13271 -18901
rect 13331 -18911 13341 -18901
rect 13581 -18901 13661 -18891
rect 13581 -18911 13591 -18901
rect 13331 -18961 13591 -18911
rect 13651 -18961 13661 -18901
rect 13261 -18971 13661 -18961
rect 13717 -18551 14117 -18541
rect 13717 -18611 13727 -18551
rect 13787 -18601 14047 -18551
rect 13787 -18611 13797 -18601
rect 13717 -18621 13797 -18611
rect 14037 -18611 14047 -18601
rect 14107 -18611 14117 -18551
rect 14037 -18621 14117 -18611
rect 13717 -18891 13777 -18621
rect 14047 -18631 14117 -18621
rect 13857 -18681 13887 -18661
rect 13837 -18721 13887 -18681
rect 13947 -18681 13977 -18661
rect 13947 -18721 13997 -18681
rect 13837 -18791 13997 -18721
rect 13837 -18831 13887 -18791
rect 13857 -18851 13887 -18831
rect 13947 -18831 13997 -18791
rect 13947 -18851 13977 -18831
rect 14057 -18891 14117 -18631
rect 13717 -18901 13797 -18891
rect 13717 -18961 13727 -18901
rect 13787 -18911 13797 -18901
rect 14037 -18901 14117 -18891
rect 14037 -18911 14047 -18901
rect 13787 -18961 14047 -18911
rect 14107 -18961 14117 -18901
rect 13717 -18971 14117 -18961
rect 14173 -18551 14573 -18541
rect 14173 -18611 14183 -18551
rect 14243 -18601 14503 -18551
rect 14243 -18611 14253 -18601
rect 14173 -18621 14253 -18611
rect 14493 -18611 14503 -18601
rect 14563 -18611 14573 -18551
rect 14493 -18621 14573 -18611
rect 14173 -18891 14233 -18621
rect 14503 -18631 14573 -18621
rect 14313 -18681 14343 -18661
rect 14293 -18721 14343 -18681
rect 14403 -18681 14433 -18661
rect 14403 -18721 14453 -18681
rect 14293 -18791 14453 -18721
rect 14293 -18831 14343 -18791
rect 14313 -18851 14343 -18831
rect 14403 -18831 14453 -18791
rect 14403 -18851 14433 -18831
rect 14513 -18891 14573 -18631
rect 14173 -18901 14253 -18891
rect 14173 -18961 14183 -18901
rect 14243 -18911 14253 -18901
rect 14493 -18901 14573 -18891
rect 14493 -18911 14503 -18901
rect 14243 -18961 14503 -18911
rect 14563 -18961 14573 -18901
rect 14173 -18971 14573 -18961
rect 14631 -18551 15031 -18541
rect 14631 -18611 14641 -18551
rect 14701 -18601 14961 -18551
rect 14701 -18611 14711 -18601
rect 14631 -18621 14711 -18611
rect 14951 -18611 14961 -18601
rect 15021 -18611 15031 -18551
rect 14951 -18621 15031 -18611
rect 14631 -18891 14691 -18621
rect 14961 -18631 15031 -18621
rect 14771 -18681 14801 -18661
rect 14751 -18721 14801 -18681
rect 14861 -18681 14891 -18661
rect 14861 -18721 14911 -18681
rect 14751 -18791 14911 -18721
rect 14751 -18831 14801 -18791
rect 14771 -18851 14801 -18831
rect 14861 -18831 14911 -18791
rect 14861 -18851 14891 -18831
rect 14971 -18891 15031 -18631
rect 14631 -18901 14711 -18891
rect 14631 -18961 14641 -18901
rect 14701 -18911 14711 -18901
rect 14951 -18901 15031 -18891
rect 14951 -18911 14961 -18901
rect 14701 -18961 14961 -18911
rect 15021 -18961 15031 -18901
rect 14631 -18971 15031 -18961
rect 15087 -18551 15487 -18541
rect 15087 -18611 15097 -18551
rect 15157 -18601 15417 -18551
rect 15157 -18611 15167 -18601
rect 15087 -18621 15167 -18611
rect 15407 -18611 15417 -18601
rect 15477 -18611 15487 -18551
rect 15407 -18621 15487 -18611
rect 15087 -18891 15147 -18621
rect 15417 -18631 15487 -18621
rect 15227 -18681 15257 -18661
rect 15207 -18721 15257 -18681
rect 15317 -18681 15347 -18661
rect 15317 -18721 15367 -18681
rect 15207 -18791 15367 -18721
rect 15207 -18831 15257 -18791
rect 15227 -18851 15257 -18831
rect 15317 -18831 15367 -18791
rect 15317 -18851 15347 -18831
rect 15427 -18891 15487 -18631
rect 15087 -18901 15167 -18891
rect 15087 -18961 15097 -18901
rect 15157 -18911 15167 -18901
rect 15407 -18901 15487 -18891
rect 15407 -18911 15417 -18901
rect 15157 -18961 15417 -18911
rect 15477 -18961 15487 -18901
rect 15087 -18971 15487 -18961
rect 1 -19043 401 -19033
rect 1 -19103 11 -19043
rect 71 -19093 331 -19043
rect 71 -19103 81 -19093
rect 1 -19113 81 -19103
rect 321 -19103 331 -19093
rect 391 -19103 401 -19043
rect 321 -19113 401 -19103
rect 1 -19383 61 -19113
rect 331 -19123 401 -19113
rect 141 -19173 171 -19153
rect 121 -19213 171 -19173
rect 231 -19173 261 -19153
rect 231 -19213 281 -19173
rect 121 -19283 281 -19213
rect 121 -19323 171 -19283
rect 141 -19343 171 -19323
rect 231 -19323 281 -19283
rect 231 -19343 261 -19323
rect 341 -19383 401 -19123
rect 1 -19393 81 -19383
rect 1 -19453 11 -19393
rect 71 -19403 81 -19393
rect 321 -19393 401 -19383
rect 321 -19403 331 -19393
rect 71 -19453 331 -19403
rect 391 -19453 401 -19393
rect 1 -19463 401 -19453
rect 457 -19043 857 -19033
rect 457 -19103 467 -19043
rect 527 -19093 787 -19043
rect 527 -19103 537 -19093
rect 457 -19113 537 -19103
rect 777 -19103 787 -19093
rect 847 -19103 857 -19043
rect 777 -19113 857 -19103
rect 457 -19383 517 -19113
rect 787 -19123 857 -19113
rect 597 -19173 627 -19153
rect 577 -19213 627 -19173
rect 687 -19173 717 -19153
rect 687 -19213 737 -19173
rect 577 -19283 737 -19213
rect 577 -19323 627 -19283
rect 597 -19343 627 -19323
rect 687 -19323 737 -19283
rect 687 -19343 717 -19323
rect 797 -19383 857 -19123
rect 457 -19393 537 -19383
rect 457 -19453 467 -19393
rect 527 -19403 537 -19393
rect 777 -19393 857 -19383
rect 777 -19403 787 -19393
rect 527 -19453 787 -19403
rect 847 -19453 857 -19393
rect 457 -19463 857 -19453
rect 913 -19043 1313 -19033
rect 913 -19103 923 -19043
rect 983 -19093 1243 -19043
rect 983 -19103 993 -19093
rect 913 -19113 993 -19103
rect 1233 -19103 1243 -19093
rect 1303 -19103 1313 -19043
rect 1233 -19113 1313 -19103
rect 913 -19383 973 -19113
rect 1243 -19123 1313 -19113
rect 1053 -19173 1083 -19153
rect 1033 -19213 1083 -19173
rect 1143 -19173 1173 -19153
rect 1143 -19213 1193 -19173
rect 1033 -19283 1193 -19213
rect 1033 -19323 1083 -19283
rect 1053 -19343 1083 -19323
rect 1143 -19323 1193 -19283
rect 1143 -19343 1173 -19323
rect 1253 -19383 1313 -19123
rect 913 -19393 993 -19383
rect 913 -19453 923 -19393
rect 983 -19403 993 -19393
rect 1233 -19393 1313 -19383
rect 1233 -19403 1243 -19393
rect 983 -19453 1243 -19403
rect 1303 -19453 1313 -19393
rect 913 -19463 1313 -19453
rect 1371 -19043 1771 -19033
rect 1371 -19103 1381 -19043
rect 1441 -19093 1701 -19043
rect 1441 -19103 1451 -19093
rect 1371 -19113 1451 -19103
rect 1691 -19103 1701 -19093
rect 1761 -19103 1771 -19043
rect 1691 -19113 1771 -19103
rect 1371 -19383 1431 -19113
rect 1701 -19123 1771 -19113
rect 1511 -19173 1541 -19153
rect 1491 -19213 1541 -19173
rect 1601 -19173 1631 -19153
rect 1601 -19213 1651 -19173
rect 1491 -19283 1651 -19213
rect 1491 -19323 1541 -19283
rect 1511 -19343 1541 -19323
rect 1601 -19323 1651 -19283
rect 1601 -19343 1631 -19323
rect 1711 -19383 1771 -19123
rect 1371 -19393 1451 -19383
rect 1371 -19453 1381 -19393
rect 1441 -19403 1451 -19393
rect 1691 -19393 1771 -19383
rect 1691 -19403 1701 -19393
rect 1441 -19453 1701 -19403
rect 1761 -19453 1771 -19393
rect 1371 -19463 1771 -19453
rect 1827 -19043 2227 -19033
rect 1827 -19103 1837 -19043
rect 1897 -19093 2157 -19043
rect 1897 -19103 1907 -19093
rect 1827 -19113 1907 -19103
rect 2147 -19103 2157 -19093
rect 2217 -19103 2227 -19043
rect 2147 -19113 2227 -19103
rect 1827 -19383 1887 -19113
rect 2157 -19123 2227 -19113
rect 1967 -19173 1997 -19153
rect 1947 -19213 1997 -19173
rect 2057 -19173 2087 -19153
rect 2057 -19213 2107 -19173
rect 1947 -19283 2107 -19213
rect 1947 -19323 1997 -19283
rect 1967 -19343 1997 -19323
rect 2057 -19323 2107 -19283
rect 2057 -19343 2087 -19323
rect 2167 -19383 2227 -19123
rect 1827 -19393 1907 -19383
rect 1827 -19453 1837 -19393
rect 1897 -19403 1907 -19393
rect 2147 -19393 2227 -19383
rect 2147 -19403 2157 -19393
rect 1897 -19453 2157 -19403
rect 2217 -19453 2227 -19393
rect 1827 -19463 2227 -19453
rect 2283 -19043 2683 -19033
rect 2283 -19103 2293 -19043
rect 2353 -19093 2613 -19043
rect 2353 -19103 2363 -19093
rect 2283 -19113 2363 -19103
rect 2603 -19103 2613 -19093
rect 2673 -19103 2683 -19043
rect 2603 -19113 2683 -19103
rect 2283 -19383 2343 -19113
rect 2613 -19123 2683 -19113
rect 2423 -19173 2453 -19153
rect 2403 -19213 2453 -19173
rect 2513 -19173 2543 -19153
rect 2513 -19213 2563 -19173
rect 2403 -19283 2563 -19213
rect 2403 -19323 2453 -19283
rect 2423 -19343 2453 -19323
rect 2513 -19323 2563 -19283
rect 2513 -19343 2543 -19323
rect 2623 -19383 2683 -19123
rect 2283 -19393 2363 -19383
rect 2283 -19453 2293 -19393
rect 2353 -19403 2363 -19393
rect 2603 -19393 2683 -19383
rect 2603 -19403 2613 -19393
rect 2353 -19453 2613 -19403
rect 2673 -19453 2683 -19393
rect 2283 -19463 2683 -19453
rect 2741 -19043 3141 -19033
rect 2741 -19103 2751 -19043
rect 2811 -19093 3071 -19043
rect 2811 -19103 2821 -19093
rect 2741 -19113 2821 -19103
rect 3061 -19103 3071 -19093
rect 3131 -19103 3141 -19043
rect 3061 -19113 3141 -19103
rect 2741 -19383 2801 -19113
rect 3071 -19123 3141 -19113
rect 2881 -19173 2911 -19153
rect 2861 -19213 2911 -19173
rect 2971 -19173 3001 -19153
rect 2971 -19213 3021 -19173
rect 2861 -19283 3021 -19213
rect 2861 -19323 2911 -19283
rect 2881 -19343 2911 -19323
rect 2971 -19323 3021 -19283
rect 2971 -19343 3001 -19323
rect 3081 -19383 3141 -19123
rect 2741 -19393 2821 -19383
rect 2741 -19453 2751 -19393
rect 2811 -19403 2821 -19393
rect 3061 -19393 3141 -19383
rect 3061 -19403 3071 -19393
rect 2811 -19453 3071 -19403
rect 3131 -19453 3141 -19393
rect 2741 -19463 3141 -19453
rect 3197 -19043 3597 -19033
rect 3197 -19103 3207 -19043
rect 3267 -19093 3527 -19043
rect 3267 -19103 3277 -19093
rect 3197 -19113 3277 -19103
rect 3517 -19103 3527 -19093
rect 3587 -19103 3597 -19043
rect 3517 -19113 3597 -19103
rect 3197 -19383 3257 -19113
rect 3527 -19123 3597 -19113
rect 3337 -19173 3367 -19153
rect 3317 -19213 3367 -19173
rect 3427 -19173 3457 -19153
rect 3427 -19213 3477 -19173
rect 3317 -19283 3477 -19213
rect 3317 -19323 3367 -19283
rect 3337 -19343 3367 -19323
rect 3427 -19323 3477 -19283
rect 3427 -19343 3457 -19323
rect 3537 -19383 3597 -19123
rect 3197 -19393 3277 -19383
rect 3197 -19453 3207 -19393
rect 3267 -19403 3277 -19393
rect 3517 -19393 3597 -19383
rect 3517 -19403 3527 -19393
rect 3267 -19453 3527 -19403
rect 3587 -19453 3597 -19393
rect 3197 -19463 3597 -19453
rect 3653 -19043 4053 -19033
rect 3653 -19103 3663 -19043
rect 3723 -19093 3983 -19043
rect 3723 -19103 3733 -19093
rect 3653 -19113 3733 -19103
rect 3973 -19103 3983 -19093
rect 4043 -19103 4053 -19043
rect 3973 -19113 4053 -19103
rect 3653 -19383 3713 -19113
rect 3983 -19123 4053 -19113
rect 3793 -19173 3823 -19153
rect 3773 -19213 3823 -19173
rect 3883 -19173 3913 -19153
rect 3883 -19213 3933 -19173
rect 3773 -19283 3933 -19213
rect 3773 -19323 3823 -19283
rect 3793 -19343 3823 -19323
rect 3883 -19323 3933 -19283
rect 3883 -19343 3913 -19323
rect 3993 -19383 4053 -19123
rect 3653 -19393 3733 -19383
rect 3653 -19453 3663 -19393
rect 3723 -19403 3733 -19393
rect 3973 -19393 4053 -19383
rect 3973 -19403 3983 -19393
rect 3723 -19453 3983 -19403
rect 4043 -19453 4053 -19393
rect 3653 -19463 4053 -19453
rect 4111 -19043 4511 -19033
rect 4111 -19103 4121 -19043
rect 4181 -19093 4441 -19043
rect 4181 -19103 4191 -19093
rect 4111 -19113 4191 -19103
rect 4431 -19103 4441 -19093
rect 4501 -19103 4511 -19043
rect 4431 -19113 4511 -19103
rect 4111 -19383 4171 -19113
rect 4441 -19123 4511 -19113
rect 4251 -19173 4281 -19153
rect 4231 -19213 4281 -19173
rect 4341 -19173 4371 -19153
rect 4341 -19213 4391 -19173
rect 4231 -19283 4391 -19213
rect 4231 -19323 4281 -19283
rect 4251 -19343 4281 -19323
rect 4341 -19323 4391 -19283
rect 4341 -19343 4371 -19323
rect 4451 -19383 4511 -19123
rect 4111 -19393 4191 -19383
rect 4111 -19453 4121 -19393
rect 4181 -19403 4191 -19393
rect 4431 -19393 4511 -19383
rect 4431 -19403 4441 -19393
rect 4181 -19453 4441 -19403
rect 4501 -19453 4511 -19393
rect 4111 -19463 4511 -19453
rect 4567 -19043 4967 -19033
rect 4567 -19103 4577 -19043
rect 4637 -19093 4897 -19043
rect 4637 -19103 4647 -19093
rect 4567 -19113 4647 -19103
rect 4887 -19103 4897 -19093
rect 4957 -19103 4967 -19043
rect 4887 -19113 4967 -19103
rect 4567 -19383 4627 -19113
rect 4897 -19123 4967 -19113
rect 4707 -19173 4737 -19153
rect 4687 -19213 4737 -19173
rect 4797 -19173 4827 -19153
rect 4797 -19213 4847 -19173
rect 4687 -19283 4847 -19213
rect 4687 -19323 4737 -19283
rect 4707 -19343 4737 -19323
rect 4797 -19323 4847 -19283
rect 4797 -19343 4827 -19323
rect 4907 -19383 4967 -19123
rect 4567 -19393 4647 -19383
rect 4567 -19453 4577 -19393
rect 4637 -19403 4647 -19393
rect 4887 -19393 4967 -19383
rect 4887 -19403 4897 -19393
rect 4637 -19453 4897 -19403
rect 4957 -19453 4967 -19393
rect 4567 -19463 4967 -19453
rect 5023 -19043 5423 -19033
rect 5023 -19103 5033 -19043
rect 5093 -19093 5353 -19043
rect 5093 -19103 5103 -19093
rect 5023 -19113 5103 -19103
rect 5343 -19103 5353 -19093
rect 5413 -19103 5423 -19043
rect 5343 -19113 5423 -19103
rect 5023 -19383 5083 -19113
rect 5353 -19123 5423 -19113
rect 5163 -19173 5193 -19153
rect 5143 -19213 5193 -19173
rect 5253 -19173 5283 -19153
rect 5253 -19213 5303 -19173
rect 5143 -19283 5303 -19213
rect 5143 -19323 5193 -19283
rect 5163 -19343 5193 -19323
rect 5253 -19323 5303 -19283
rect 5253 -19343 5283 -19323
rect 5363 -19383 5423 -19123
rect 5023 -19393 5103 -19383
rect 5023 -19453 5033 -19393
rect 5093 -19403 5103 -19393
rect 5343 -19393 5423 -19383
rect 5343 -19403 5353 -19393
rect 5093 -19453 5353 -19403
rect 5413 -19453 5423 -19393
rect 5023 -19463 5423 -19453
rect 5481 -19043 5881 -19033
rect 5481 -19103 5491 -19043
rect 5551 -19093 5811 -19043
rect 5551 -19103 5561 -19093
rect 5481 -19113 5561 -19103
rect 5801 -19103 5811 -19093
rect 5871 -19103 5881 -19043
rect 5801 -19113 5881 -19103
rect 5481 -19383 5541 -19113
rect 5811 -19123 5881 -19113
rect 5621 -19173 5651 -19153
rect 5601 -19213 5651 -19173
rect 5711 -19173 5741 -19153
rect 5711 -19213 5761 -19173
rect 5601 -19283 5761 -19213
rect 5601 -19323 5651 -19283
rect 5621 -19343 5651 -19323
rect 5711 -19323 5761 -19283
rect 5711 -19343 5741 -19323
rect 5821 -19383 5881 -19123
rect 5481 -19393 5561 -19383
rect 5481 -19453 5491 -19393
rect 5551 -19403 5561 -19393
rect 5801 -19393 5881 -19383
rect 5801 -19403 5811 -19393
rect 5551 -19453 5811 -19403
rect 5871 -19453 5881 -19393
rect 5481 -19463 5881 -19453
rect 5937 -19043 6337 -19033
rect 5937 -19103 5947 -19043
rect 6007 -19093 6267 -19043
rect 6007 -19103 6017 -19093
rect 5937 -19113 6017 -19103
rect 6257 -19103 6267 -19093
rect 6327 -19103 6337 -19043
rect 6257 -19113 6337 -19103
rect 5937 -19383 5997 -19113
rect 6267 -19123 6337 -19113
rect 6077 -19173 6107 -19153
rect 6057 -19213 6107 -19173
rect 6167 -19173 6197 -19153
rect 6167 -19213 6217 -19173
rect 6057 -19283 6217 -19213
rect 6057 -19323 6107 -19283
rect 6077 -19343 6107 -19323
rect 6167 -19323 6217 -19283
rect 6167 -19343 6197 -19323
rect 6277 -19383 6337 -19123
rect 5937 -19393 6017 -19383
rect 5937 -19453 5947 -19393
rect 6007 -19403 6017 -19393
rect 6257 -19393 6337 -19383
rect 6257 -19403 6267 -19393
rect 6007 -19453 6267 -19403
rect 6327 -19453 6337 -19393
rect 5937 -19463 6337 -19453
rect 6393 -19043 6793 -19033
rect 6393 -19103 6403 -19043
rect 6463 -19093 6723 -19043
rect 6463 -19103 6473 -19093
rect 6393 -19113 6473 -19103
rect 6713 -19103 6723 -19093
rect 6783 -19103 6793 -19043
rect 6713 -19113 6793 -19103
rect 6393 -19383 6453 -19113
rect 6723 -19123 6793 -19113
rect 6533 -19173 6563 -19153
rect 6513 -19213 6563 -19173
rect 6623 -19173 6653 -19153
rect 6623 -19213 6673 -19173
rect 6513 -19283 6673 -19213
rect 6513 -19323 6563 -19283
rect 6533 -19343 6563 -19323
rect 6623 -19323 6673 -19283
rect 6623 -19343 6653 -19323
rect 6733 -19383 6793 -19123
rect 6393 -19393 6473 -19383
rect 6393 -19453 6403 -19393
rect 6463 -19403 6473 -19393
rect 6713 -19393 6793 -19383
rect 6713 -19403 6723 -19393
rect 6463 -19453 6723 -19403
rect 6783 -19453 6793 -19393
rect 6393 -19463 6793 -19453
rect 6851 -19043 7251 -19033
rect 6851 -19103 6861 -19043
rect 6921 -19093 7181 -19043
rect 6921 -19103 6931 -19093
rect 6851 -19113 6931 -19103
rect 7171 -19103 7181 -19093
rect 7241 -19103 7251 -19043
rect 7171 -19113 7251 -19103
rect 6851 -19383 6911 -19113
rect 7181 -19123 7251 -19113
rect 6991 -19173 7021 -19153
rect 6971 -19213 7021 -19173
rect 7081 -19173 7111 -19153
rect 7081 -19213 7131 -19173
rect 6971 -19283 7131 -19213
rect 6971 -19323 7021 -19283
rect 6991 -19343 7021 -19323
rect 7081 -19323 7131 -19283
rect 7081 -19343 7111 -19323
rect 7191 -19383 7251 -19123
rect 6851 -19393 6931 -19383
rect 6851 -19453 6861 -19393
rect 6921 -19403 6931 -19393
rect 7171 -19393 7251 -19383
rect 7171 -19403 7181 -19393
rect 6921 -19453 7181 -19403
rect 7241 -19453 7251 -19393
rect 6851 -19463 7251 -19453
rect 7307 -19043 7707 -19033
rect 7307 -19103 7317 -19043
rect 7377 -19093 7637 -19043
rect 7377 -19103 7387 -19093
rect 7307 -19113 7387 -19103
rect 7627 -19103 7637 -19093
rect 7697 -19103 7707 -19043
rect 7627 -19113 7707 -19103
rect 7307 -19383 7367 -19113
rect 7637 -19123 7707 -19113
rect 7447 -19173 7477 -19153
rect 7427 -19213 7477 -19173
rect 7537 -19173 7567 -19153
rect 7537 -19213 7587 -19173
rect 7427 -19283 7587 -19213
rect 7427 -19323 7477 -19283
rect 7447 -19343 7477 -19323
rect 7537 -19323 7587 -19283
rect 7537 -19343 7567 -19323
rect 7647 -19383 7707 -19123
rect 7307 -19393 7387 -19383
rect 7307 -19453 7317 -19393
rect 7377 -19403 7387 -19393
rect 7627 -19393 7707 -19383
rect 7627 -19403 7637 -19393
rect 7377 -19453 7637 -19403
rect 7697 -19453 7707 -19393
rect 7307 -19463 7707 -19453
rect 7763 -19043 8163 -19033
rect 7763 -19103 7773 -19043
rect 7833 -19093 8093 -19043
rect 7833 -19103 7843 -19093
rect 7763 -19113 7843 -19103
rect 8083 -19103 8093 -19093
rect 8153 -19103 8163 -19043
rect 8083 -19113 8163 -19103
rect 7763 -19383 7823 -19113
rect 8093 -19123 8163 -19113
rect 7903 -19173 7933 -19153
rect 7883 -19213 7933 -19173
rect 7993 -19173 8023 -19153
rect 7993 -19213 8043 -19173
rect 7883 -19283 8043 -19213
rect 7883 -19323 7933 -19283
rect 7903 -19343 7933 -19323
rect 7993 -19323 8043 -19283
rect 7993 -19343 8023 -19323
rect 8103 -19383 8163 -19123
rect 7763 -19393 7843 -19383
rect 7763 -19453 7773 -19393
rect 7833 -19403 7843 -19393
rect 8083 -19393 8163 -19383
rect 8083 -19403 8093 -19393
rect 7833 -19453 8093 -19403
rect 8153 -19453 8163 -19393
rect 7763 -19463 8163 -19453
rect 8237 -19043 8637 -19033
rect 8237 -19103 8247 -19043
rect 8307 -19093 8567 -19043
rect 8307 -19103 8317 -19093
rect 8237 -19113 8317 -19103
rect 8557 -19103 8567 -19093
rect 8627 -19103 8637 -19043
rect 8557 -19113 8637 -19103
rect 8237 -19383 8297 -19113
rect 8567 -19123 8637 -19113
rect 8377 -19173 8407 -19153
rect 8357 -19213 8407 -19173
rect 8467 -19173 8497 -19153
rect 8467 -19213 8517 -19173
rect 8357 -19283 8517 -19213
rect 8357 -19323 8407 -19283
rect 8377 -19343 8407 -19323
rect 8467 -19323 8517 -19283
rect 8467 -19343 8497 -19323
rect 8577 -19383 8637 -19123
rect 8237 -19393 8317 -19383
rect 8237 -19453 8247 -19393
rect 8307 -19403 8317 -19393
rect 8557 -19393 8637 -19383
rect 8557 -19403 8567 -19393
rect 8307 -19453 8567 -19403
rect 8627 -19453 8637 -19393
rect 8237 -19463 8637 -19453
rect 8693 -19043 9093 -19033
rect 8693 -19103 8703 -19043
rect 8763 -19093 9023 -19043
rect 8763 -19103 8773 -19093
rect 8693 -19113 8773 -19103
rect 9013 -19103 9023 -19093
rect 9083 -19103 9093 -19043
rect 9013 -19113 9093 -19103
rect 8693 -19383 8753 -19113
rect 9023 -19123 9093 -19113
rect 8833 -19173 8863 -19153
rect 8813 -19213 8863 -19173
rect 8923 -19173 8953 -19153
rect 8923 -19213 8973 -19173
rect 8813 -19283 8973 -19213
rect 8813 -19323 8863 -19283
rect 8833 -19343 8863 -19323
rect 8923 -19323 8973 -19283
rect 8923 -19343 8953 -19323
rect 9033 -19383 9093 -19123
rect 8693 -19393 8773 -19383
rect 8693 -19453 8703 -19393
rect 8763 -19403 8773 -19393
rect 9013 -19393 9093 -19383
rect 9013 -19403 9023 -19393
rect 8763 -19453 9023 -19403
rect 9083 -19453 9093 -19393
rect 8693 -19463 9093 -19453
rect 9151 -19043 9551 -19033
rect 9151 -19103 9161 -19043
rect 9221 -19093 9481 -19043
rect 9221 -19103 9231 -19093
rect 9151 -19113 9231 -19103
rect 9471 -19103 9481 -19093
rect 9541 -19103 9551 -19043
rect 9471 -19113 9551 -19103
rect 9151 -19383 9211 -19113
rect 9481 -19123 9551 -19113
rect 9291 -19173 9321 -19153
rect 9271 -19213 9321 -19173
rect 9381 -19173 9411 -19153
rect 9381 -19213 9431 -19173
rect 9271 -19283 9431 -19213
rect 9271 -19323 9321 -19283
rect 9291 -19343 9321 -19323
rect 9381 -19323 9431 -19283
rect 9381 -19343 9411 -19323
rect 9491 -19383 9551 -19123
rect 9151 -19393 9231 -19383
rect 9151 -19453 9161 -19393
rect 9221 -19403 9231 -19393
rect 9471 -19393 9551 -19383
rect 9471 -19403 9481 -19393
rect 9221 -19453 9481 -19403
rect 9541 -19453 9551 -19393
rect 9151 -19463 9551 -19453
rect 9607 -19043 10007 -19033
rect 9607 -19103 9617 -19043
rect 9677 -19093 9937 -19043
rect 9677 -19103 9687 -19093
rect 9607 -19113 9687 -19103
rect 9927 -19103 9937 -19093
rect 9997 -19103 10007 -19043
rect 9927 -19113 10007 -19103
rect 9607 -19383 9667 -19113
rect 9937 -19123 10007 -19113
rect 9747 -19173 9777 -19153
rect 9727 -19213 9777 -19173
rect 9837 -19173 9867 -19153
rect 9837 -19213 9887 -19173
rect 9727 -19283 9887 -19213
rect 9727 -19323 9777 -19283
rect 9747 -19343 9777 -19323
rect 9837 -19323 9887 -19283
rect 9837 -19343 9867 -19323
rect 9947 -19383 10007 -19123
rect 9607 -19393 9687 -19383
rect 9607 -19453 9617 -19393
rect 9677 -19403 9687 -19393
rect 9927 -19393 10007 -19383
rect 9927 -19403 9937 -19393
rect 9677 -19453 9937 -19403
rect 9997 -19453 10007 -19393
rect 9607 -19463 10007 -19453
rect 10063 -19043 10463 -19033
rect 10063 -19103 10073 -19043
rect 10133 -19093 10393 -19043
rect 10133 -19103 10143 -19093
rect 10063 -19113 10143 -19103
rect 10383 -19103 10393 -19093
rect 10453 -19103 10463 -19043
rect 10383 -19113 10463 -19103
rect 10063 -19383 10123 -19113
rect 10393 -19123 10463 -19113
rect 10203 -19173 10233 -19153
rect 10183 -19213 10233 -19173
rect 10293 -19173 10323 -19153
rect 10293 -19213 10343 -19173
rect 10183 -19283 10343 -19213
rect 10183 -19323 10233 -19283
rect 10203 -19343 10233 -19323
rect 10293 -19323 10343 -19283
rect 10293 -19343 10323 -19323
rect 10403 -19383 10463 -19123
rect 10063 -19393 10143 -19383
rect 10063 -19453 10073 -19393
rect 10133 -19403 10143 -19393
rect 10383 -19393 10463 -19383
rect 10383 -19403 10393 -19393
rect 10133 -19453 10393 -19403
rect 10453 -19453 10463 -19393
rect 10063 -19463 10463 -19453
rect 10521 -19043 10921 -19033
rect 10521 -19103 10531 -19043
rect 10591 -19093 10851 -19043
rect 10591 -19103 10601 -19093
rect 10521 -19113 10601 -19103
rect 10841 -19103 10851 -19093
rect 10911 -19103 10921 -19043
rect 10841 -19113 10921 -19103
rect 10521 -19383 10581 -19113
rect 10851 -19123 10921 -19113
rect 10661 -19173 10691 -19153
rect 10641 -19213 10691 -19173
rect 10751 -19173 10781 -19153
rect 10751 -19213 10801 -19173
rect 10641 -19283 10801 -19213
rect 10641 -19323 10691 -19283
rect 10661 -19343 10691 -19323
rect 10751 -19323 10801 -19283
rect 10751 -19343 10781 -19323
rect 10861 -19383 10921 -19123
rect 10521 -19393 10601 -19383
rect 10521 -19453 10531 -19393
rect 10591 -19403 10601 -19393
rect 10841 -19393 10921 -19383
rect 10841 -19403 10851 -19393
rect 10591 -19453 10851 -19403
rect 10911 -19453 10921 -19393
rect 10521 -19463 10921 -19453
rect 10977 -19043 11377 -19033
rect 10977 -19103 10987 -19043
rect 11047 -19093 11307 -19043
rect 11047 -19103 11057 -19093
rect 10977 -19113 11057 -19103
rect 11297 -19103 11307 -19093
rect 11367 -19103 11377 -19043
rect 11297 -19113 11377 -19103
rect 10977 -19383 11037 -19113
rect 11307 -19123 11377 -19113
rect 11117 -19173 11147 -19153
rect 11097 -19213 11147 -19173
rect 11207 -19173 11237 -19153
rect 11207 -19213 11257 -19173
rect 11097 -19283 11257 -19213
rect 11097 -19323 11147 -19283
rect 11117 -19343 11147 -19323
rect 11207 -19323 11257 -19283
rect 11207 -19343 11237 -19323
rect 11317 -19383 11377 -19123
rect 10977 -19393 11057 -19383
rect 10977 -19453 10987 -19393
rect 11047 -19403 11057 -19393
rect 11297 -19393 11377 -19383
rect 11297 -19403 11307 -19393
rect 11047 -19453 11307 -19403
rect 11367 -19453 11377 -19393
rect 10977 -19463 11377 -19453
rect 11433 -19043 11833 -19033
rect 11433 -19103 11443 -19043
rect 11503 -19093 11763 -19043
rect 11503 -19103 11513 -19093
rect 11433 -19113 11513 -19103
rect 11753 -19103 11763 -19093
rect 11823 -19103 11833 -19043
rect 11753 -19113 11833 -19103
rect 11433 -19383 11493 -19113
rect 11763 -19123 11833 -19113
rect 11573 -19173 11603 -19153
rect 11553 -19213 11603 -19173
rect 11663 -19173 11693 -19153
rect 11663 -19213 11713 -19173
rect 11553 -19283 11713 -19213
rect 11553 -19323 11603 -19283
rect 11573 -19343 11603 -19323
rect 11663 -19323 11713 -19283
rect 11663 -19343 11693 -19323
rect 11773 -19383 11833 -19123
rect 11433 -19393 11513 -19383
rect 11433 -19453 11443 -19393
rect 11503 -19403 11513 -19393
rect 11753 -19393 11833 -19383
rect 11753 -19403 11763 -19393
rect 11503 -19453 11763 -19403
rect 11823 -19453 11833 -19393
rect 11433 -19463 11833 -19453
rect 11891 -19043 12291 -19033
rect 11891 -19103 11901 -19043
rect 11961 -19093 12221 -19043
rect 11961 -19103 11971 -19093
rect 11891 -19113 11971 -19103
rect 12211 -19103 12221 -19093
rect 12281 -19103 12291 -19043
rect 12211 -19113 12291 -19103
rect 11891 -19383 11951 -19113
rect 12221 -19123 12291 -19113
rect 12031 -19173 12061 -19153
rect 12011 -19213 12061 -19173
rect 12121 -19173 12151 -19153
rect 12121 -19213 12171 -19173
rect 12011 -19283 12171 -19213
rect 12011 -19323 12061 -19283
rect 12031 -19343 12061 -19323
rect 12121 -19323 12171 -19283
rect 12121 -19343 12151 -19323
rect 12231 -19383 12291 -19123
rect 11891 -19393 11971 -19383
rect 11891 -19453 11901 -19393
rect 11961 -19403 11971 -19393
rect 12211 -19393 12291 -19383
rect 12211 -19403 12221 -19393
rect 11961 -19453 12221 -19403
rect 12281 -19453 12291 -19393
rect 11891 -19463 12291 -19453
rect 12347 -19043 12747 -19033
rect 12347 -19103 12357 -19043
rect 12417 -19093 12677 -19043
rect 12417 -19103 12427 -19093
rect 12347 -19113 12427 -19103
rect 12667 -19103 12677 -19093
rect 12737 -19103 12747 -19043
rect 12667 -19113 12747 -19103
rect 12347 -19383 12407 -19113
rect 12677 -19123 12747 -19113
rect 12487 -19173 12517 -19153
rect 12467 -19213 12517 -19173
rect 12577 -19173 12607 -19153
rect 12577 -19213 12627 -19173
rect 12467 -19283 12627 -19213
rect 12467 -19323 12517 -19283
rect 12487 -19343 12517 -19323
rect 12577 -19323 12627 -19283
rect 12577 -19343 12607 -19323
rect 12687 -19383 12747 -19123
rect 12347 -19393 12427 -19383
rect 12347 -19453 12357 -19393
rect 12417 -19403 12427 -19393
rect 12667 -19393 12747 -19383
rect 12667 -19403 12677 -19393
rect 12417 -19453 12677 -19403
rect 12737 -19453 12747 -19393
rect 12347 -19463 12747 -19453
rect 12803 -19043 13203 -19033
rect 12803 -19103 12813 -19043
rect 12873 -19093 13133 -19043
rect 12873 -19103 12883 -19093
rect 12803 -19113 12883 -19103
rect 13123 -19103 13133 -19093
rect 13193 -19103 13203 -19043
rect 13123 -19113 13203 -19103
rect 12803 -19383 12863 -19113
rect 13133 -19123 13203 -19113
rect 12943 -19173 12973 -19153
rect 12923 -19213 12973 -19173
rect 13033 -19173 13063 -19153
rect 13033 -19213 13083 -19173
rect 12923 -19283 13083 -19213
rect 12923 -19323 12973 -19283
rect 12943 -19343 12973 -19323
rect 13033 -19323 13083 -19283
rect 13033 -19343 13063 -19323
rect 13143 -19383 13203 -19123
rect 12803 -19393 12883 -19383
rect 12803 -19453 12813 -19393
rect 12873 -19403 12883 -19393
rect 13123 -19393 13203 -19383
rect 13123 -19403 13133 -19393
rect 12873 -19453 13133 -19403
rect 13193 -19453 13203 -19393
rect 12803 -19463 13203 -19453
rect 13261 -19043 13661 -19033
rect 13261 -19103 13271 -19043
rect 13331 -19093 13591 -19043
rect 13331 -19103 13341 -19093
rect 13261 -19113 13341 -19103
rect 13581 -19103 13591 -19093
rect 13651 -19103 13661 -19043
rect 13581 -19113 13661 -19103
rect 13261 -19383 13321 -19113
rect 13591 -19123 13661 -19113
rect 13401 -19173 13431 -19153
rect 13381 -19213 13431 -19173
rect 13491 -19173 13521 -19153
rect 13491 -19213 13541 -19173
rect 13381 -19283 13541 -19213
rect 13381 -19323 13431 -19283
rect 13401 -19343 13431 -19323
rect 13491 -19323 13541 -19283
rect 13491 -19343 13521 -19323
rect 13601 -19383 13661 -19123
rect 13261 -19393 13341 -19383
rect 13261 -19453 13271 -19393
rect 13331 -19403 13341 -19393
rect 13581 -19393 13661 -19383
rect 13581 -19403 13591 -19393
rect 13331 -19453 13591 -19403
rect 13651 -19453 13661 -19393
rect 13261 -19463 13661 -19453
rect 13717 -19043 14117 -19033
rect 13717 -19103 13727 -19043
rect 13787 -19093 14047 -19043
rect 13787 -19103 13797 -19093
rect 13717 -19113 13797 -19103
rect 14037 -19103 14047 -19093
rect 14107 -19103 14117 -19043
rect 14037 -19113 14117 -19103
rect 13717 -19383 13777 -19113
rect 14047 -19123 14117 -19113
rect 13857 -19173 13887 -19153
rect 13837 -19213 13887 -19173
rect 13947 -19173 13977 -19153
rect 13947 -19213 13997 -19173
rect 13837 -19283 13997 -19213
rect 13837 -19323 13887 -19283
rect 13857 -19343 13887 -19323
rect 13947 -19323 13997 -19283
rect 13947 -19343 13977 -19323
rect 14057 -19383 14117 -19123
rect 13717 -19393 13797 -19383
rect 13717 -19453 13727 -19393
rect 13787 -19403 13797 -19393
rect 14037 -19393 14117 -19383
rect 14037 -19403 14047 -19393
rect 13787 -19453 14047 -19403
rect 14107 -19453 14117 -19393
rect 13717 -19463 14117 -19453
rect 14173 -19043 14573 -19033
rect 14173 -19103 14183 -19043
rect 14243 -19093 14503 -19043
rect 14243 -19103 14253 -19093
rect 14173 -19113 14253 -19103
rect 14493 -19103 14503 -19093
rect 14563 -19103 14573 -19043
rect 14493 -19113 14573 -19103
rect 14173 -19383 14233 -19113
rect 14503 -19123 14573 -19113
rect 14313 -19173 14343 -19153
rect 14293 -19213 14343 -19173
rect 14403 -19173 14433 -19153
rect 14403 -19213 14453 -19173
rect 14293 -19283 14453 -19213
rect 14293 -19323 14343 -19283
rect 14313 -19343 14343 -19323
rect 14403 -19323 14453 -19283
rect 14403 -19343 14433 -19323
rect 14513 -19383 14573 -19123
rect 14173 -19393 14253 -19383
rect 14173 -19453 14183 -19393
rect 14243 -19403 14253 -19393
rect 14493 -19393 14573 -19383
rect 14493 -19403 14503 -19393
rect 14243 -19453 14503 -19403
rect 14563 -19453 14573 -19393
rect 14173 -19463 14573 -19453
rect 14631 -19043 15031 -19033
rect 14631 -19103 14641 -19043
rect 14701 -19093 14961 -19043
rect 14701 -19103 14711 -19093
rect 14631 -19113 14711 -19103
rect 14951 -19103 14961 -19093
rect 15021 -19103 15031 -19043
rect 14951 -19113 15031 -19103
rect 14631 -19383 14691 -19113
rect 14961 -19123 15031 -19113
rect 14771 -19173 14801 -19153
rect 14751 -19213 14801 -19173
rect 14861 -19173 14891 -19153
rect 14861 -19213 14911 -19173
rect 14751 -19283 14911 -19213
rect 14751 -19323 14801 -19283
rect 14771 -19343 14801 -19323
rect 14861 -19323 14911 -19283
rect 14861 -19343 14891 -19323
rect 14971 -19383 15031 -19123
rect 14631 -19393 14711 -19383
rect 14631 -19453 14641 -19393
rect 14701 -19403 14711 -19393
rect 14951 -19393 15031 -19383
rect 14951 -19403 14961 -19393
rect 14701 -19453 14961 -19403
rect 15021 -19453 15031 -19393
rect 14631 -19463 15031 -19453
rect 15087 -19043 15487 -19033
rect 15087 -19103 15097 -19043
rect 15157 -19093 15417 -19043
rect 15157 -19103 15167 -19093
rect 15087 -19113 15167 -19103
rect 15407 -19103 15417 -19093
rect 15477 -19103 15487 -19043
rect 15407 -19113 15487 -19103
rect 15087 -19383 15147 -19113
rect 15417 -19123 15487 -19113
rect 15227 -19173 15257 -19153
rect 15207 -19213 15257 -19173
rect 15317 -19173 15347 -19153
rect 15317 -19213 15367 -19173
rect 15207 -19283 15367 -19213
rect 15207 -19323 15257 -19283
rect 15227 -19343 15257 -19323
rect 15317 -19323 15367 -19283
rect 15317 -19343 15347 -19323
rect 15427 -19383 15487 -19123
rect 15087 -19393 15167 -19383
rect 15087 -19453 15097 -19393
rect 15157 -19403 15167 -19393
rect 15407 -19393 15487 -19383
rect 15407 -19403 15417 -19393
rect 15157 -19453 15417 -19403
rect 15477 -19453 15487 -19393
rect 15087 -19463 15487 -19453
rect 1 -19537 401 -19527
rect 1 -19597 11 -19537
rect 71 -19587 331 -19537
rect 71 -19597 81 -19587
rect 1 -19607 81 -19597
rect 321 -19597 331 -19587
rect 391 -19597 401 -19537
rect 321 -19607 401 -19597
rect 1 -19877 61 -19607
rect 331 -19617 401 -19607
rect 141 -19667 171 -19647
rect 121 -19707 171 -19667
rect 231 -19667 261 -19647
rect 231 -19707 281 -19667
rect 121 -19777 281 -19707
rect 121 -19817 171 -19777
rect 141 -19837 171 -19817
rect 231 -19817 281 -19777
rect 231 -19837 261 -19817
rect 341 -19877 401 -19617
rect 1 -19887 81 -19877
rect 1 -19947 11 -19887
rect 71 -19897 81 -19887
rect 321 -19887 401 -19877
rect 321 -19897 331 -19887
rect 71 -19947 331 -19897
rect 391 -19947 401 -19887
rect 1 -19957 401 -19947
rect 457 -19537 857 -19527
rect 457 -19597 467 -19537
rect 527 -19587 787 -19537
rect 527 -19597 537 -19587
rect 457 -19607 537 -19597
rect 777 -19597 787 -19587
rect 847 -19597 857 -19537
rect 777 -19607 857 -19597
rect 457 -19877 517 -19607
rect 787 -19617 857 -19607
rect 597 -19667 627 -19647
rect 577 -19707 627 -19667
rect 687 -19667 717 -19647
rect 687 -19707 737 -19667
rect 577 -19777 737 -19707
rect 577 -19817 627 -19777
rect 597 -19837 627 -19817
rect 687 -19817 737 -19777
rect 687 -19837 717 -19817
rect 797 -19877 857 -19617
rect 457 -19887 537 -19877
rect 457 -19947 467 -19887
rect 527 -19897 537 -19887
rect 777 -19887 857 -19877
rect 777 -19897 787 -19887
rect 527 -19947 787 -19897
rect 847 -19947 857 -19887
rect 457 -19957 857 -19947
rect 913 -19537 1313 -19527
rect 913 -19597 923 -19537
rect 983 -19587 1243 -19537
rect 983 -19597 993 -19587
rect 913 -19607 993 -19597
rect 1233 -19597 1243 -19587
rect 1303 -19597 1313 -19537
rect 1233 -19607 1313 -19597
rect 913 -19877 973 -19607
rect 1243 -19617 1313 -19607
rect 1053 -19667 1083 -19647
rect 1033 -19707 1083 -19667
rect 1143 -19667 1173 -19647
rect 1143 -19707 1193 -19667
rect 1033 -19777 1193 -19707
rect 1033 -19817 1083 -19777
rect 1053 -19837 1083 -19817
rect 1143 -19817 1193 -19777
rect 1143 -19837 1173 -19817
rect 1253 -19877 1313 -19617
rect 913 -19887 993 -19877
rect 913 -19947 923 -19887
rect 983 -19897 993 -19887
rect 1233 -19887 1313 -19877
rect 1233 -19897 1243 -19887
rect 983 -19947 1243 -19897
rect 1303 -19947 1313 -19887
rect 913 -19957 1313 -19947
rect 1371 -19537 1771 -19527
rect 1371 -19597 1381 -19537
rect 1441 -19587 1701 -19537
rect 1441 -19597 1451 -19587
rect 1371 -19607 1451 -19597
rect 1691 -19597 1701 -19587
rect 1761 -19597 1771 -19537
rect 1691 -19607 1771 -19597
rect 1371 -19877 1431 -19607
rect 1701 -19617 1771 -19607
rect 1511 -19667 1541 -19647
rect 1491 -19707 1541 -19667
rect 1601 -19667 1631 -19647
rect 1601 -19707 1651 -19667
rect 1491 -19777 1651 -19707
rect 1491 -19817 1541 -19777
rect 1511 -19837 1541 -19817
rect 1601 -19817 1651 -19777
rect 1601 -19837 1631 -19817
rect 1711 -19877 1771 -19617
rect 1371 -19887 1451 -19877
rect 1371 -19947 1381 -19887
rect 1441 -19897 1451 -19887
rect 1691 -19887 1771 -19877
rect 1691 -19897 1701 -19887
rect 1441 -19947 1701 -19897
rect 1761 -19947 1771 -19887
rect 1371 -19957 1771 -19947
rect 1827 -19537 2227 -19527
rect 1827 -19597 1837 -19537
rect 1897 -19587 2157 -19537
rect 1897 -19597 1907 -19587
rect 1827 -19607 1907 -19597
rect 2147 -19597 2157 -19587
rect 2217 -19597 2227 -19537
rect 2147 -19607 2227 -19597
rect 1827 -19877 1887 -19607
rect 2157 -19617 2227 -19607
rect 1967 -19667 1997 -19647
rect 1947 -19707 1997 -19667
rect 2057 -19667 2087 -19647
rect 2057 -19707 2107 -19667
rect 1947 -19777 2107 -19707
rect 1947 -19817 1997 -19777
rect 1967 -19837 1997 -19817
rect 2057 -19817 2107 -19777
rect 2057 -19837 2087 -19817
rect 2167 -19877 2227 -19617
rect 1827 -19887 1907 -19877
rect 1827 -19947 1837 -19887
rect 1897 -19897 1907 -19887
rect 2147 -19887 2227 -19877
rect 2147 -19897 2157 -19887
rect 1897 -19947 2157 -19897
rect 2217 -19947 2227 -19887
rect 1827 -19957 2227 -19947
rect 2283 -19537 2683 -19527
rect 2283 -19597 2293 -19537
rect 2353 -19587 2613 -19537
rect 2353 -19597 2363 -19587
rect 2283 -19607 2363 -19597
rect 2603 -19597 2613 -19587
rect 2673 -19597 2683 -19537
rect 2603 -19607 2683 -19597
rect 2283 -19877 2343 -19607
rect 2613 -19617 2683 -19607
rect 2423 -19667 2453 -19647
rect 2403 -19707 2453 -19667
rect 2513 -19667 2543 -19647
rect 2513 -19707 2563 -19667
rect 2403 -19777 2563 -19707
rect 2403 -19817 2453 -19777
rect 2423 -19837 2453 -19817
rect 2513 -19817 2563 -19777
rect 2513 -19837 2543 -19817
rect 2623 -19877 2683 -19617
rect 2283 -19887 2363 -19877
rect 2283 -19947 2293 -19887
rect 2353 -19897 2363 -19887
rect 2603 -19887 2683 -19877
rect 2603 -19897 2613 -19887
rect 2353 -19947 2613 -19897
rect 2673 -19947 2683 -19887
rect 2283 -19957 2683 -19947
rect 2741 -19537 3141 -19527
rect 2741 -19597 2751 -19537
rect 2811 -19587 3071 -19537
rect 2811 -19597 2821 -19587
rect 2741 -19607 2821 -19597
rect 3061 -19597 3071 -19587
rect 3131 -19597 3141 -19537
rect 3061 -19607 3141 -19597
rect 2741 -19877 2801 -19607
rect 3071 -19617 3141 -19607
rect 2881 -19667 2911 -19647
rect 2861 -19707 2911 -19667
rect 2971 -19667 3001 -19647
rect 2971 -19707 3021 -19667
rect 2861 -19777 3021 -19707
rect 2861 -19817 2911 -19777
rect 2881 -19837 2911 -19817
rect 2971 -19817 3021 -19777
rect 2971 -19837 3001 -19817
rect 3081 -19877 3141 -19617
rect 2741 -19887 2821 -19877
rect 2741 -19947 2751 -19887
rect 2811 -19897 2821 -19887
rect 3061 -19887 3141 -19877
rect 3061 -19897 3071 -19887
rect 2811 -19947 3071 -19897
rect 3131 -19947 3141 -19887
rect 2741 -19957 3141 -19947
rect 3197 -19537 3597 -19527
rect 3197 -19597 3207 -19537
rect 3267 -19587 3527 -19537
rect 3267 -19597 3277 -19587
rect 3197 -19607 3277 -19597
rect 3517 -19597 3527 -19587
rect 3587 -19597 3597 -19537
rect 3517 -19607 3597 -19597
rect 3197 -19877 3257 -19607
rect 3527 -19617 3597 -19607
rect 3337 -19667 3367 -19647
rect 3317 -19707 3367 -19667
rect 3427 -19667 3457 -19647
rect 3427 -19707 3477 -19667
rect 3317 -19777 3477 -19707
rect 3317 -19817 3367 -19777
rect 3337 -19837 3367 -19817
rect 3427 -19817 3477 -19777
rect 3427 -19837 3457 -19817
rect 3537 -19877 3597 -19617
rect 3197 -19887 3277 -19877
rect 3197 -19947 3207 -19887
rect 3267 -19897 3277 -19887
rect 3517 -19887 3597 -19877
rect 3517 -19897 3527 -19887
rect 3267 -19947 3527 -19897
rect 3587 -19947 3597 -19887
rect 3197 -19957 3597 -19947
rect 3653 -19537 4053 -19527
rect 3653 -19597 3663 -19537
rect 3723 -19587 3983 -19537
rect 3723 -19597 3733 -19587
rect 3653 -19607 3733 -19597
rect 3973 -19597 3983 -19587
rect 4043 -19597 4053 -19537
rect 3973 -19607 4053 -19597
rect 3653 -19877 3713 -19607
rect 3983 -19617 4053 -19607
rect 3793 -19667 3823 -19647
rect 3773 -19707 3823 -19667
rect 3883 -19667 3913 -19647
rect 3883 -19707 3933 -19667
rect 3773 -19777 3933 -19707
rect 3773 -19817 3823 -19777
rect 3793 -19837 3823 -19817
rect 3883 -19817 3933 -19777
rect 3883 -19837 3913 -19817
rect 3993 -19877 4053 -19617
rect 3653 -19887 3733 -19877
rect 3653 -19947 3663 -19887
rect 3723 -19897 3733 -19887
rect 3973 -19887 4053 -19877
rect 3973 -19897 3983 -19887
rect 3723 -19947 3983 -19897
rect 4043 -19947 4053 -19887
rect 3653 -19957 4053 -19947
rect 4111 -19537 4511 -19527
rect 4111 -19597 4121 -19537
rect 4181 -19587 4441 -19537
rect 4181 -19597 4191 -19587
rect 4111 -19607 4191 -19597
rect 4431 -19597 4441 -19587
rect 4501 -19597 4511 -19537
rect 4431 -19607 4511 -19597
rect 4111 -19877 4171 -19607
rect 4441 -19617 4511 -19607
rect 4251 -19667 4281 -19647
rect 4231 -19707 4281 -19667
rect 4341 -19667 4371 -19647
rect 4341 -19707 4391 -19667
rect 4231 -19777 4391 -19707
rect 4231 -19817 4281 -19777
rect 4251 -19837 4281 -19817
rect 4341 -19817 4391 -19777
rect 4341 -19837 4371 -19817
rect 4451 -19877 4511 -19617
rect 4111 -19887 4191 -19877
rect 4111 -19947 4121 -19887
rect 4181 -19897 4191 -19887
rect 4431 -19887 4511 -19877
rect 4431 -19897 4441 -19887
rect 4181 -19947 4441 -19897
rect 4501 -19947 4511 -19887
rect 4111 -19957 4511 -19947
rect 4567 -19537 4967 -19527
rect 4567 -19597 4577 -19537
rect 4637 -19587 4897 -19537
rect 4637 -19597 4647 -19587
rect 4567 -19607 4647 -19597
rect 4887 -19597 4897 -19587
rect 4957 -19597 4967 -19537
rect 4887 -19607 4967 -19597
rect 4567 -19877 4627 -19607
rect 4897 -19617 4967 -19607
rect 4707 -19667 4737 -19647
rect 4687 -19707 4737 -19667
rect 4797 -19667 4827 -19647
rect 4797 -19707 4847 -19667
rect 4687 -19777 4847 -19707
rect 4687 -19817 4737 -19777
rect 4707 -19837 4737 -19817
rect 4797 -19817 4847 -19777
rect 4797 -19837 4827 -19817
rect 4907 -19877 4967 -19617
rect 4567 -19887 4647 -19877
rect 4567 -19947 4577 -19887
rect 4637 -19897 4647 -19887
rect 4887 -19887 4967 -19877
rect 4887 -19897 4897 -19887
rect 4637 -19947 4897 -19897
rect 4957 -19947 4967 -19887
rect 4567 -19957 4967 -19947
rect 5023 -19537 5423 -19527
rect 5023 -19597 5033 -19537
rect 5093 -19587 5353 -19537
rect 5093 -19597 5103 -19587
rect 5023 -19607 5103 -19597
rect 5343 -19597 5353 -19587
rect 5413 -19597 5423 -19537
rect 5343 -19607 5423 -19597
rect 5023 -19877 5083 -19607
rect 5353 -19617 5423 -19607
rect 5163 -19667 5193 -19647
rect 5143 -19707 5193 -19667
rect 5253 -19667 5283 -19647
rect 5253 -19707 5303 -19667
rect 5143 -19777 5303 -19707
rect 5143 -19817 5193 -19777
rect 5163 -19837 5193 -19817
rect 5253 -19817 5303 -19777
rect 5253 -19837 5283 -19817
rect 5363 -19877 5423 -19617
rect 5023 -19887 5103 -19877
rect 5023 -19947 5033 -19887
rect 5093 -19897 5103 -19887
rect 5343 -19887 5423 -19877
rect 5343 -19897 5353 -19887
rect 5093 -19947 5353 -19897
rect 5413 -19947 5423 -19887
rect 5023 -19957 5423 -19947
rect 5481 -19537 5881 -19527
rect 5481 -19597 5491 -19537
rect 5551 -19587 5811 -19537
rect 5551 -19597 5561 -19587
rect 5481 -19607 5561 -19597
rect 5801 -19597 5811 -19587
rect 5871 -19597 5881 -19537
rect 5801 -19607 5881 -19597
rect 5481 -19877 5541 -19607
rect 5811 -19617 5881 -19607
rect 5621 -19667 5651 -19647
rect 5601 -19707 5651 -19667
rect 5711 -19667 5741 -19647
rect 5711 -19707 5761 -19667
rect 5601 -19777 5761 -19707
rect 5601 -19817 5651 -19777
rect 5621 -19837 5651 -19817
rect 5711 -19817 5761 -19777
rect 5711 -19837 5741 -19817
rect 5821 -19877 5881 -19617
rect 5481 -19887 5561 -19877
rect 5481 -19947 5491 -19887
rect 5551 -19897 5561 -19887
rect 5801 -19887 5881 -19877
rect 5801 -19897 5811 -19887
rect 5551 -19947 5811 -19897
rect 5871 -19947 5881 -19887
rect 5481 -19957 5881 -19947
rect 5937 -19537 6337 -19527
rect 5937 -19597 5947 -19537
rect 6007 -19587 6267 -19537
rect 6007 -19597 6017 -19587
rect 5937 -19607 6017 -19597
rect 6257 -19597 6267 -19587
rect 6327 -19597 6337 -19537
rect 6257 -19607 6337 -19597
rect 5937 -19877 5997 -19607
rect 6267 -19617 6337 -19607
rect 6077 -19667 6107 -19647
rect 6057 -19707 6107 -19667
rect 6167 -19667 6197 -19647
rect 6167 -19707 6217 -19667
rect 6057 -19777 6217 -19707
rect 6057 -19817 6107 -19777
rect 6077 -19837 6107 -19817
rect 6167 -19817 6217 -19777
rect 6167 -19837 6197 -19817
rect 6277 -19877 6337 -19617
rect 5937 -19887 6017 -19877
rect 5937 -19947 5947 -19887
rect 6007 -19897 6017 -19887
rect 6257 -19887 6337 -19877
rect 6257 -19897 6267 -19887
rect 6007 -19947 6267 -19897
rect 6327 -19947 6337 -19887
rect 5937 -19957 6337 -19947
rect 6393 -19537 6793 -19527
rect 6393 -19597 6403 -19537
rect 6463 -19587 6723 -19537
rect 6463 -19597 6473 -19587
rect 6393 -19607 6473 -19597
rect 6713 -19597 6723 -19587
rect 6783 -19597 6793 -19537
rect 6713 -19607 6793 -19597
rect 6393 -19877 6453 -19607
rect 6723 -19617 6793 -19607
rect 6533 -19667 6563 -19647
rect 6513 -19707 6563 -19667
rect 6623 -19667 6653 -19647
rect 6623 -19707 6673 -19667
rect 6513 -19777 6673 -19707
rect 6513 -19817 6563 -19777
rect 6533 -19837 6563 -19817
rect 6623 -19817 6673 -19777
rect 6623 -19837 6653 -19817
rect 6733 -19877 6793 -19617
rect 6393 -19887 6473 -19877
rect 6393 -19947 6403 -19887
rect 6463 -19897 6473 -19887
rect 6713 -19887 6793 -19877
rect 6713 -19897 6723 -19887
rect 6463 -19947 6723 -19897
rect 6783 -19947 6793 -19887
rect 6393 -19957 6793 -19947
rect 6851 -19537 7251 -19527
rect 6851 -19597 6861 -19537
rect 6921 -19587 7181 -19537
rect 6921 -19597 6931 -19587
rect 6851 -19607 6931 -19597
rect 7171 -19597 7181 -19587
rect 7241 -19597 7251 -19537
rect 7171 -19607 7251 -19597
rect 6851 -19877 6911 -19607
rect 7181 -19617 7251 -19607
rect 6991 -19667 7021 -19647
rect 6971 -19707 7021 -19667
rect 7081 -19667 7111 -19647
rect 7081 -19707 7131 -19667
rect 6971 -19777 7131 -19707
rect 6971 -19817 7021 -19777
rect 6991 -19837 7021 -19817
rect 7081 -19817 7131 -19777
rect 7081 -19837 7111 -19817
rect 7191 -19877 7251 -19617
rect 6851 -19887 6931 -19877
rect 6851 -19947 6861 -19887
rect 6921 -19897 6931 -19887
rect 7171 -19887 7251 -19877
rect 7171 -19897 7181 -19887
rect 6921 -19947 7181 -19897
rect 7241 -19947 7251 -19887
rect 6851 -19957 7251 -19947
rect 7307 -19537 7707 -19527
rect 7307 -19597 7317 -19537
rect 7377 -19587 7637 -19537
rect 7377 -19597 7387 -19587
rect 7307 -19607 7387 -19597
rect 7627 -19597 7637 -19587
rect 7697 -19597 7707 -19537
rect 7627 -19607 7707 -19597
rect 7307 -19877 7367 -19607
rect 7637 -19617 7707 -19607
rect 7447 -19667 7477 -19647
rect 7427 -19707 7477 -19667
rect 7537 -19667 7567 -19647
rect 7537 -19707 7587 -19667
rect 7427 -19777 7587 -19707
rect 7427 -19817 7477 -19777
rect 7447 -19837 7477 -19817
rect 7537 -19817 7587 -19777
rect 7537 -19837 7567 -19817
rect 7647 -19877 7707 -19617
rect 7307 -19887 7387 -19877
rect 7307 -19947 7317 -19887
rect 7377 -19897 7387 -19887
rect 7627 -19887 7707 -19877
rect 7627 -19897 7637 -19887
rect 7377 -19947 7637 -19897
rect 7697 -19947 7707 -19887
rect 7307 -19957 7707 -19947
rect 7763 -19537 8163 -19527
rect 7763 -19597 7773 -19537
rect 7833 -19587 8093 -19537
rect 7833 -19597 7843 -19587
rect 7763 -19607 7843 -19597
rect 8083 -19597 8093 -19587
rect 8153 -19597 8163 -19537
rect 8083 -19607 8163 -19597
rect 7763 -19877 7823 -19607
rect 8093 -19617 8163 -19607
rect 7903 -19667 7933 -19647
rect 7883 -19707 7933 -19667
rect 7993 -19667 8023 -19647
rect 7993 -19707 8043 -19667
rect 7883 -19777 8043 -19707
rect 7883 -19817 7933 -19777
rect 7903 -19837 7933 -19817
rect 7993 -19817 8043 -19777
rect 7993 -19837 8023 -19817
rect 8103 -19877 8163 -19617
rect 7763 -19887 7843 -19877
rect 7763 -19947 7773 -19887
rect 7833 -19897 7843 -19887
rect 8083 -19887 8163 -19877
rect 8083 -19897 8093 -19887
rect 7833 -19947 8093 -19897
rect 8153 -19947 8163 -19887
rect 7763 -19957 8163 -19947
rect 8237 -19537 8637 -19527
rect 8237 -19597 8247 -19537
rect 8307 -19587 8567 -19537
rect 8307 -19597 8317 -19587
rect 8237 -19607 8317 -19597
rect 8557 -19597 8567 -19587
rect 8627 -19597 8637 -19537
rect 8557 -19607 8637 -19597
rect 8237 -19877 8297 -19607
rect 8567 -19617 8637 -19607
rect 8377 -19667 8407 -19647
rect 8357 -19707 8407 -19667
rect 8467 -19667 8497 -19647
rect 8467 -19707 8517 -19667
rect 8357 -19777 8517 -19707
rect 8357 -19817 8407 -19777
rect 8377 -19837 8407 -19817
rect 8467 -19817 8517 -19777
rect 8467 -19837 8497 -19817
rect 8577 -19877 8637 -19617
rect 8237 -19887 8317 -19877
rect 8237 -19947 8247 -19887
rect 8307 -19897 8317 -19887
rect 8557 -19887 8637 -19877
rect 8557 -19897 8567 -19887
rect 8307 -19947 8567 -19897
rect 8627 -19947 8637 -19887
rect 8237 -19957 8637 -19947
rect 8693 -19537 9093 -19527
rect 8693 -19597 8703 -19537
rect 8763 -19587 9023 -19537
rect 8763 -19597 8773 -19587
rect 8693 -19607 8773 -19597
rect 9013 -19597 9023 -19587
rect 9083 -19597 9093 -19537
rect 9013 -19607 9093 -19597
rect 8693 -19877 8753 -19607
rect 9023 -19617 9093 -19607
rect 8833 -19667 8863 -19647
rect 8813 -19707 8863 -19667
rect 8923 -19667 8953 -19647
rect 8923 -19707 8973 -19667
rect 8813 -19777 8973 -19707
rect 8813 -19817 8863 -19777
rect 8833 -19837 8863 -19817
rect 8923 -19817 8973 -19777
rect 8923 -19837 8953 -19817
rect 9033 -19877 9093 -19617
rect 8693 -19887 8773 -19877
rect 8693 -19947 8703 -19887
rect 8763 -19897 8773 -19887
rect 9013 -19887 9093 -19877
rect 9013 -19897 9023 -19887
rect 8763 -19947 9023 -19897
rect 9083 -19947 9093 -19887
rect 8693 -19957 9093 -19947
rect 9151 -19537 9551 -19527
rect 9151 -19597 9161 -19537
rect 9221 -19587 9481 -19537
rect 9221 -19597 9231 -19587
rect 9151 -19607 9231 -19597
rect 9471 -19597 9481 -19587
rect 9541 -19597 9551 -19537
rect 9471 -19607 9551 -19597
rect 9151 -19877 9211 -19607
rect 9481 -19617 9551 -19607
rect 9291 -19667 9321 -19647
rect 9271 -19707 9321 -19667
rect 9381 -19667 9411 -19647
rect 9381 -19707 9431 -19667
rect 9271 -19777 9431 -19707
rect 9271 -19817 9321 -19777
rect 9291 -19837 9321 -19817
rect 9381 -19817 9431 -19777
rect 9381 -19837 9411 -19817
rect 9491 -19877 9551 -19617
rect 9151 -19887 9231 -19877
rect 9151 -19947 9161 -19887
rect 9221 -19897 9231 -19887
rect 9471 -19887 9551 -19877
rect 9471 -19897 9481 -19887
rect 9221 -19947 9481 -19897
rect 9541 -19947 9551 -19887
rect 9151 -19957 9551 -19947
rect 9607 -19537 10007 -19527
rect 9607 -19597 9617 -19537
rect 9677 -19587 9937 -19537
rect 9677 -19597 9687 -19587
rect 9607 -19607 9687 -19597
rect 9927 -19597 9937 -19587
rect 9997 -19597 10007 -19537
rect 9927 -19607 10007 -19597
rect 9607 -19877 9667 -19607
rect 9937 -19617 10007 -19607
rect 9747 -19667 9777 -19647
rect 9727 -19707 9777 -19667
rect 9837 -19667 9867 -19647
rect 9837 -19707 9887 -19667
rect 9727 -19777 9887 -19707
rect 9727 -19817 9777 -19777
rect 9747 -19837 9777 -19817
rect 9837 -19817 9887 -19777
rect 9837 -19837 9867 -19817
rect 9947 -19877 10007 -19617
rect 9607 -19887 9687 -19877
rect 9607 -19947 9617 -19887
rect 9677 -19897 9687 -19887
rect 9927 -19887 10007 -19877
rect 9927 -19897 9937 -19887
rect 9677 -19947 9937 -19897
rect 9997 -19947 10007 -19887
rect 9607 -19957 10007 -19947
rect 10063 -19537 10463 -19527
rect 10063 -19597 10073 -19537
rect 10133 -19587 10393 -19537
rect 10133 -19597 10143 -19587
rect 10063 -19607 10143 -19597
rect 10383 -19597 10393 -19587
rect 10453 -19597 10463 -19537
rect 10383 -19607 10463 -19597
rect 10063 -19877 10123 -19607
rect 10393 -19617 10463 -19607
rect 10203 -19667 10233 -19647
rect 10183 -19707 10233 -19667
rect 10293 -19667 10323 -19647
rect 10293 -19707 10343 -19667
rect 10183 -19777 10343 -19707
rect 10183 -19817 10233 -19777
rect 10203 -19837 10233 -19817
rect 10293 -19817 10343 -19777
rect 10293 -19837 10323 -19817
rect 10403 -19877 10463 -19617
rect 10063 -19887 10143 -19877
rect 10063 -19947 10073 -19887
rect 10133 -19897 10143 -19887
rect 10383 -19887 10463 -19877
rect 10383 -19897 10393 -19887
rect 10133 -19947 10393 -19897
rect 10453 -19947 10463 -19887
rect 10063 -19957 10463 -19947
rect 10521 -19537 10921 -19527
rect 10521 -19597 10531 -19537
rect 10591 -19587 10851 -19537
rect 10591 -19597 10601 -19587
rect 10521 -19607 10601 -19597
rect 10841 -19597 10851 -19587
rect 10911 -19597 10921 -19537
rect 10841 -19607 10921 -19597
rect 10521 -19877 10581 -19607
rect 10851 -19617 10921 -19607
rect 10661 -19667 10691 -19647
rect 10641 -19707 10691 -19667
rect 10751 -19667 10781 -19647
rect 10751 -19707 10801 -19667
rect 10641 -19777 10801 -19707
rect 10641 -19817 10691 -19777
rect 10661 -19837 10691 -19817
rect 10751 -19817 10801 -19777
rect 10751 -19837 10781 -19817
rect 10861 -19877 10921 -19617
rect 10521 -19887 10601 -19877
rect 10521 -19947 10531 -19887
rect 10591 -19897 10601 -19887
rect 10841 -19887 10921 -19877
rect 10841 -19897 10851 -19887
rect 10591 -19947 10851 -19897
rect 10911 -19947 10921 -19887
rect 10521 -19957 10921 -19947
rect 10977 -19537 11377 -19527
rect 10977 -19597 10987 -19537
rect 11047 -19587 11307 -19537
rect 11047 -19597 11057 -19587
rect 10977 -19607 11057 -19597
rect 11297 -19597 11307 -19587
rect 11367 -19597 11377 -19537
rect 11297 -19607 11377 -19597
rect 10977 -19877 11037 -19607
rect 11307 -19617 11377 -19607
rect 11117 -19667 11147 -19647
rect 11097 -19707 11147 -19667
rect 11207 -19667 11237 -19647
rect 11207 -19707 11257 -19667
rect 11097 -19777 11257 -19707
rect 11097 -19817 11147 -19777
rect 11117 -19837 11147 -19817
rect 11207 -19817 11257 -19777
rect 11207 -19837 11237 -19817
rect 11317 -19877 11377 -19617
rect 10977 -19887 11057 -19877
rect 10977 -19947 10987 -19887
rect 11047 -19897 11057 -19887
rect 11297 -19887 11377 -19877
rect 11297 -19897 11307 -19887
rect 11047 -19947 11307 -19897
rect 11367 -19947 11377 -19887
rect 10977 -19957 11377 -19947
rect 11433 -19537 11833 -19527
rect 11433 -19597 11443 -19537
rect 11503 -19587 11763 -19537
rect 11503 -19597 11513 -19587
rect 11433 -19607 11513 -19597
rect 11753 -19597 11763 -19587
rect 11823 -19597 11833 -19537
rect 11753 -19607 11833 -19597
rect 11433 -19877 11493 -19607
rect 11763 -19617 11833 -19607
rect 11573 -19667 11603 -19647
rect 11553 -19707 11603 -19667
rect 11663 -19667 11693 -19647
rect 11663 -19707 11713 -19667
rect 11553 -19777 11713 -19707
rect 11553 -19817 11603 -19777
rect 11573 -19837 11603 -19817
rect 11663 -19817 11713 -19777
rect 11663 -19837 11693 -19817
rect 11773 -19877 11833 -19617
rect 11433 -19887 11513 -19877
rect 11433 -19947 11443 -19887
rect 11503 -19897 11513 -19887
rect 11753 -19887 11833 -19877
rect 11753 -19897 11763 -19887
rect 11503 -19947 11763 -19897
rect 11823 -19947 11833 -19887
rect 11433 -19957 11833 -19947
rect 11891 -19537 12291 -19527
rect 11891 -19597 11901 -19537
rect 11961 -19587 12221 -19537
rect 11961 -19597 11971 -19587
rect 11891 -19607 11971 -19597
rect 12211 -19597 12221 -19587
rect 12281 -19597 12291 -19537
rect 12211 -19607 12291 -19597
rect 11891 -19877 11951 -19607
rect 12221 -19617 12291 -19607
rect 12031 -19667 12061 -19647
rect 12011 -19707 12061 -19667
rect 12121 -19667 12151 -19647
rect 12121 -19707 12171 -19667
rect 12011 -19777 12171 -19707
rect 12011 -19817 12061 -19777
rect 12031 -19837 12061 -19817
rect 12121 -19817 12171 -19777
rect 12121 -19837 12151 -19817
rect 12231 -19877 12291 -19617
rect 11891 -19887 11971 -19877
rect 11891 -19947 11901 -19887
rect 11961 -19897 11971 -19887
rect 12211 -19887 12291 -19877
rect 12211 -19897 12221 -19887
rect 11961 -19947 12221 -19897
rect 12281 -19947 12291 -19887
rect 11891 -19957 12291 -19947
rect 12347 -19537 12747 -19527
rect 12347 -19597 12357 -19537
rect 12417 -19587 12677 -19537
rect 12417 -19597 12427 -19587
rect 12347 -19607 12427 -19597
rect 12667 -19597 12677 -19587
rect 12737 -19597 12747 -19537
rect 12667 -19607 12747 -19597
rect 12347 -19877 12407 -19607
rect 12677 -19617 12747 -19607
rect 12487 -19667 12517 -19647
rect 12467 -19707 12517 -19667
rect 12577 -19667 12607 -19647
rect 12577 -19707 12627 -19667
rect 12467 -19777 12627 -19707
rect 12467 -19817 12517 -19777
rect 12487 -19837 12517 -19817
rect 12577 -19817 12627 -19777
rect 12577 -19837 12607 -19817
rect 12687 -19877 12747 -19617
rect 12347 -19887 12427 -19877
rect 12347 -19947 12357 -19887
rect 12417 -19897 12427 -19887
rect 12667 -19887 12747 -19877
rect 12667 -19897 12677 -19887
rect 12417 -19947 12677 -19897
rect 12737 -19947 12747 -19887
rect 12347 -19957 12747 -19947
rect 12803 -19537 13203 -19527
rect 12803 -19597 12813 -19537
rect 12873 -19587 13133 -19537
rect 12873 -19597 12883 -19587
rect 12803 -19607 12883 -19597
rect 13123 -19597 13133 -19587
rect 13193 -19597 13203 -19537
rect 13123 -19607 13203 -19597
rect 12803 -19877 12863 -19607
rect 13133 -19617 13203 -19607
rect 12943 -19667 12973 -19647
rect 12923 -19707 12973 -19667
rect 13033 -19667 13063 -19647
rect 13033 -19707 13083 -19667
rect 12923 -19777 13083 -19707
rect 12923 -19817 12973 -19777
rect 12943 -19837 12973 -19817
rect 13033 -19817 13083 -19777
rect 13033 -19837 13063 -19817
rect 13143 -19877 13203 -19617
rect 12803 -19887 12883 -19877
rect 12803 -19947 12813 -19887
rect 12873 -19897 12883 -19887
rect 13123 -19887 13203 -19877
rect 13123 -19897 13133 -19887
rect 12873 -19947 13133 -19897
rect 13193 -19947 13203 -19887
rect 12803 -19957 13203 -19947
rect 13261 -19537 13661 -19527
rect 13261 -19597 13271 -19537
rect 13331 -19587 13591 -19537
rect 13331 -19597 13341 -19587
rect 13261 -19607 13341 -19597
rect 13581 -19597 13591 -19587
rect 13651 -19597 13661 -19537
rect 13581 -19607 13661 -19597
rect 13261 -19877 13321 -19607
rect 13591 -19617 13661 -19607
rect 13401 -19667 13431 -19647
rect 13381 -19707 13431 -19667
rect 13491 -19667 13521 -19647
rect 13491 -19707 13541 -19667
rect 13381 -19777 13541 -19707
rect 13381 -19817 13431 -19777
rect 13401 -19837 13431 -19817
rect 13491 -19817 13541 -19777
rect 13491 -19837 13521 -19817
rect 13601 -19877 13661 -19617
rect 13261 -19887 13341 -19877
rect 13261 -19947 13271 -19887
rect 13331 -19897 13341 -19887
rect 13581 -19887 13661 -19877
rect 13581 -19897 13591 -19887
rect 13331 -19947 13591 -19897
rect 13651 -19947 13661 -19887
rect 13261 -19957 13661 -19947
rect 13717 -19537 14117 -19527
rect 13717 -19597 13727 -19537
rect 13787 -19587 14047 -19537
rect 13787 -19597 13797 -19587
rect 13717 -19607 13797 -19597
rect 14037 -19597 14047 -19587
rect 14107 -19597 14117 -19537
rect 14037 -19607 14117 -19597
rect 13717 -19877 13777 -19607
rect 14047 -19617 14117 -19607
rect 13857 -19667 13887 -19647
rect 13837 -19707 13887 -19667
rect 13947 -19667 13977 -19647
rect 13947 -19707 13997 -19667
rect 13837 -19777 13997 -19707
rect 13837 -19817 13887 -19777
rect 13857 -19837 13887 -19817
rect 13947 -19817 13997 -19777
rect 13947 -19837 13977 -19817
rect 14057 -19877 14117 -19617
rect 13717 -19887 13797 -19877
rect 13717 -19947 13727 -19887
rect 13787 -19897 13797 -19887
rect 14037 -19887 14117 -19877
rect 14037 -19897 14047 -19887
rect 13787 -19947 14047 -19897
rect 14107 -19947 14117 -19887
rect 13717 -19957 14117 -19947
rect 14173 -19537 14573 -19527
rect 14173 -19597 14183 -19537
rect 14243 -19587 14503 -19537
rect 14243 -19597 14253 -19587
rect 14173 -19607 14253 -19597
rect 14493 -19597 14503 -19587
rect 14563 -19597 14573 -19537
rect 14493 -19607 14573 -19597
rect 14173 -19877 14233 -19607
rect 14503 -19617 14573 -19607
rect 14313 -19667 14343 -19647
rect 14293 -19707 14343 -19667
rect 14403 -19667 14433 -19647
rect 14403 -19707 14453 -19667
rect 14293 -19777 14453 -19707
rect 14293 -19817 14343 -19777
rect 14313 -19837 14343 -19817
rect 14403 -19817 14453 -19777
rect 14403 -19837 14433 -19817
rect 14513 -19877 14573 -19617
rect 14173 -19887 14253 -19877
rect 14173 -19947 14183 -19887
rect 14243 -19897 14253 -19887
rect 14493 -19887 14573 -19877
rect 14493 -19897 14503 -19887
rect 14243 -19947 14503 -19897
rect 14563 -19947 14573 -19887
rect 14173 -19957 14573 -19947
rect 14631 -19537 15031 -19527
rect 14631 -19597 14641 -19537
rect 14701 -19587 14961 -19537
rect 14701 -19597 14711 -19587
rect 14631 -19607 14711 -19597
rect 14951 -19597 14961 -19587
rect 15021 -19597 15031 -19537
rect 14951 -19607 15031 -19597
rect 14631 -19877 14691 -19607
rect 14961 -19617 15031 -19607
rect 14771 -19667 14801 -19647
rect 14751 -19707 14801 -19667
rect 14861 -19667 14891 -19647
rect 14861 -19707 14911 -19667
rect 14751 -19777 14911 -19707
rect 14751 -19817 14801 -19777
rect 14771 -19837 14801 -19817
rect 14861 -19817 14911 -19777
rect 14861 -19837 14891 -19817
rect 14971 -19877 15031 -19617
rect 14631 -19887 14711 -19877
rect 14631 -19947 14641 -19887
rect 14701 -19897 14711 -19887
rect 14951 -19887 15031 -19877
rect 14951 -19897 14961 -19887
rect 14701 -19947 14961 -19897
rect 15021 -19947 15031 -19887
rect 14631 -19957 15031 -19947
rect 15087 -19537 15487 -19527
rect 15087 -19597 15097 -19537
rect 15157 -19587 15417 -19537
rect 15157 -19597 15167 -19587
rect 15087 -19607 15167 -19597
rect 15407 -19597 15417 -19587
rect 15477 -19597 15487 -19537
rect 15407 -19607 15487 -19597
rect 15087 -19877 15147 -19607
rect 15417 -19617 15487 -19607
rect 15227 -19667 15257 -19647
rect 15207 -19707 15257 -19667
rect 15317 -19667 15347 -19647
rect 15317 -19707 15367 -19667
rect 15207 -19777 15367 -19707
rect 15207 -19817 15257 -19777
rect 15227 -19837 15257 -19817
rect 15317 -19817 15367 -19777
rect 15317 -19837 15347 -19817
rect 15427 -19877 15487 -19617
rect 15087 -19887 15167 -19877
rect 15087 -19947 15097 -19887
rect 15157 -19897 15167 -19887
rect 15407 -19887 15487 -19877
rect 15407 -19897 15417 -19887
rect 15157 -19947 15417 -19897
rect 15477 -19947 15487 -19887
rect 15087 -19957 15487 -19947
rect 1 -20039 401 -20029
rect 1 -20099 11 -20039
rect 71 -20089 331 -20039
rect 71 -20099 81 -20089
rect 1 -20109 81 -20099
rect 321 -20099 331 -20089
rect 391 -20099 401 -20039
rect 321 -20109 401 -20099
rect 1 -20379 61 -20109
rect 331 -20119 401 -20109
rect 141 -20169 171 -20149
rect 121 -20209 171 -20169
rect 231 -20169 261 -20149
rect 231 -20209 281 -20169
rect 121 -20279 281 -20209
rect 121 -20319 171 -20279
rect 141 -20339 171 -20319
rect 231 -20319 281 -20279
rect 231 -20339 261 -20319
rect 341 -20379 401 -20119
rect 1 -20389 81 -20379
rect 1 -20449 11 -20389
rect 71 -20399 81 -20389
rect 321 -20389 401 -20379
rect 321 -20399 331 -20389
rect 71 -20449 331 -20399
rect 391 -20449 401 -20389
rect 1 -20459 401 -20449
rect 457 -20039 857 -20029
rect 457 -20099 467 -20039
rect 527 -20089 787 -20039
rect 527 -20099 537 -20089
rect 457 -20109 537 -20099
rect 777 -20099 787 -20089
rect 847 -20099 857 -20039
rect 777 -20109 857 -20099
rect 457 -20379 517 -20109
rect 787 -20119 857 -20109
rect 597 -20169 627 -20149
rect 577 -20209 627 -20169
rect 687 -20169 717 -20149
rect 687 -20209 737 -20169
rect 577 -20279 737 -20209
rect 577 -20319 627 -20279
rect 597 -20339 627 -20319
rect 687 -20319 737 -20279
rect 687 -20339 717 -20319
rect 797 -20379 857 -20119
rect 457 -20389 537 -20379
rect 457 -20449 467 -20389
rect 527 -20399 537 -20389
rect 777 -20389 857 -20379
rect 777 -20399 787 -20389
rect 527 -20449 787 -20399
rect 847 -20449 857 -20389
rect 457 -20459 857 -20449
rect 913 -20039 1313 -20029
rect 913 -20099 923 -20039
rect 983 -20089 1243 -20039
rect 983 -20099 993 -20089
rect 913 -20109 993 -20099
rect 1233 -20099 1243 -20089
rect 1303 -20099 1313 -20039
rect 1233 -20109 1313 -20099
rect 913 -20379 973 -20109
rect 1243 -20119 1313 -20109
rect 1053 -20169 1083 -20149
rect 1033 -20209 1083 -20169
rect 1143 -20169 1173 -20149
rect 1143 -20209 1193 -20169
rect 1033 -20279 1193 -20209
rect 1033 -20319 1083 -20279
rect 1053 -20339 1083 -20319
rect 1143 -20319 1193 -20279
rect 1143 -20339 1173 -20319
rect 1253 -20379 1313 -20119
rect 913 -20389 993 -20379
rect 913 -20449 923 -20389
rect 983 -20399 993 -20389
rect 1233 -20389 1313 -20379
rect 1233 -20399 1243 -20389
rect 983 -20449 1243 -20399
rect 1303 -20449 1313 -20389
rect 913 -20459 1313 -20449
rect 1371 -20039 1771 -20029
rect 1371 -20099 1381 -20039
rect 1441 -20089 1701 -20039
rect 1441 -20099 1451 -20089
rect 1371 -20109 1451 -20099
rect 1691 -20099 1701 -20089
rect 1761 -20099 1771 -20039
rect 1691 -20109 1771 -20099
rect 1371 -20379 1431 -20109
rect 1701 -20119 1771 -20109
rect 1511 -20169 1541 -20149
rect 1491 -20209 1541 -20169
rect 1601 -20169 1631 -20149
rect 1601 -20209 1651 -20169
rect 1491 -20279 1651 -20209
rect 1491 -20319 1541 -20279
rect 1511 -20339 1541 -20319
rect 1601 -20319 1651 -20279
rect 1601 -20339 1631 -20319
rect 1711 -20379 1771 -20119
rect 1371 -20389 1451 -20379
rect 1371 -20449 1381 -20389
rect 1441 -20399 1451 -20389
rect 1691 -20389 1771 -20379
rect 1691 -20399 1701 -20389
rect 1441 -20449 1701 -20399
rect 1761 -20449 1771 -20389
rect 1371 -20459 1771 -20449
rect 1827 -20039 2227 -20029
rect 1827 -20099 1837 -20039
rect 1897 -20089 2157 -20039
rect 1897 -20099 1907 -20089
rect 1827 -20109 1907 -20099
rect 2147 -20099 2157 -20089
rect 2217 -20099 2227 -20039
rect 2147 -20109 2227 -20099
rect 1827 -20379 1887 -20109
rect 2157 -20119 2227 -20109
rect 1967 -20169 1997 -20149
rect 1947 -20209 1997 -20169
rect 2057 -20169 2087 -20149
rect 2057 -20209 2107 -20169
rect 1947 -20279 2107 -20209
rect 1947 -20319 1997 -20279
rect 1967 -20339 1997 -20319
rect 2057 -20319 2107 -20279
rect 2057 -20339 2087 -20319
rect 2167 -20379 2227 -20119
rect 1827 -20389 1907 -20379
rect 1827 -20449 1837 -20389
rect 1897 -20399 1907 -20389
rect 2147 -20389 2227 -20379
rect 2147 -20399 2157 -20389
rect 1897 -20449 2157 -20399
rect 2217 -20449 2227 -20389
rect 1827 -20459 2227 -20449
rect 2283 -20039 2683 -20029
rect 2283 -20099 2293 -20039
rect 2353 -20089 2613 -20039
rect 2353 -20099 2363 -20089
rect 2283 -20109 2363 -20099
rect 2603 -20099 2613 -20089
rect 2673 -20099 2683 -20039
rect 2603 -20109 2683 -20099
rect 2283 -20379 2343 -20109
rect 2613 -20119 2683 -20109
rect 2423 -20169 2453 -20149
rect 2403 -20209 2453 -20169
rect 2513 -20169 2543 -20149
rect 2513 -20209 2563 -20169
rect 2403 -20279 2563 -20209
rect 2403 -20319 2453 -20279
rect 2423 -20339 2453 -20319
rect 2513 -20319 2563 -20279
rect 2513 -20339 2543 -20319
rect 2623 -20379 2683 -20119
rect 2283 -20389 2363 -20379
rect 2283 -20449 2293 -20389
rect 2353 -20399 2363 -20389
rect 2603 -20389 2683 -20379
rect 2603 -20399 2613 -20389
rect 2353 -20449 2613 -20399
rect 2673 -20449 2683 -20389
rect 2283 -20459 2683 -20449
rect 2741 -20039 3141 -20029
rect 2741 -20099 2751 -20039
rect 2811 -20089 3071 -20039
rect 2811 -20099 2821 -20089
rect 2741 -20109 2821 -20099
rect 3061 -20099 3071 -20089
rect 3131 -20099 3141 -20039
rect 3061 -20109 3141 -20099
rect 2741 -20379 2801 -20109
rect 3071 -20119 3141 -20109
rect 2881 -20169 2911 -20149
rect 2861 -20209 2911 -20169
rect 2971 -20169 3001 -20149
rect 2971 -20209 3021 -20169
rect 2861 -20279 3021 -20209
rect 2861 -20319 2911 -20279
rect 2881 -20339 2911 -20319
rect 2971 -20319 3021 -20279
rect 2971 -20339 3001 -20319
rect 3081 -20379 3141 -20119
rect 2741 -20389 2821 -20379
rect 2741 -20449 2751 -20389
rect 2811 -20399 2821 -20389
rect 3061 -20389 3141 -20379
rect 3061 -20399 3071 -20389
rect 2811 -20449 3071 -20399
rect 3131 -20449 3141 -20389
rect 2741 -20459 3141 -20449
rect 3197 -20039 3597 -20029
rect 3197 -20099 3207 -20039
rect 3267 -20089 3527 -20039
rect 3267 -20099 3277 -20089
rect 3197 -20109 3277 -20099
rect 3517 -20099 3527 -20089
rect 3587 -20099 3597 -20039
rect 3517 -20109 3597 -20099
rect 3197 -20379 3257 -20109
rect 3527 -20119 3597 -20109
rect 3337 -20169 3367 -20149
rect 3317 -20209 3367 -20169
rect 3427 -20169 3457 -20149
rect 3427 -20209 3477 -20169
rect 3317 -20279 3477 -20209
rect 3317 -20319 3367 -20279
rect 3337 -20339 3367 -20319
rect 3427 -20319 3477 -20279
rect 3427 -20339 3457 -20319
rect 3537 -20379 3597 -20119
rect 3197 -20389 3277 -20379
rect 3197 -20449 3207 -20389
rect 3267 -20399 3277 -20389
rect 3517 -20389 3597 -20379
rect 3517 -20399 3527 -20389
rect 3267 -20449 3527 -20399
rect 3587 -20449 3597 -20389
rect 3197 -20459 3597 -20449
rect 3653 -20039 4053 -20029
rect 3653 -20099 3663 -20039
rect 3723 -20089 3983 -20039
rect 3723 -20099 3733 -20089
rect 3653 -20109 3733 -20099
rect 3973 -20099 3983 -20089
rect 4043 -20099 4053 -20039
rect 3973 -20109 4053 -20099
rect 3653 -20379 3713 -20109
rect 3983 -20119 4053 -20109
rect 3793 -20169 3823 -20149
rect 3773 -20209 3823 -20169
rect 3883 -20169 3913 -20149
rect 3883 -20209 3933 -20169
rect 3773 -20279 3933 -20209
rect 3773 -20319 3823 -20279
rect 3793 -20339 3823 -20319
rect 3883 -20319 3933 -20279
rect 3883 -20339 3913 -20319
rect 3993 -20379 4053 -20119
rect 3653 -20389 3733 -20379
rect 3653 -20449 3663 -20389
rect 3723 -20399 3733 -20389
rect 3973 -20389 4053 -20379
rect 3973 -20399 3983 -20389
rect 3723 -20449 3983 -20399
rect 4043 -20449 4053 -20389
rect 3653 -20459 4053 -20449
rect 4111 -20039 4511 -20029
rect 4111 -20099 4121 -20039
rect 4181 -20089 4441 -20039
rect 4181 -20099 4191 -20089
rect 4111 -20109 4191 -20099
rect 4431 -20099 4441 -20089
rect 4501 -20099 4511 -20039
rect 4431 -20109 4511 -20099
rect 4111 -20379 4171 -20109
rect 4441 -20119 4511 -20109
rect 4251 -20169 4281 -20149
rect 4231 -20209 4281 -20169
rect 4341 -20169 4371 -20149
rect 4341 -20209 4391 -20169
rect 4231 -20279 4391 -20209
rect 4231 -20319 4281 -20279
rect 4251 -20339 4281 -20319
rect 4341 -20319 4391 -20279
rect 4341 -20339 4371 -20319
rect 4451 -20379 4511 -20119
rect 4111 -20389 4191 -20379
rect 4111 -20449 4121 -20389
rect 4181 -20399 4191 -20389
rect 4431 -20389 4511 -20379
rect 4431 -20399 4441 -20389
rect 4181 -20449 4441 -20399
rect 4501 -20449 4511 -20389
rect 4111 -20459 4511 -20449
rect 4567 -20039 4967 -20029
rect 4567 -20099 4577 -20039
rect 4637 -20089 4897 -20039
rect 4637 -20099 4647 -20089
rect 4567 -20109 4647 -20099
rect 4887 -20099 4897 -20089
rect 4957 -20099 4967 -20039
rect 4887 -20109 4967 -20099
rect 4567 -20379 4627 -20109
rect 4897 -20119 4967 -20109
rect 4707 -20169 4737 -20149
rect 4687 -20209 4737 -20169
rect 4797 -20169 4827 -20149
rect 4797 -20209 4847 -20169
rect 4687 -20279 4847 -20209
rect 4687 -20319 4737 -20279
rect 4707 -20339 4737 -20319
rect 4797 -20319 4847 -20279
rect 4797 -20339 4827 -20319
rect 4907 -20379 4967 -20119
rect 4567 -20389 4647 -20379
rect 4567 -20449 4577 -20389
rect 4637 -20399 4647 -20389
rect 4887 -20389 4967 -20379
rect 4887 -20399 4897 -20389
rect 4637 -20449 4897 -20399
rect 4957 -20449 4967 -20389
rect 4567 -20459 4967 -20449
rect 5023 -20039 5423 -20029
rect 5023 -20099 5033 -20039
rect 5093 -20089 5353 -20039
rect 5093 -20099 5103 -20089
rect 5023 -20109 5103 -20099
rect 5343 -20099 5353 -20089
rect 5413 -20099 5423 -20039
rect 5343 -20109 5423 -20099
rect 5023 -20379 5083 -20109
rect 5353 -20119 5423 -20109
rect 5163 -20169 5193 -20149
rect 5143 -20209 5193 -20169
rect 5253 -20169 5283 -20149
rect 5253 -20209 5303 -20169
rect 5143 -20279 5303 -20209
rect 5143 -20319 5193 -20279
rect 5163 -20339 5193 -20319
rect 5253 -20319 5303 -20279
rect 5253 -20339 5283 -20319
rect 5363 -20379 5423 -20119
rect 5023 -20389 5103 -20379
rect 5023 -20449 5033 -20389
rect 5093 -20399 5103 -20389
rect 5343 -20389 5423 -20379
rect 5343 -20399 5353 -20389
rect 5093 -20449 5353 -20399
rect 5413 -20449 5423 -20389
rect 5023 -20459 5423 -20449
rect 5481 -20039 5881 -20029
rect 5481 -20099 5491 -20039
rect 5551 -20089 5811 -20039
rect 5551 -20099 5561 -20089
rect 5481 -20109 5561 -20099
rect 5801 -20099 5811 -20089
rect 5871 -20099 5881 -20039
rect 5801 -20109 5881 -20099
rect 5481 -20379 5541 -20109
rect 5811 -20119 5881 -20109
rect 5621 -20169 5651 -20149
rect 5601 -20209 5651 -20169
rect 5711 -20169 5741 -20149
rect 5711 -20209 5761 -20169
rect 5601 -20279 5761 -20209
rect 5601 -20319 5651 -20279
rect 5621 -20339 5651 -20319
rect 5711 -20319 5761 -20279
rect 5711 -20339 5741 -20319
rect 5821 -20379 5881 -20119
rect 5481 -20389 5561 -20379
rect 5481 -20449 5491 -20389
rect 5551 -20399 5561 -20389
rect 5801 -20389 5881 -20379
rect 5801 -20399 5811 -20389
rect 5551 -20449 5811 -20399
rect 5871 -20449 5881 -20389
rect 5481 -20459 5881 -20449
rect 5937 -20039 6337 -20029
rect 5937 -20099 5947 -20039
rect 6007 -20089 6267 -20039
rect 6007 -20099 6017 -20089
rect 5937 -20109 6017 -20099
rect 6257 -20099 6267 -20089
rect 6327 -20099 6337 -20039
rect 6257 -20109 6337 -20099
rect 5937 -20379 5997 -20109
rect 6267 -20119 6337 -20109
rect 6077 -20169 6107 -20149
rect 6057 -20209 6107 -20169
rect 6167 -20169 6197 -20149
rect 6167 -20209 6217 -20169
rect 6057 -20279 6217 -20209
rect 6057 -20319 6107 -20279
rect 6077 -20339 6107 -20319
rect 6167 -20319 6217 -20279
rect 6167 -20339 6197 -20319
rect 6277 -20379 6337 -20119
rect 5937 -20389 6017 -20379
rect 5937 -20449 5947 -20389
rect 6007 -20399 6017 -20389
rect 6257 -20389 6337 -20379
rect 6257 -20399 6267 -20389
rect 6007 -20449 6267 -20399
rect 6327 -20449 6337 -20389
rect 5937 -20459 6337 -20449
rect 6393 -20039 6793 -20029
rect 6393 -20099 6403 -20039
rect 6463 -20089 6723 -20039
rect 6463 -20099 6473 -20089
rect 6393 -20109 6473 -20099
rect 6713 -20099 6723 -20089
rect 6783 -20099 6793 -20039
rect 6713 -20109 6793 -20099
rect 6393 -20379 6453 -20109
rect 6723 -20119 6793 -20109
rect 6533 -20169 6563 -20149
rect 6513 -20209 6563 -20169
rect 6623 -20169 6653 -20149
rect 6623 -20209 6673 -20169
rect 6513 -20279 6673 -20209
rect 6513 -20319 6563 -20279
rect 6533 -20339 6563 -20319
rect 6623 -20319 6673 -20279
rect 6623 -20339 6653 -20319
rect 6733 -20379 6793 -20119
rect 6393 -20389 6473 -20379
rect 6393 -20449 6403 -20389
rect 6463 -20399 6473 -20389
rect 6713 -20389 6793 -20379
rect 6713 -20399 6723 -20389
rect 6463 -20449 6723 -20399
rect 6783 -20449 6793 -20389
rect 6393 -20459 6793 -20449
rect 6851 -20039 7251 -20029
rect 6851 -20099 6861 -20039
rect 6921 -20089 7181 -20039
rect 6921 -20099 6931 -20089
rect 6851 -20109 6931 -20099
rect 7171 -20099 7181 -20089
rect 7241 -20099 7251 -20039
rect 7171 -20109 7251 -20099
rect 6851 -20379 6911 -20109
rect 7181 -20119 7251 -20109
rect 6991 -20169 7021 -20149
rect 6971 -20209 7021 -20169
rect 7081 -20169 7111 -20149
rect 7081 -20209 7131 -20169
rect 6971 -20279 7131 -20209
rect 6971 -20319 7021 -20279
rect 6991 -20339 7021 -20319
rect 7081 -20319 7131 -20279
rect 7081 -20339 7111 -20319
rect 7191 -20379 7251 -20119
rect 6851 -20389 6931 -20379
rect 6851 -20449 6861 -20389
rect 6921 -20399 6931 -20389
rect 7171 -20389 7251 -20379
rect 7171 -20399 7181 -20389
rect 6921 -20449 7181 -20399
rect 7241 -20449 7251 -20389
rect 6851 -20459 7251 -20449
rect 7307 -20039 7707 -20029
rect 7307 -20099 7317 -20039
rect 7377 -20089 7637 -20039
rect 7377 -20099 7387 -20089
rect 7307 -20109 7387 -20099
rect 7627 -20099 7637 -20089
rect 7697 -20099 7707 -20039
rect 7627 -20109 7707 -20099
rect 7307 -20379 7367 -20109
rect 7637 -20119 7707 -20109
rect 7447 -20169 7477 -20149
rect 7427 -20209 7477 -20169
rect 7537 -20169 7567 -20149
rect 7537 -20209 7587 -20169
rect 7427 -20279 7587 -20209
rect 7427 -20319 7477 -20279
rect 7447 -20339 7477 -20319
rect 7537 -20319 7587 -20279
rect 7537 -20339 7567 -20319
rect 7647 -20379 7707 -20119
rect 7307 -20389 7387 -20379
rect 7307 -20449 7317 -20389
rect 7377 -20399 7387 -20389
rect 7627 -20389 7707 -20379
rect 7627 -20399 7637 -20389
rect 7377 -20449 7637 -20399
rect 7697 -20449 7707 -20389
rect 7307 -20459 7707 -20449
rect 7763 -20039 8163 -20029
rect 7763 -20099 7773 -20039
rect 7833 -20089 8093 -20039
rect 7833 -20099 7843 -20089
rect 7763 -20109 7843 -20099
rect 8083 -20099 8093 -20089
rect 8153 -20099 8163 -20039
rect 8083 -20109 8163 -20099
rect 7763 -20379 7823 -20109
rect 8093 -20119 8163 -20109
rect 7903 -20169 7933 -20149
rect 7883 -20209 7933 -20169
rect 7993 -20169 8023 -20149
rect 7993 -20209 8043 -20169
rect 7883 -20279 8043 -20209
rect 7883 -20319 7933 -20279
rect 7903 -20339 7933 -20319
rect 7993 -20319 8043 -20279
rect 7993 -20339 8023 -20319
rect 8103 -20379 8163 -20119
rect 7763 -20389 7843 -20379
rect 7763 -20449 7773 -20389
rect 7833 -20399 7843 -20389
rect 8083 -20389 8163 -20379
rect 8083 -20399 8093 -20389
rect 7833 -20449 8093 -20399
rect 8153 -20449 8163 -20389
rect 7763 -20459 8163 -20449
rect 8237 -20039 8637 -20029
rect 8237 -20099 8247 -20039
rect 8307 -20089 8567 -20039
rect 8307 -20099 8317 -20089
rect 8237 -20109 8317 -20099
rect 8557 -20099 8567 -20089
rect 8627 -20099 8637 -20039
rect 8557 -20109 8637 -20099
rect 8237 -20379 8297 -20109
rect 8567 -20119 8637 -20109
rect 8377 -20169 8407 -20149
rect 8357 -20209 8407 -20169
rect 8467 -20169 8497 -20149
rect 8467 -20209 8517 -20169
rect 8357 -20279 8517 -20209
rect 8357 -20319 8407 -20279
rect 8377 -20339 8407 -20319
rect 8467 -20319 8517 -20279
rect 8467 -20339 8497 -20319
rect 8577 -20379 8637 -20119
rect 8237 -20389 8317 -20379
rect 8237 -20449 8247 -20389
rect 8307 -20399 8317 -20389
rect 8557 -20389 8637 -20379
rect 8557 -20399 8567 -20389
rect 8307 -20449 8567 -20399
rect 8627 -20449 8637 -20389
rect 8237 -20459 8637 -20449
rect 8693 -20039 9093 -20029
rect 8693 -20099 8703 -20039
rect 8763 -20089 9023 -20039
rect 8763 -20099 8773 -20089
rect 8693 -20109 8773 -20099
rect 9013 -20099 9023 -20089
rect 9083 -20099 9093 -20039
rect 9013 -20109 9093 -20099
rect 8693 -20379 8753 -20109
rect 9023 -20119 9093 -20109
rect 8833 -20169 8863 -20149
rect 8813 -20209 8863 -20169
rect 8923 -20169 8953 -20149
rect 8923 -20209 8973 -20169
rect 8813 -20279 8973 -20209
rect 8813 -20319 8863 -20279
rect 8833 -20339 8863 -20319
rect 8923 -20319 8973 -20279
rect 8923 -20339 8953 -20319
rect 9033 -20379 9093 -20119
rect 8693 -20389 8773 -20379
rect 8693 -20449 8703 -20389
rect 8763 -20399 8773 -20389
rect 9013 -20389 9093 -20379
rect 9013 -20399 9023 -20389
rect 8763 -20449 9023 -20399
rect 9083 -20449 9093 -20389
rect 8693 -20459 9093 -20449
rect 9151 -20039 9551 -20029
rect 9151 -20099 9161 -20039
rect 9221 -20089 9481 -20039
rect 9221 -20099 9231 -20089
rect 9151 -20109 9231 -20099
rect 9471 -20099 9481 -20089
rect 9541 -20099 9551 -20039
rect 9471 -20109 9551 -20099
rect 9151 -20379 9211 -20109
rect 9481 -20119 9551 -20109
rect 9291 -20169 9321 -20149
rect 9271 -20209 9321 -20169
rect 9381 -20169 9411 -20149
rect 9381 -20209 9431 -20169
rect 9271 -20279 9431 -20209
rect 9271 -20319 9321 -20279
rect 9291 -20339 9321 -20319
rect 9381 -20319 9431 -20279
rect 9381 -20339 9411 -20319
rect 9491 -20379 9551 -20119
rect 9151 -20389 9231 -20379
rect 9151 -20449 9161 -20389
rect 9221 -20399 9231 -20389
rect 9471 -20389 9551 -20379
rect 9471 -20399 9481 -20389
rect 9221 -20449 9481 -20399
rect 9541 -20449 9551 -20389
rect 9151 -20459 9551 -20449
rect 9607 -20039 10007 -20029
rect 9607 -20099 9617 -20039
rect 9677 -20089 9937 -20039
rect 9677 -20099 9687 -20089
rect 9607 -20109 9687 -20099
rect 9927 -20099 9937 -20089
rect 9997 -20099 10007 -20039
rect 9927 -20109 10007 -20099
rect 9607 -20379 9667 -20109
rect 9937 -20119 10007 -20109
rect 9747 -20169 9777 -20149
rect 9727 -20209 9777 -20169
rect 9837 -20169 9867 -20149
rect 9837 -20209 9887 -20169
rect 9727 -20279 9887 -20209
rect 9727 -20319 9777 -20279
rect 9747 -20339 9777 -20319
rect 9837 -20319 9887 -20279
rect 9837 -20339 9867 -20319
rect 9947 -20379 10007 -20119
rect 9607 -20389 9687 -20379
rect 9607 -20449 9617 -20389
rect 9677 -20399 9687 -20389
rect 9927 -20389 10007 -20379
rect 9927 -20399 9937 -20389
rect 9677 -20449 9937 -20399
rect 9997 -20449 10007 -20389
rect 9607 -20459 10007 -20449
rect 10063 -20039 10463 -20029
rect 10063 -20099 10073 -20039
rect 10133 -20089 10393 -20039
rect 10133 -20099 10143 -20089
rect 10063 -20109 10143 -20099
rect 10383 -20099 10393 -20089
rect 10453 -20099 10463 -20039
rect 10383 -20109 10463 -20099
rect 10063 -20379 10123 -20109
rect 10393 -20119 10463 -20109
rect 10203 -20169 10233 -20149
rect 10183 -20209 10233 -20169
rect 10293 -20169 10323 -20149
rect 10293 -20209 10343 -20169
rect 10183 -20279 10343 -20209
rect 10183 -20319 10233 -20279
rect 10203 -20339 10233 -20319
rect 10293 -20319 10343 -20279
rect 10293 -20339 10323 -20319
rect 10403 -20379 10463 -20119
rect 10063 -20389 10143 -20379
rect 10063 -20449 10073 -20389
rect 10133 -20399 10143 -20389
rect 10383 -20389 10463 -20379
rect 10383 -20399 10393 -20389
rect 10133 -20449 10393 -20399
rect 10453 -20449 10463 -20389
rect 10063 -20459 10463 -20449
rect 10521 -20039 10921 -20029
rect 10521 -20099 10531 -20039
rect 10591 -20089 10851 -20039
rect 10591 -20099 10601 -20089
rect 10521 -20109 10601 -20099
rect 10841 -20099 10851 -20089
rect 10911 -20099 10921 -20039
rect 10841 -20109 10921 -20099
rect 10521 -20379 10581 -20109
rect 10851 -20119 10921 -20109
rect 10661 -20169 10691 -20149
rect 10641 -20209 10691 -20169
rect 10751 -20169 10781 -20149
rect 10751 -20209 10801 -20169
rect 10641 -20279 10801 -20209
rect 10641 -20319 10691 -20279
rect 10661 -20339 10691 -20319
rect 10751 -20319 10801 -20279
rect 10751 -20339 10781 -20319
rect 10861 -20379 10921 -20119
rect 10521 -20389 10601 -20379
rect 10521 -20449 10531 -20389
rect 10591 -20399 10601 -20389
rect 10841 -20389 10921 -20379
rect 10841 -20399 10851 -20389
rect 10591 -20449 10851 -20399
rect 10911 -20449 10921 -20389
rect 10521 -20459 10921 -20449
rect 10977 -20039 11377 -20029
rect 10977 -20099 10987 -20039
rect 11047 -20089 11307 -20039
rect 11047 -20099 11057 -20089
rect 10977 -20109 11057 -20099
rect 11297 -20099 11307 -20089
rect 11367 -20099 11377 -20039
rect 11297 -20109 11377 -20099
rect 10977 -20379 11037 -20109
rect 11307 -20119 11377 -20109
rect 11117 -20169 11147 -20149
rect 11097 -20209 11147 -20169
rect 11207 -20169 11237 -20149
rect 11207 -20209 11257 -20169
rect 11097 -20279 11257 -20209
rect 11097 -20319 11147 -20279
rect 11117 -20339 11147 -20319
rect 11207 -20319 11257 -20279
rect 11207 -20339 11237 -20319
rect 11317 -20379 11377 -20119
rect 10977 -20389 11057 -20379
rect 10977 -20449 10987 -20389
rect 11047 -20399 11057 -20389
rect 11297 -20389 11377 -20379
rect 11297 -20399 11307 -20389
rect 11047 -20449 11307 -20399
rect 11367 -20449 11377 -20389
rect 10977 -20459 11377 -20449
rect 11433 -20039 11833 -20029
rect 11433 -20099 11443 -20039
rect 11503 -20089 11763 -20039
rect 11503 -20099 11513 -20089
rect 11433 -20109 11513 -20099
rect 11753 -20099 11763 -20089
rect 11823 -20099 11833 -20039
rect 11753 -20109 11833 -20099
rect 11433 -20379 11493 -20109
rect 11763 -20119 11833 -20109
rect 11573 -20169 11603 -20149
rect 11553 -20209 11603 -20169
rect 11663 -20169 11693 -20149
rect 11663 -20209 11713 -20169
rect 11553 -20279 11713 -20209
rect 11553 -20319 11603 -20279
rect 11573 -20339 11603 -20319
rect 11663 -20319 11713 -20279
rect 11663 -20339 11693 -20319
rect 11773 -20379 11833 -20119
rect 11433 -20389 11513 -20379
rect 11433 -20449 11443 -20389
rect 11503 -20399 11513 -20389
rect 11753 -20389 11833 -20379
rect 11753 -20399 11763 -20389
rect 11503 -20449 11763 -20399
rect 11823 -20449 11833 -20389
rect 11433 -20459 11833 -20449
rect 11891 -20039 12291 -20029
rect 11891 -20099 11901 -20039
rect 11961 -20089 12221 -20039
rect 11961 -20099 11971 -20089
rect 11891 -20109 11971 -20099
rect 12211 -20099 12221 -20089
rect 12281 -20099 12291 -20039
rect 12211 -20109 12291 -20099
rect 11891 -20379 11951 -20109
rect 12221 -20119 12291 -20109
rect 12031 -20169 12061 -20149
rect 12011 -20209 12061 -20169
rect 12121 -20169 12151 -20149
rect 12121 -20209 12171 -20169
rect 12011 -20279 12171 -20209
rect 12011 -20319 12061 -20279
rect 12031 -20339 12061 -20319
rect 12121 -20319 12171 -20279
rect 12121 -20339 12151 -20319
rect 12231 -20379 12291 -20119
rect 11891 -20389 11971 -20379
rect 11891 -20449 11901 -20389
rect 11961 -20399 11971 -20389
rect 12211 -20389 12291 -20379
rect 12211 -20399 12221 -20389
rect 11961 -20449 12221 -20399
rect 12281 -20449 12291 -20389
rect 11891 -20459 12291 -20449
rect 12347 -20039 12747 -20029
rect 12347 -20099 12357 -20039
rect 12417 -20089 12677 -20039
rect 12417 -20099 12427 -20089
rect 12347 -20109 12427 -20099
rect 12667 -20099 12677 -20089
rect 12737 -20099 12747 -20039
rect 12667 -20109 12747 -20099
rect 12347 -20379 12407 -20109
rect 12677 -20119 12747 -20109
rect 12487 -20169 12517 -20149
rect 12467 -20209 12517 -20169
rect 12577 -20169 12607 -20149
rect 12577 -20209 12627 -20169
rect 12467 -20279 12627 -20209
rect 12467 -20319 12517 -20279
rect 12487 -20339 12517 -20319
rect 12577 -20319 12627 -20279
rect 12577 -20339 12607 -20319
rect 12687 -20379 12747 -20119
rect 12347 -20389 12427 -20379
rect 12347 -20449 12357 -20389
rect 12417 -20399 12427 -20389
rect 12667 -20389 12747 -20379
rect 12667 -20399 12677 -20389
rect 12417 -20449 12677 -20399
rect 12737 -20449 12747 -20389
rect 12347 -20459 12747 -20449
rect 12803 -20039 13203 -20029
rect 12803 -20099 12813 -20039
rect 12873 -20089 13133 -20039
rect 12873 -20099 12883 -20089
rect 12803 -20109 12883 -20099
rect 13123 -20099 13133 -20089
rect 13193 -20099 13203 -20039
rect 13123 -20109 13203 -20099
rect 12803 -20379 12863 -20109
rect 13133 -20119 13203 -20109
rect 12943 -20169 12973 -20149
rect 12923 -20209 12973 -20169
rect 13033 -20169 13063 -20149
rect 13033 -20209 13083 -20169
rect 12923 -20279 13083 -20209
rect 12923 -20319 12973 -20279
rect 12943 -20339 12973 -20319
rect 13033 -20319 13083 -20279
rect 13033 -20339 13063 -20319
rect 13143 -20379 13203 -20119
rect 12803 -20389 12883 -20379
rect 12803 -20449 12813 -20389
rect 12873 -20399 12883 -20389
rect 13123 -20389 13203 -20379
rect 13123 -20399 13133 -20389
rect 12873 -20449 13133 -20399
rect 13193 -20449 13203 -20389
rect 12803 -20459 13203 -20449
rect 13261 -20039 13661 -20029
rect 13261 -20099 13271 -20039
rect 13331 -20089 13591 -20039
rect 13331 -20099 13341 -20089
rect 13261 -20109 13341 -20099
rect 13581 -20099 13591 -20089
rect 13651 -20099 13661 -20039
rect 13581 -20109 13661 -20099
rect 13261 -20379 13321 -20109
rect 13591 -20119 13661 -20109
rect 13401 -20169 13431 -20149
rect 13381 -20209 13431 -20169
rect 13491 -20169 13521 -20149
rect 13491 -20209 13541 -20169
rect 13381 -20279 13541 -20209
rect 13381 -20319 13431 -20279
rect 13401 -20339 13431 -20319
rect 13491 -20319 13541 -20279
rect 13491 -20339 13521 -20319
rect 13601 -20379 13661 -20119
rect 13261 -20389 13341 -20379
rect 13261 -20449 13271 -20389
rect 13331 -20399 13341 -20389
rect 13581 -20389 13661 -20379
rect 13581 -20399 13591 -20389
rect 13331 -20449 13591 -20399
rect 13651 -20449 13661 -20389
rect 13261 -20459 13661 -20449
rect 13717 -20039 14117 -20029
rect 13717 -20099 13727 -20039
rect 13787 -20089 14047 -20039
rect 13787 -20099 13797 -20089
rect 13717 -20109 13797 -20099
rect 14037 -20099 14047 -20089
rect 14107 -20099 14117 -20039
rect 14037 -20109 14117 -20099
rect 13717 -20379 13777 -20109
rect 14047 -20119 14117 -20109
rect 13857 -20169 13887 -20149
rect 13837 -20209 13887 -20169
rect 13947 -20169 13977 -20149
rect 13947 -20209 13997 -20169
rect 13837 -20279 13997 -20209
rect 13837 -20319 13887 -20279
rect 13857 -20339 13887 -20319
rect 13947 -20319 13997 -20279
rect 13947 -20339 13977 -20319
rect 14057 -20379 14117 -20119
rect 13717 -20389 13797 -20379
rect 13717 -20449 13727 -20389
rect 13787 -20399 13797 -20389
rect 14037 -20389 14117 -20379
rect 14037 -20399 14047 -20389
rect 13787 -20449 14047 -20399
rect 14107 -20449 14117 -20389
rect 13717 -20459 14117 -20449
rect 14173 -20039 14573 -20029
rect 14173 -20099 14183 -20039
rect 14243 -20089 14503 -20039
rect 14243 -20099 14253 -20089
rect 14173 -20109 14253 -20099
rect 14493 -20099 14503 -20089
rect 14563 -20099 14573 -20039
rect 14493 -20109 14573 -20099
rect 14173 -20379 14233 -20109
rect 14503 -20119 14573 -20109
rect 14313 -20169 14343 -20149
rect 14293 -20209 14343 -20169
rect 14403 -20169 14433 -20149
rect 14403 -20209 14453 -20169
rect 14293 -20279 14453 -20209
rect 14293 -20319 14343 -20279
rect 14313 -20339 14343 -20319
rect 14403 -20319 14453 -20279
rect 14403 -20339 14433 -20319
rect 14513 -20379 14573 -20119
rect 14173 -20389 14253 -20379
rect 14173 -20449 14183 -20389
rect 14243 -20399 14253 -20389
rect 14493 -20389 14573 -20379
rect 14493 -20399 14503 -20389
rect 14243 -20449 14503 -20399
rect 14563 -20449 14573 -20389
rect 14173 -20459 14573 -20449
rect 14631 -20039 15031 -20029
rect 14631 -20099 14641 -20039
rect 14701 -20089 14961 -20039
rect 14701 -20099 14711 -20089
rect 14631 -20109 14711 -20099
rect 14951 -20099 14961 -20089
rect 15021 -20099 15031 -20039
rect 14951 -20109 15031 -20099
rect 14631 -20379 14691 -20109
rect 14961 -20119 15031 -20109
rect 14771 -20169 14801 -20149
rect 14751 -20209 14801 -20169
rect 14861 -20169 14891 -20149
rect 14861 -20209 14911 -20169
rect 14751 -20279 14911 -20209
rect 14751 -20319 14801 -20279
rect 14771 -20339 14801 -20319
rect 14861 -20319 14911 -20279
rect 14861 -20339 14891 -20319
rect 14971 -20379 15031 -20119
rect 14631 -20389 14711 -20379
rect 14631 -20449 14641 -20389
rect 14701 -20399 14711 -20389
rect 14951 -20389 15031 -20379
rect 14951 -20399 14961 -20389
rect 14701 -20449 14961 -20399
rect 15021 -20449 15031 -20389
rect 14631 -20459 15031 -20449
rect 15087 -20039 15487 -20029
rect 15087 -20099 15097 -20039
rect 15157 -20089 15417 -20039
rect 15157 -20099 15167 -20089
rect 15087 -20109 15167 -20099
rect 15407 -20099 15417 -20089
rect 15477 -20099 15487 -20039
rect 15407 -20109 15487 -20099
rect 15087 -20379 15147 -20109
rect 15417 -20119 15487 -20109
rect 15227 -20169 15257 -20149
rect 15207 -20209 15257 -20169
rect 15317 -20169 15347 -20149
rect 15317 -20209 15367 -20169
rect 15207 -20279 15367 -20209
rect 15207 -20319 15257 -20279
rect 15227 -20339 15257 -20319
rect 15317 -20319 15367 -20279
rect 15317 -20339 15347 -20319
rect 15427 -20379 15487 -20119
rect 15087 -20389 15167 -20379
rect 15087 -20449 15097 -20389
rect 15157 -20399 15167 -20389
rect 15407 -20389 15487 -20379
rect 15407 -20399 15417 -20389
rect 15157 -20449 15417 -20399
rect 15477 -20449 15487 -20389
rect 15087 -20459 15487 -20449
rect 1 -20531 401 -20521
rect 1 -20591 11 -20531
rect 71 -20581 331 -20531
rect 71 -20591 81 -20581
rect 1 -20601 81 -20591
rect 321 -20591 331 -20581
rect 391 -20591 401 -20531
rect 321 -20601 401 -20591
rect 1 -20871 61 -20601
rect 331 -20611 401 -20601
rect 141 -20661 171 -20641
rect 121 -20701 171 -20661
rect 231 -20661 261 -20641
rect 231 -20701 281 -20661
rect 121 -20771 281 -20701
rect 121 -20811 171 -20771
rect 141 -20831 171 -20811
rect 231 -20811 281 -20771
rect 231 -20831 261 -20811
rect 341 -20871 401 -20611
rect 1 -20881 81 -20871
rect 1 -20941 11 -20881
rect 71 -20891 81 -20881
rect 321 -20881 401 -20871
rect 321 -20891 331 -20881
rect 71 -20941 331 -20891
rect 391 -20941 401 -20881
rect 1 -20951 401 -20941
rect 457 -20531 857 -20521
rect 457 -20591 467 -20531
rect 527 -20581 787 -20531
rect 527 -20591 537 -20581
rect 457 -20601 537 -20591
rect 777 -20591 787 -20581
rect 847 -20591 857 -20531
rect 777 -20601 857 -20591
rect 457 -20871 517 -20601
rect 787 -20611 857 -20601
rect 597 -20661 627 -20641
rect 577 -20701 627 -20661
rect 687 -20661 717 -20641
rect 687 -20701 737 -20661
rect 577 -20771 737 -20701
rect 577 -20811 627 -20771
rect 597 -20831 627 -20811
rect 687 -20811 737 -20771
rect 687 -20831 717 -20811
rect 797 -20871 857 -20611
rect 457 -20881 537 -20871
rect 457 -20941 467 -20881
rect 527 -20891 537 -20881
rect 777 -20881 857 -20871
rect 777 -20891 787 -20881
rect 527 -20941 787 -20891
rect 847 -20941 857 -20881
rect 457 -20951 857 -20941
rect 913 -20531 1313 -20521
rect 913 -20591 923 -20531
rect 983 -20581 1243 -20531
rect 983 -20591 993 -20581
rect 913 -20601 993 -20591
rect 1233 -20591 1243 -20581
rect 1303 -20591 1313 -20531
rect 1233 -20601 1313 -20591
rect 913 -20871 973 -20601
rect 1243 -20611 1313 -20601
rect 1053 -20661 1083 -20641
rect 1033 -20701 1083 -20661
rect 1143 -20661 1173 -20641
rect 1143 -20701 1193 -20661
rect 1033 -20771 1193 -20701
rect 1033 -20811 1083 -20771
rect 1053 -20831 1083 -20811
rect 1143 -20811 1193 -20771
rect 1143 -20831 1173 -20811
rect 1253 -20871 1313 -20611
rect 913 -20881 993 -20871
rect 913 -20941 923 -20881
rect 983 -20891 993 -20881
rect 1233 -20881 1313 -20871
rect 1233 -20891 1243 -20881
rect 983 -20941 1243 -20891
rect 1303 -20941 1313 -20881
rect 913 -20951 1313 -20941
rect 1371 -20531 1771 -20521
rect 1371 -20591 1381 -20531
rect 1441 -20581 1701 -20531
rect 1441 -20591 1451 -20581
rect 1371 -20601 1451 -20591
rect 1691 -20591 1701 -20581
rect 1761 -20591 1771 -20531
rect 1691 -20601 1771 -20591
rect 1371 -20871 1431 -20601
rect 1701 -20611 1771 -20601
rect 1511 -20661 1541 -20641
rect 1491 -20701 1541 -20661
rect 1601 -20661 1631 -20641
rect 1601 -20701 1651 -20661
rect 1491 -20771 1651 -20701
rect 1491 -20811 1541 -20771
rect 1511 -20831 1541 -20811
rect 1601 -20811 1651 -20771
rect 1601 -20831 1631 -20811
rect 1711 -20871 1771 -20611
rect 1371 -20881 1451 -20871
rect 1371 -20941 1381 -20881
rect 1441 -20891 1451 -20881
rect 1691 -20881 1771 -20871
rect 1691 -20891 1701 -20881
rect 1441 -20941 1701 -20891
rect 1761 -20941 1771 -20881
rect 1371 -20951 1771 -20941
rect 1827 -20531 2227 -20521
rect 1827 -20591 1837 -20531
rect 1897 -20581 2157 -20531
rect 1897 -20591 1907 -20581
rect 1827 -20601 1907 -20591
rect 2147 -20591 2157 -20581
rect 2217 -20591 2227 -20531
rect 2147 -20601 2227 -20591
rect 1827 -20871 1887 -20601
rect 2157 -20611 2227 -20601
rect 1967 -20661 1997 -20641
rect 1947 -20701 1997 -20661
rect 2057 -20661 2087 -20641
rect 2057 -20701 2107 -20661
rect 1947 -20771 2107 -20701
rect 1947 -20811 1997 -20771
rect 1967 -20831 1997 -20811
rect 2057 -20811 2107 -20771
rect 2057 -20831 2087 -20811
rect 2167 -20871 2227 -20611
rect 1827 -20881 1907 -20871
rect 1827 -20941 1837 -20881
rect 1897 -20891 1907 -20881
rect 2147 -20881 2227 -20871
rect 2147 -20891 2157 -20881
rect 1897 -20941 2157 -20891
rect 2217 -20941 2227 -20881
rect 1827 -20951 2227 -20941
rect 2283 -20531 2683 -20521
rect 2283 -20591 2293 -20531
rect 2353 -20581 2613 -20531
rect 2353 -20591 2363 -20581
rect 2283 -20601 2363 -20591
rect 2603 -20591 2613 -20581
rect 2673 -20591 2683 -20531
rect 2603 -20601 2683 -20591
rect 2283 -20871 2343 -20601
rect 2613 -20611 2683 -20601
rect 2423 -20661 2453 -20641
rect 2403 -20701 2453 -20661
rect 2513 -20661 2543 -20641
rect 2513 -20701 2563 -20661
rect 2403 -20771 2563 -20701
rect 2403 -20811 2453 -20771
rect 2423 -20831 2453 -20811
rect 2513 -20811 2563 -20771
rect 2513 -20831 2543 -20811
rect 2623 -20871 2683 -20611
rect 2283 -20881 2363 -20871
rect 2283 -20941 2293 -20881
rect 2353 -20891 2363 -20881
rect 2603 -20881 2683 -20871
rect 2603 -20891 2613 -20881
rect 2353 -20941 2613 -20891
rect 2673 -20941 2683 -20881
rect 2283 -20951 2683 -20941
rect 2741 -20531 3141 -20521
rect 2741 -20591 2751 -20531
rect 2811 -20581 3071 -20531
rect 2811 -20591 2821 -20581
rect 2741 -20601 2821 -20591
rect 3061 -20591 3071 -20581
rect 3131 -20591 3141 -20531
rect 3061 -20601 3141 -20591
rect 2741 -20871 2801 -20601
rect 3071 -20611 3141 -20601
rect 2881 -20661 2911 -20641
rect 2861 -20701 2911 -20661
rect 2971 -20661 3001 -20641
rect 2971 -20701 3021 -20661
rect 2861 -20771 3021 -20701
rect 2861 -20811 2911 -20771
rect 2881 -20831 2911 -20811
rect 2971 -20811 3021 -20771
rect 2971 -20831 3001 -20811
rect 3081 -20871 3141 -20611
rect 2741 -20881 2821 -20871
rect 2741 -20941 2751 -20881
rect 2811 -20891 2821 -20881
rect 3061 -20881 3141 -20871
rect 3061 -20891 3071 -20881
rect 2811 -20941 3071 -20891
rect 3131 -20941 3141 -20881
rect 2741 -20951 3141 -20941
rect 3197 -20531 3597 -20521
rect 3197 -20591 3207 -20531
rect 3267 -20581 3527 -20531
rect 3267 -20591 3277 -20581
rect 3197 -20601 3277 -20591
rect 3517 -20591 3527 -20581
rect 3587 -20591 3597 -20531
rect 3517 -20601 3597 -20591
rect 3197 -20871 3257 -20601
rect 3527 -20611 3597 -20601
rect 3337 -20661 3367 -20641
rect 3317 -20701 3367 -20661
rect 3427 -20661 3457 -20641
rect 3427 -20701 3477 -20661
rect 3317 -20771 3477 -20701
rect 3317 -20811 3367 -20771
rect 3337 -20831 3367 -20811
rect 3427 -20811 3477 -20771
rect 3427 -20831 3457 -20811
rect 3537 -20871 3597 -20611
rect 3197 -20881 3277 -20871
rect 3197 -20941 3207 -20881
rect 3267 -20891 3277 -20881
rect 3517 -20881 3597 -20871
rect 3517 -20891 3527 -20881
rect 3267 -20941 3527 -20891
rect 3587 -20941 3597 -20881
rect 3197 -20951 3597 -20941
rect 3653 -20531 4053 -20521
rect 3653 -20591 3663 -20531
rect 3723 -20581 3983 -20531
rect 3723 -20591 3733 -20581
rect 3653 -20601 3733 -20591
rect 3973 -20591 3983 -20581
rect 4043 -20591 4053 -20531
rect 3973 -20601 4053 -20591
rect 3653 -20871 3713 -20601
rect 3983 -20611 4053 -20601
rect 3793 -20661 3823 -20641
rect 3773 -20701 3823 -20661
rect 3883 -20661 3913 -20641
rect 3883 -20701 3933 -20661
rect 3773 -20771 3933 -20701
rect 3773 -20811 3823 -20771
rect 3793 -20831 3823 -20811
rect 3883 -20811 3933 -20771
rect 3883 -20831 3913 -20811
rect 3993 -20871 4053 -20611
rect 3653 -20881 3733 -20871
rect 3653 -20941 3663 -20881
rect 3723 -20891 3733 -20881
rect 3973 -20881 4053 -20871
rect 3973 -20891 3983 -20881
rect 3723 -20941 3983 -20891
rect 4043 -20941 4053 -20881
rect 3653 -20951 4053 -20941
rect 4111 -20531 4511 -20521
rect 4111 -20591 4121 -20531
rect 4181 -20581 4441 -20531
rect 4181 -20591 4191 -20581
rect 4111 -20601 4191 -20591
rect 4431 -20591 4441 -20581
rect 4501 -20591 4511 -20531
rect 4431 -20601 4511 -20591
rect 4111 -20871 4171 -20601
rect 4441 -20611 4511 -20601
rect 4251 -20661 4281 -20641
rect 4231 -20701 4281 -20661
rect 4341 -20661 4371 -20641
rect 4341 -20701 4391 -20661
rect 4231 -20771 4391 -20701
rect 4231 -20811 4281 -20771
rect 4251 -20831 4281 -20811
rect 4341 -20811 4391 -20771
rect 4341 -20831 4371 -20811
rect 4451 -20871 4511 -20611
rect 4111 -20881 4191 -20871
rect 4111 -20941 4121 -20881
rect 4181 -20891 4191 -20881
rect 4431 -20881 4511 -20871
rect 4431 -20891 4441 -20881
rect 4181 -20941 4441 -20891
rect 4501 -20941 4511 -20881
rect 4111 -20951 4511 -20941
rect 4567 -20531 4967 -20521
rect 4567 -20591 4577 -20531
rect 4637 -20581 4897 -20531
rect 4637 -20591 4647 -20581
rect 4567 -20601 4647 -20591
rect 4887 -20591 4897 -20581
rect 4957 -20591 4967 -20531
rect 4887 -20601 4967 -20591
rect 4567 -20871 4627 -20601
rect 4897 -20611 4967 -20601
rect 4707 -20661 4737 -20641
rect 4687 -20701 4737 -20661
rect 4797 -20661 4827 -20641
rect 4797 -20701 4847 -20661
rect 4687 -20771 4847 -20701
rect 4687 -20811 4737 -20771
rect 4707 -20831 4737 -20811
rect 4797 -20811 4847 -20771
rect 4797 -20831 4827 -20811
rect 4907 -20871 4967 -20611
rect 4567 -20881 4647 -20871
rect 4567 -20941 4577 -20881
rect 4637 -20891 4647 -20881
rect 4887 -20881 4967 -20871
rect 4887 -20891 4897 -20881
rect 4637 -20941 4897 -20891
rect 4957 -20941 4967 -20881
rect 4567 -20951 4967 -20941
rect 5023 -20531 5423 -20521
rect 5023 -20591 5033 -20531
rect 5093 -20581 5353 -20531
rect 5093 -20591 5103 -20581
rect 5023 -20601 5103 -20591
rect 5343 -20591 5353 -20581
rect 5413 -20591 5423 -20531
rect 5343 -20601 5423 -20591
rect 5023 -20871 5083 -20601
rect 5353 -20611 5423 -20601
rect 5163 -20661 5193 -20641
rect 5143 -20701 5193 -20661
rect 5253 -20661 5283 -20641
rect 5253 -20701 5303 -20661
rect 5143 -20771 5303 -20701
rect 5143 -20811 5193 -20771
rect 5163 -20831 5193 -20811
rect 5253 -20811 5303 -20771
rect 5253 -20831 5283 -20811
rect 5363 -20871 5423 -20611
rect 5023 -20881 5103 -20871
rect 5023 -20941 5033 -20881
rect 5093 -20891 5103 -20881
rect 5343 -20881 5423 -20871
rect 5343 -20891 5353 -20881
rect 5093 -20941 5353 -20891
rect 5413 -20941 5423 -20881
rect 5023 -20951 5423 -20941
rect 5481 -20531 5881 -20521
rect 5481 -20591 5491 -20531
rect 5551 -20581 5811 -20531
rect 5551 -20591 5561 -20581
rect 5481 -20601 5561 -20591
rect 5801 -20591 5811 -20581
rect 5871 -20591 5881 -20531
rect 5801 -20601 5881 -20591
rect 5481 -20871 5541 -20601
rect 5811 -20611 5881 -20601
rect 5621 -20661 5651 -20641
rect 5601 -20701 5651 -20661
rect 5711 -20661 5741 -20641
rect 5711 -20701 5761 -20661
rect 5601 -20771 5761 -20701
rect 5601 -20811 5651 -20771
rect 5621 -20831 5651 -20811
rect 5711 -20811 5761 -20771
rect 5711 -20831 5741 -20811
rect 5821 -20871 5881 -20611
rect 5481 -20881 5561 -20871
rect 5481 -20941 5491 -20881
rect 5551 -20891 5561 -20881
rect 5801 -20881 5881 -20871
rect 5801 -20891 5811 -20881
rect 5551 -20941 5811 -20891
rect 5871 -20941 5881 -20881
rect 5481 -20951 5881 -20941
rect 5937 -20531 6337 -20521
rect 5937 -20591 5947 -20531
rect 6007 -20581 6267 -20531
rect 6007 -20591 6017 -20581
rect 5937 -20601 6017 -20591
rect 6257 -20591 6267 -20581
rect 6327 -20591 6337 -20531
rect 6257 -20601 6337 -20591
rect 5937 -20871 5997 -20601
rect 6267 -20611 6337 -20601
rect 6077 -20661 6107 -20641
rect 6057 -20701 6107 -20661
rect 6167 -20661 6197 -20641
rect 6167 -20701 6217 -20661
rect 6057 -20771 6217 -20701
rect 6057 -20811 6107 -20771
rect 6077 -20831 6107 -20811
rect 6167 -20811 6217 -20771
rect 6167 -20831 6197 -20811
rect 6277 -20871 6337 -20611
rect 5937 -20881 6017 -20871
rect 5937 -20941 5947 -20881
rect 6007 -20891 6017 -20881
rect 6257 -20881 6337 -20871
rect 6257 -20891 6267 -20881
rect 6007 -20941 6267 -20891
rect 6327 -20941 6337 -20881
rect 5937 -20951 6337 -20941
rect 6393 -20531 6793 -20521
rect 6393 -20591 6403 -20531
rect 6463 -20581 6723 -20531
rect 6463 -20591 6473 -20581
rect 6393 -20601 6473 -20591
rect 6713 -20591 6723 -20581
rect 6783 -20591 6793 -20531
rect 6713 -20601 6793 -20591
rect 6393 -20871 6453 -20601
rect 6723 -20611 6793 -20601
rect 6533 -20661 6563 -20641
rect 6513 -20701 6563 -20661
rect 6623 -20661 6653 -20641
rect 6623 -20701 6673 -20661
rect 6513 -20771 6673 -20701
rect 6513 -20811 6563 -20771
rect 6533 -20831 6563 -20811
rect 6623 -20811 6673 -20771
rect 6623 -20831 6653 -20811
rect 6733 -20871 6793 -20611
rect 6393 -20881 6473 -20871
rect 6393 -20941 6403 -20881
rect 6463 -20891 6473 -20881
rect 6713 -20881 6793 -20871
rect 6713 -20891 6723 -20881
rect 6463 -20941 6723 -20891
rect 6783 -20941 6793 -20881
rect 6393 -20951 6793 -20941
rect 6851 -20531 7251 -20521
rect 6851 -20591 6861 -20531
rect 6921 -20581 7181 -20531
rect 6921 -20591 6931 -20581
rect 6851 -20601 6931 -20591
rect 7171 -20591 7181 -20581
rect 7241 -20591 7251 -20531
rect 7171 -20601 7251 -20591
rect 6851 -20871 6911 -20601
rect 7181 -20611 7251 -20601
rect 6991 -20661 7021 -20641
rect 6971 -20701 7021 -20661
rect 7081 -20661 7111 -20641
rect 7081 -20701 7131 -20661
rect 6971 -20771 7131 -20701
rect 6971 -20811 7021 -20771
rect 6991 -20831 7021 -20811
rect 7081 -20811 7131 -20771
rect 7081 -20831 7111 -20811
rect 7191 -20871 7251 -20611
rect 6851 -20881 6931 -20871
rect 6851 -20941 6861 -20881
rect 6921 -20891 6931 -20881
rect 7171 -20881 7251 -20871
rect 7171 -20891 7181 -20881
rect 6921 -20941 7181 -20891
rect 7241 -20941 7251 -20881
rect 6851 -20951 7251 -20941
rect 7307 -20531 7707 -20521
rect 7307 -20591 7317 -20531
rect 7377 -20581 7637 -20531
rect 7377 -20591 7387 -20581
rect 7307 -20601 7387 -20591
rect 7627 -20591 7637 -20581
rect 7697 -20591 7707 -20531
rect 7627 -20601 7707 -20591
rect 7307 -20871 7367 -20601
rect 7637 -20611 7707 -20601
rect 7447 -20661 7477 -20641
rect 7427 -20701 7477 -20661
rect 7537 -20661 7567 -20641
rect 7537 -20701 7587 -20661
rect 7427 -20771 7587 -20701
rect 7427 -20811 7477 -20771
rect 7447 -20831 7477 -20811
rect 7537 -20811 7587 -20771
rect 7537 -20831 7567 -20811
rect 7647 -20871 7707 -20611
rect 7307 -20881 7387 -20871
rect 7307 -20941 7317 -20881
rect 7377 -20891 7387 -20881
rect 7627 -20881 7707 -20871
rect 7627 -20891 7637 -20881
rect 7377 -20941 7637 -20891
rect 7697 -20941 7707 -20881
rect 7307 -20951 7707 -20941
rect 7763 -20531 8163 -20521
rect 7763 -20591 7773 -20531
rect 7833 -20581 8093 -20531
rect 7833 -20591 7843 -20581
rect 7763 -20601 7843 -20591
rect 8083 -20591 8093 -20581
rect 8153 -20591 8163 -20531
rect 8083 -20601 8163 -20591
rect 7763 -20871 7823 -20601
rect 8093 -20611 8163 -20601
rect 7903 -20661 7933 -20641
rect 7883 -20701 7933 -20661
rect 7993 -20661 8023 -20641
rect 7993 -20701 8043 -20661
rect 7883 -20771 8043 -20701
rect 7883 -20811 7933 -20771
rect 7903 -20831 7933 -20811
rect 7993 -20811 8043 -20771
rect 7993 -20831 8023 -20811
rect 8103 -20871 8163 -20611
rect 7763 -20881 7843 -20871
rect 7763 -20941 7773 -20881
rect 7833 -20891 7843 -20881
rect 8083 -20881 8163 -20871
rect 8083 -20891 8093 -20881
rect 7833 -20941 8093 -20891
rect 8153 -20941 8163 -20881
rect 7763 -20951 8163 -20941
rect 8237 -20531 8637 -20521
rect 8237 -20591 8247 -20531
rect 8307 -20581 8567 -20531
rect 8307 -20591 8317 -20581
rect 8237 -20601 8317 -20591
rect 8557 -20591 8567 -20581
rect 8627 -20591 8637 -20531
rect 8557 -20601 8637 -20591
rect 8237 -20871 8297 -20601
rect 8567 -20611 8637 -20601
rect 8377 -20661 8407 -20641
rect 8357 -20701 8407 -20661
rect 8467 -20661 8497 -20641
rect 8467 -20701 8517 -20661
rect 8357 -20771 8517 -20701
rect 8357 -20811 8407 -20771
rect 8377 -20831 8407 -20811
rect 8467 -20811 8517 -20771
rect 8467 -20831 8497 -20811
rect 8577 -20871 8637 -20611
rect 8237 -20881 8317 -20871
rect 8237 -20941 8247 -20881
rect 8307 -20891 8317 -20881
rect 8557 -20881 8637 -20871
rect 8557 -20891 8567 -20881
rect 8307 -20941 8567 -20891
rect 8627 -20941 8637 -20881
rect 8237 -20951 8637 -20941
rect 8693 -20531 9093 -20521
rect 8693 -20591 8703 -20531
rect 8763 -20581 9023 -20531
rect 8763 -20591 8773 -20581
rect 8693 -20601 8773 -20591
rect 9013 -20591 9023 -20581
rect 9083 -20591 9093 -20531
rect 9013 -20601 9093 -20591
rect 8693 -20871 8753 -20601
rect 9023 -20611 9093 -20601
rect 8833 -20661 8863 -20641
rect 8813 -20701 8863 -20661
rect 8923 -20661 8953 -20641
rect 8923 -20701 8973 -20661
rect 8813 -20771 8973 -20701
rect 8813 -20811 8863 -20771
rect 8833 -20831 8863 -20811
rect 8923 -20811 8973 -20771
rect 8923 -20831 8953 -20811
rect 9033 -20871 9093 -20611
rect 8693 -20881 8773 -20871
rect 8693 -20941 8703 -20881
rect 8763 -20891 8773 -20881
rect 9013 -20881 9093 -20871
rect 9013 -20891 9023 -20881
rect 8763 -20941 9023 -20891
rect 9083 -20941 9093 -20881
rect 8693 -20951 9093 -20941
rect 9151 -20531 9551 -20521
rect 9151 -20591 9161 -20531
rect 9221 -20581 9481 -20531
rect 9221 -20591 9231 -20581
rect 9151 -20601 9231 -20591
rect 9471 -20591 9481 -20581
rect 9541 -20591 9551 -20531
rect 9471 -20601 9551 -20591
rect 9151 -20871 9211 -20601
rect 9481 -20611 9551 -20601
rect 9291 -20661 9321 -20641
rect 9271 -20701 9321 -20661
rect 9381 -20661 9411 -20641
rect 9381 -20701 9431 -20661
rect 9271 -20771 9431 -20701
rect 9271 -20811 9321 -20771
rect 9291 -20831 9321 -20811
rect 9381 -20811 9431 -20771
rect 9381 -20831 9411 -20811
rect 9491 -20871 9551 -20611
rect 9151 -20881 9231 -20871
rect 9151 -20941 9161 -20881
rect 9221 -20891 9231 -20881
rect 9471 -20881 9551 -20871
rect 9471 -20891 9481 -20881
rect 9221 -20941 9481 -20891
rect 9541 -20941 9551 -20881
rect 9151 -20951 9551 -20941
rect 9607 -20531 10007 -20521
rect 9607 -20591 9617 -20531
rect 9677 -20581 9937 -20531
rect 9677 -20591 9687 -20581
rect 9607 -20601 9687 -20591
rect 9927 -20591 9937 -20581
rect 9997 -20591 10007 -20531
rect 9927 -20601 10007 -20591
rect 9607 -20871 9667 -20601
rect 9937 -20611 10007 -20601
rect 9747 -20661 9777 -20641
rect 9727 -20701 9777 -20661
rect 9837 -20661 9867 -20641
rect 9837 -20701 9887 -20661
rect 9727 -20771 9887 -20701
rect 9727 -20811 9777 -20771
rect 9747 -20831 9777 -20811
rect 9837 -20811 9887 -20771
rect 9837 -20831 9867 -20811
rect 9947 -20871 10007 -20611
rect 9607 -20881 9687 -20871
rect 9607 -20941 9617 -20881
rect 9677 -20891 9687 -20881
rect 9927 -20881 10007 -20871
rect 9927 -20891 9937 -20881
rect 9677 -20941 9937 -20891
rect 9997 -20941 10007 -20881
rect 9607 -20951 10007 -20941
rect 10063 -20531 10463 -20521
rect 10063 -20591 10073 -20531
rect 10133 -20581 10393 -20531
rect 10133 -20591 10143 -20581
rect 10063 -20601 10143 -20591
rect 10383 -20591 10393 -20581
rect 10453 -20591 10463 -20531
rect 10383 -20601 10463 -20591
rect 10063 -20871 10123 -20601
rect 10393 -20611 10463 -20601
rect 10203 -20661 10233 -20641
rect 10183 -20701 10233 -20661
rect 10293 -20661 10323 -20641
rect 10293 -20701 10343 -20661
rect 10183 -20771 10343 -20701
rect 10183 -20811 10233 -20771
rect 10203 -20831 10233 -20811
rect 10293 -20811 10343 -20771
rect 10293 -20831 10323 -20811
rect 10403 -20871 10463 -20611
rect 10063 -20881 10143 -20871
rect 10063 -20941 10073 -20881
rect 10133 -20891 10143 -20881
rect 10383 -20881 10463 -20871
rect 10383 -20891 10393 -20881
rect 10133 -20941 10393 -20891
rect 10453 -20941 10463 -20881
rect 10063 -20951 10463 -20941
rect 10521 -20531 10921 -20521
rect 10521 -20591 10531 -20531
rect 10591 -20581 10851 -20531
rect 10591 -20591 10601 -20581
rect 10521 -20601 10601 -20591
rect 10841 -20591 10851 -20581
rect 10911 -20591 10921 -20531
rect 10841 -20601 10921 -20591
rect 10521 -20871 10581 -20601
rect 10851 -20611 10921 -20601
rect 10661 -20661 10691 -20641
rect 10641 -20701 10691 -20661
rect 10751 -20661 10781 -20641
rect 10751 -20701 10801 -20661
rect 10641 -20771 10801 -20701
rect 10641 -20811 10691 -20771
rect 10661 -20831 10691 -20811
rect 10751 -20811 10801 -20771
rect 10751 -20831 10781 -20811
rect 10861 -20871 10921 -20611
rect 10521 -20881 10601 -20871
rect 10521 -20941 10531 -20881
rect 10591 -20891 10601 -20881
rect 10841 -20881 10921 -20871
rect 10841 -20891 10851 -20881
rect 10591 -20941 10851 -20891
rect 10911 -20941 10921 -20881
rect 10521 -20951 10921 -20941
rect 10977 -20531 11377 -20521
rect 10977 -20591 10987 -20531
rect 11047 -20581 11307 -20531
rect 11047 -20591 11057 -20581
rect 10977 -20601 11057 -20591
rect 11297 -20591 11307 -20581
rect 11367 -20591 11377 -20531
rect 11297 -20601 11377 -20591
rect 10977 -20871 11037 -20601
rect 11307 -20611 11377 -20601
rect 11117 -20661 11147 -20641
rect 11097 -20701 11147 -20661
rect 11207 -20661 11237 -20641
rect 11207 -20701 11257 -20661
rect 11097 -20771 11257 -20701
rect 11097 -20811 11147 -20771
rect 11117 -20831 11147 -20811
rect 11207 -20811 11257 -20771
rect 11207 -20831 11237 -20811
rect 11317 -20871 11377 -20611
rect 10977 -20881 11057 -20871
rect 10977 -20941 10987 -20881
rect 11047 -20891 11057 -20881
rect 11297 -20881 11377 -20871
rect 11297 -20891 11307 -20881
rect 11047 -20941 11307 -20891
rect 11367 -20941 11377 -20881
rect 10977 -20951 11377 -20941
rect 11433 -20531 11833 -20521
rect 11433 -20591 11443 -20531
rect 11503 -20581 11763 -20531
rect 11503 -20591 11513 -20581
rect 11433 -20601 11513 -20591
rect 11753 -20591 11763 -20581
rect 11823 -20591 11833 -20531
rect 11753 -20601 11833 -20591
rect 11433 -20871 11493 -20601
rect 11763 -20611 11833 -20601
rect 11573 -20661 11603 -20641
rect 11553 -20701 11603 -20661
rect 11663 -20661 11693 -20641
rect 11663 -20701 11713 -20661
rect 11553 -20771 11713 -20701
rect 11553 -20811 11603 -20771
rect 11573 -20831 11603 -20811
rect 11663 -20811 11713 -20771
rect 11663 -20831 11693 -20811
rect 11773 -20871 11833 -20611
rect 11433 -20881 11513 -20871
rect 11433 -20941 11443 -20881
rect 11503 -20891 11513 -20881
rect 11753 -20881 11833 -20871
rect 11753 -20891 11763 -20881
rect 11503 -20941 11763 -20891
rect 11823 -20941 11833 -20881
rect 11433 -20951 11833 -20941
rect 11891 -20531 12291 -20521
rect 11891 -20591 11901 -20531
rect 11961 -20581 12221 -20531
rect 11961 -20591 11971 -20581
rect 11891 -20601 11971 -20591
rect 12211 -20591 12221 -20581
rect 12281 -20591 12291 -20531
rect 12211 -20601 12291 -20591
rect 11891 -20871 11951 -20601
rect 12221 -20611 12291 -20601
rect 12031 -20661 12061 -20641
rect 12011 -20701 12061 -20661
rect 12121 -20661 12151 -20641
rect 12121 -20701 12171 -20661
rect 12011 -20771 12171 -20701
rect 12011 -20811 12061 -20771
rect 12031 -20831 12061 -20811
rect 12121 -20811 12171 -20771
rect 12121 -20831 12151 -20811
rect 12231 -20871 12291 -20611
rect 11891 -20881 11971 -20871
rect 11891 -20941 11901 -20881
rect 11961 -20891 11971 -20881
rect 12211 -20881 12291 -20871
rect 12211 -20891 12221 -20881
rect 11961 -20941 12221 -20891
rect 12281 -20941 12291 -20881
rect 11891 -20951 12291 -20941
rect 12347 -20531 12747 -20521
rect 12347 -20591 12357 -20531
rect 12417 -20581 12677 -20531
rect 12417 -20591 12427 -20581
rect 12347 -20601 12427 -20591
rect 12667 -20591 12677 -20581
rect 12737 -20591 12747 -20531
rect 12667 -20601 12747 -20591
rect 12347 -20871 12407 -20601
rect 12677 -20611 12747 -20601
rect 12487 -20661 12517 -20641
rect 12467 -20701 12517 -20661
rect 12577 -20661 12607 -20641
rect 12577 -20701 12627 -20661
rect 12467 -20771 12627 -20701
rect 12467 -20811 12517 -20771
rect 12487 -20831 12517 -20811
rect 12577 -20811 12627 -20771
rect 12577 -20831 12607 -20811
rect 12687 -20871 12747 -20611
rect 12347 -20881 12427 -20871
rect 12347 -20941 12357 -20881
rect 12417 -20891 12427 -20881
rect 12667 -20881 12747 -20871
rect 12667 -20891 12677 -20881
rect 12417 -20941 12677 -20891
rect 12737 -20941 12747 -20881
rect 12347 -20951 12747 -20941
rect 12803 -20531 13203 -20521
rect 12803 -20591 12813 -20531
rect 12873 -20581 13133 -20531
rect 12873 -20591 12883 -20581
rect 12803 -20601 12883 -20591
rect 13123 -20591 13133 -20581
rect 13193 -20591 13203 -20531
rect 13123 -20601 13203 -20591
rect 12803 -20871 12863 -20601
rect 13133 -20611 13203 -20601
rect 12943 -20661 12973 -20641
rect 12923 -20701 12973 -20661
rect 13033 -20661 13063 -20641
rect 13033 -20701 13083 -20661
rect 12923 -20771 13083 -20701
rect 12923 -20811 12973 -20771
rect 12943 -20831 12973 -20811
rect 13033 -20811 13083 -20771
rect 13033 -20831 13063 -20811
rect 13143 -20871 13203 -20611
rect 12803 -20881 12883 -20871
rect 12803 -20941 12813 -20881
rect 12873 -20891 12883 -20881
rect 13123 -20881 13203 -20871
rect 13123 -20891 13133 -20881
rect 12873 -20941 13133 -20891
rect 13193 -20941 13203 -20881
rect 12803 -20951 13203 -20941
rect 13261 -20531 13661 -20521
rect 13261 -20591 13271 -20531
rect 13331 -20581 13591 -20531
rect 13331 -20591 13341 -20581
rect 13261 -20601 13341 -20591
rect 13581 -20591 13591 -20581
rect 13651 -20591 13661 -20531
rect 13581 -20601 13661 -20591
rect 13261 -20871 13321 -20601
rect 13591 -20611 13661 -20601
rect 13401 -20661 13431 -20641
rect 13381 -20701 13431 -20661
rect 13491 -20661 13521 -20641
rect 13491 -20701 13541 -20661
rect 13381 -20771 13541 -20701
rect 13381 -20811 13431 -20771
rect 13401 -20831 13431 -20811
rect 13491 -20811 13541 -20771
rect 13491 -20831 13521 -20811
rect 13601 -20871 13661 -20611
rect 13261 -20881 13341 -20871
rect 13261 -20941 13271 -20881
rect 13331 -20891 13341 -20881
rect 13581 -20881 13661 -20871
rect 13581 -20891 13591 -20881
rect 13331 -20941 13591 -20891
rect 13651 -20941 13661 -20881
rect 13261 -20951 13661 -20941
rect 13717 -20531 14117 -20521
rect 13717 -20591 13727 -20531
rect 13787 -20581 14047 -20531
rect 13787 -20591 13797 -20581
rect 13717 -20601 13797 -20591
rect 14037 -20591 14047 -20581
rect 14107 -20591 14117 -20531
rect 14037 -20601 14117 -20591
rect 13717 -20871 13777 -20601
rect 14047 -20611 14117 -20601
rect 13857 -20661 13887 -20641
rect 13837 -20701 13887 -20661
rect 13947 -20661 13977 -20641
rect 13947 -20701 13997 -20661
rect 13837 -20771 13997 -20701
rect 13837 -20811 13887 -20771
rect 13857 -20831 13887 -20811
rect 13947 -20811 13997 -20771
rect 13947 -20831 13977 -20811
rect 14057 -20871 14117 -20611
rect 13717 -20881 13797 -20871
rect 13717 -20941 13727 -20881
rect 13787 -20891 13797 -20881
rect 14037 -20881 14117 -20871
rect 14037 -20891 14047 -20881
rect 13787 -20941 14047 -20891
rect 14107 -20941 14117 -20881
rect 13717 -20951 14117 -20941
rect 14173 -20531 14573 -20521
rect 14173 -20591 14183 -20531
rect 14243 -20581 14503 -20531
rect 14243 -20591 14253 -20581
rect 14173 -20601 14253 -20591
rect 14493 -20591 14503 -20581
rect 14563 -20591 14573 -20531
rect 14493 -20601 14573 -20591
rect 14173 -20871 14233 -20601
rect 14503 -20611 14573 -20601
rect 14313 -20661 14343 -20641
rect 14293 -20701 14343 -20661
rect 14403 -20661 14433 -20641
rect 14403 -20701 14453 -20661
rect 14293 -20771 14453 -20701
rect 14293 -20811 14343 -20771
rect 14313 -20831 14343 -20811
rect 14403 -20811 14453 -20771
rect 14403 -20831 14433 -20811
rect 14513 -20871 14573 -20611
rect 14173 -20881 14253 -20871
rect 14173 -20941 14183 -20881
rect 14243 -20891 14253 -20881
rect 14493 -20881 14573 -20871
rect 14493 -20891 14503 -20881
rect 14243 -20941 14503 -20891
rect 14563 -20941 14573 -20881
rect 14173 -20951 14573 -20941
rect 14631 -20531 15031 -20521
rect 14631 -20591 14641 -20531
rect 14701 -20581 14961 -20531
rect 14701 -20591 14711 -20581
rect 14631 -20601 14711 -20591
rect 14951 -20591 14961 -20581
rect 15021 -20591 15031 -20531
rect 14951 -20601 15031 -20591
rect 14631 -20871 14691 -20601
rect 14961 -20611 15031 -20601
rect 14771 -20661 14801 -20641
rect 14751 -20701 14801 -20661
rect 14861 -20661 14891 -20641
rect 14861 -20701 14911 -20661
rect 14751 -20771 14911 -20701
rect 14751 -20811 14801 -20771
rect 14771 -20831 14801 -20811
rect 14861 -20811 14911 -20771
rect 14861 -20831 14891 -20811
rect 14971 -20871 15031 -20611
rect 14631 -20881 14711 -20871
rect 14631 -20941 14641 -20881
rect 14701 -20891 14711 -20881
rect 14951 -20881 15031 -20871
rect 14951 -20891 14961 -20881
rect 14701 -20941 14961 -20891
rect 15021 -20941 15031 -20881
rect 14631 -20951 15031 -20941
rect 15087 -20531 15487 -20521
rect 15087 -20591 15097 -20531
rect 15157 -20581 15417 -20531
rect 15157 -20591 15167 -20581
rect 15087 -20601 15167 -20591
rect 15407 -20591 15417 -20581
rect 15477 -20591 15487 -20531
rect 15407 -20601 15487 -20591
rect 15087 -20871 15147 -20601
rect 15417 -20611 15487 -20601
rect 15227 -20661 15257 -20641
rect 15207 -20701 15257 -20661
rect 15317 -20661 15347 -20641
rect 15317 -20701 15367 -20661
rect 15207 -20771 15367 -20701
rect 15207 -20811 15257 -20771
rect 15227 -20831 15257 -20811
rect 15317 -20811 15367 -20771
rect 15317 -20831 15347 -20811
rect 15427 -20871 15487 -20611
rect 15087 -20881 15167 -20871
rect 15087 -20941 15097 -20881
rect 15157 -20891 15167 -20881
rect 15407 -20881 15487 -20871
rect 15407 -20891 15417 -20881
rect 15157 -20941 15417 -20891
rect 15477 -20941 15487 -20881
rect 15087 -20951 15487 -20941
rect 1 -21047 401 -21037
rect 1 -21107 11 -21047
rect 71 -21097 331 -21047
rect 71 -21107 81 -21097
rect 1 -21117 81 -21107
rect 321 -21107 331 -21097
rect 391 -21107 401 -21047
rect 321 -21117 401 -21107
rect 1 -21387 61 -21117
rect 331 -21127 401 -21117
rect 141 -21177 171 -21157
rect 121 -21217 171 -21177
rect 231 -21177 261 -21157
rect 231 -21217 281 -21177
rect 121 -21287 281 -21217
rect 121 -21327 171 -21287
rect 141 -21347 171 -21327
rect 231 -21327 281 -21287
rect 231 -21347 261 -21327
rect 341 -21387 401 -21127
rect 1 -21397 81 -21387
rect 1 -21457 11 -21397
rect 71 -21407 81 -21397
rect 321 -21397 401 -21387
rect 321 -21407 331 -21397
rect 71 -21457 331 -21407
rect 391 -21457 401 -21397
rect 1 -21467 401 -21457
rect 457 -21047 857 -21037
rect 457 -21107 467 -21047
rect 527 -21097 787 -21047
rect 527 -21107 537 -21097
rect 457 -21117 537 -21107
rect 777 -21107 787 -21097
rect 847 -21107 857 -21047
rect 777 -21117 857 -21107
rect 457 -21387 517 -21117
rect 787 -21127 857 -21117
rect 597 -21177 627 -21157
rect 577 -21217 627 -21177
rect 687 -21177 717 -21157
rect 687 -21217 737 -21177
rect 577 -21287 737 -21217
rect 577 -21327 627 -21287
rect 597 -21347 627 -21327
rect 687 -21327 737 -21287
rect 687 -21347 717 -21327
rect 797 -21387 857 -21127
rect 457 -21397 537 -21387
rect 457 -21457 467 -21397
rect 527 -21407 537 -21397
rect 777 -21397 857 -21387
rect 777 -21407 787 -21397
rect 527 -21457 787 -21407
rect 847 -21457 857 -21397
rect 457 -21467 857 -21457
rect 913 -21047 1313 -21037
rect 913 -21107 923 -21047
rect 983 -21097 1243 -21047
rect 983 -21107 993 -21097
rect 913 -21117 993 -21107
rect 1233 -21107 1243 -21097
rect 1303 -21107 1313 -21047
rect 1233 -21117 1313 -21107
rect 913 -21387 973 -21117
rect 1243 -21127 1313 -21117
rect 1053 -21177 1083 -21157
rect 1033 -21217 1083 -21177
rect 1143 -21177 1173 -21157
rect 1143 -21217 1193 -21177
rect 1033 -21287 1193 -21217
rect 1033 -21327 1083 -21287
rect 1053 -21347 1083 -21327
rect 1143 -21327 1193 -21287
rect 1143 -21347 1173 -21327
rect 1253 -21387 1313 -21127
rect 913 -21397 993 -21387
rect 913 -21457 923 -21397
rect 983 -21407 993 -21397
rect 1233 -21397 1313 -21387
rect 1233 -21407 1243 -21397
rect 983 -21457 1243 -21407
rect 1303 -21457 1313 -21397
rect 913 -21467 1313 -21457
rect 1371 -21047 1771 -21037
rect 1371 -21107 1381 -21047
rect 1441 -21097 1701 -21047
rect 1441 -21107 1451 -21097
rect 1371 -21117 1451 -21107
rect 1691 -21107 1701 -21097
rect 1761 -21107 1771 -21047
rect 1691 -21117 1771 -21107
rect 1371 -21387 1431 -21117
rect 1701 -21127 1771 -21117
rect 1511 -21177 1541 -21157
rect 1491 -21217 1541 -21177
rect 1601 -21177 1631 -21157
rect 1601 -21217 1651 -21177
rect 1491 -21287 1651 -21217
rect 1491 -21327 1541 -21287
rect 1511 -21347 1541 -21327
rect 1601 -21327 1651 -21287
rect 1601 -21347 1631 -21327
rect 1711 -21387 1771 -21127
rect 1371 -21397 1451 -21387
rect 1371 -21457 1381 -21397
rect 1441 -21407 1451 -21397
rect 1691 -21397 1771 -21387
rect 1691 -21407 1701 -21397
rect 1441 -21457 1701 -21407
rect 1761 -21457 1771 -21397
rect 1371 -21467 1771 -21457
rect 1827 -21047 2227 -21037
rect 1827 -21107 1837 -21047
rect 1897 -21097 2157 -21047
rect 1897 -21107 1907 -21097
rect 1827 -21117 1907 -21107
rect 2147 -21107 2157 -21097
rect 2217 -21107 2227 -21047
rect 2147 -21117 2227 -21107
rect 1827 -21387 1887 -21117
rect 2157 -21127 2227 -21117
rect 1967 -21177 1997 -21157
rect 1947 -21217 1997 -21177
rect 2057 -21177 2087 -21157
rect 2057 -21217 2107 -21177
rect 1947 -21287 2107 -21217
rect 1947 -21327 1997 -21287
rect 1967 -21347 1997 -21327
rect 2057 -21327 2107 -21287
rect 2057 -21347 2087 -21327
rect 2167 -21387 2227 -21127
rect 1827 -21397 1907 -21387
rect 1827 -21457 1837 -21397
rect 1897 -21407 1907 -21397
rect 2147 -21397 2227 -21387
rect 2147 -21407 2157 -21397
rect 1897 -21457 2157 -21407
rect 2217 -21457 2227 -21397
rect 1827 -21467 2227 -21457
rect 2283 -21047 2683 -21037
rect 2283 -21107 2293 -21047
rect 2353 -21097 2613 -21047
rect 2353 -21107 2363 -21097
rect 2283 -21117 2363 -21107
rect 2603 -21107 2613 -21097
rect 2673 -21107 2683 -21047
rect 2603 -21117 2683 -21107
rect 2283 -21387 2343 -21117
rect 2613 -21127 2683 -21117
rect 2423 -21177 2453 -21157
rect 2403 -21217 2453 -21177
rect 2513 -21177 2543 -21157
rect 2513 -21217 2563 -21177
rect 2403 -21287 2563 -21217
rect 2403 -21327 2453 -21287
rect 2423 -21347 2453 -21327
rect 2513 -21327 2563 -21287
rect 2513 -21347 2543 -21327
rect 2623 -21387 2683 -21127
rect 2283 -21397 2363 -21387
rect 2283 -21457 2293 -21397
rect 2353 -21407 2363 -21397
rect 2603 -21397 2683 -21387
rect 2603 -21407 2613 -21397
rect 2353 -21457 2613 -21407
rect 2673 -21457 2683 -21397
rect 2283 -21467 2683 -21457
rect 2741 -21047 3141 -21037
rect 2741 -21107 2751 -21047
rect 2811 -21097 3071 -21047
rect 2811 -21107 2821 -21097
rect 2741 -21117 2821 -21107
rect 3061 -21107 3071 -21097
rect 3131 -21107 3141 -21047
rect 3061 -21117 3141 -21107
rect 2741 -21387 2801 -21117
rect 3071 -21127 3141 -21117
rect 2881 -21177 2911 -21157
rect 2861 -21217 2911 -21177
rect 2971 -21177 3001 -21157
rect 2971 -21217 3021 -21177
rect 2861 -21287 3021 -21217
rect 2861 -21327 2911 -21287
rect 2881 -21347 2911 -21327
rect 2971 -21327 3021 -21287
rect 2971 -21347 3001 -21327
rect 3081 -21387 3141 -21127
rect 2741 -21397 2821 -21387
rect 2741 -21457 2751 -21397
rect 2811 -21407 2821 -21397
rect 3061 -21397 3141 -21387
rect 3061 -21407 3071 -21397
rect 2811 -21457 3071 -21407
rect 3131 -21457 3141 -21397
rect 2741 -21467 3141 -21457
rect 3197 -21047 3597 -21037
rect 3197 -21107 3207 -21047
rect 3267 -21097 3527 -21047
rect 3267 -21107 3277 -21097
rect 3197 -21117 3277 -21107
rect 3517 -21107 3527 -21097
rect 3587 -21107 3597 -21047
rect 3517 -21117 3597 -21107
rect 3197 -21387 3257 -21117
rect 3527 -21127 3597 -21117
rect 3337 -21177 3367 -21157
rect 3317 -21217 3367 -21177
rect 3427 -21177 3457 -21157
rect 3427 -21217 3477 -21177
rect 3317 -21287 3477 -21217
rect 3317 -21327 3367 -21287
rect 3337 -21347 3367 -21327
rect 3427 -21327 3477 -21287
rect 3427 -21347 3457 -21327
rect 3537 -21387 3597 -21127
rect 3197 -21397 3277 -21387
rect 3197 -21457 3207 -21397
rect 3267 -21407 3277 -21397
rect 3517 -21397 3597 -21387
rect 3517 -21407 3527 -21397
rect 3267 -21457 3527 -21407
rect 3587 -21457 3597 -21397
rect 3197 -21467 3597 -21457
rect 3653 -21047 4053 -21037
rect 3653 -21107 3663 -21047
rect 3723 -21097 3983 -21047
rect 3723 -21107 3733 -21097
rect 3653 -21117 3733 -21107
rect 3973 -21107 3983 -21097
rect 4043 -21107 4053 -21047
rect 3973 -21117 4053 -21107
rect 3653 -21387 3713 -21117
rect 3983 -21127 4053 -21117
rect 3793 -21177 3823 -21157
rect 3773 -21217 3823 -21177
rect 3883 -21177 3913 -21157
rect 3883 -21217 3933 -21177
rect 3773 -21287 3933 -21217
rect 3773 -21327 3823 -21287
rect 3793 -21347 3823 -21327
rect 3883 -21327 3933 -21287
rect 3883 -21347 3913 -21327
rect 3993 -21387 4053 -21127
rect 3653 -21397 3733 -21387
rect 3653 -21457 3663 -21397
rect 3723 -21407 3733 -21397
rect 3973 -21397 4053 -21387
rect 3973 -21407 3983 -21397
rect 3723 -21457 3983 -21407
rect 4043 -21457 4053 -21397
rect 3653 -21467 4053 -21457
rect 4111 -21047 4511 -21037
rect 4111 -21107 4121 -21047
rect 4181 -21097 4441 -21047
rect 4181 -21107 4191 -21097
rect 4111 -21117 4191 -21107
rect 4431 -21107 4441 -21097
rect 4501 -21107 4511 -21047
rect 4431 -21117 4511 -21107
rect 4111 -21387 4171 -21117
rect 4441 -21127 4511 -21117
rect 4251 -21177 4281 -21157
rect 4231 -21217 4281 -21177
rect 4341 -21177 4371 -21157
rect 4341 -21217 4391 -21177
rect 4231 -21287 4391 -21217
rect 4231 -21327 4281 -21287
rect 4251 -21347 4281 -21327
rect 4341 -21327 4391 -21287
rect 4341 -21347 4371 -21327
rect 4451 -21387 4511 -21127
rect 4111 -21397 4191 -21387
rect 4111 -21457 4121 -21397
rect 4181 -21407 4191 -21397
rect 4431 -21397 4511 -21387
rect 4431 -21407 4441 -21397
rect 4181 -21457 4441 -21407
rect 4501 -21457 4511 -21397
rect 4111 -21467 4511 -21457
rect 4567 -21047 4967 -21037
rect 4567 -21107 4577 -21047
rect 4637 -21097 4897 -21047
rect 4637 -21107 4647 -21097
rect 4567 -21117 4647 -21107
rect 4887 -21107 4897 -21097
rect 4957 -21107 4967 -21047
rect 4887 -21117 4967 -21107
rect 4567 -21387 4627 -21117
rect 4897 -21127 4967 -21117
rect 4707 -21177 4737 -21157
rect 4687 -21217 4737 -21177
rect 4797 -21177 4827 -21157
rect 4797 -21217 4847 -21177
rect 4687 -21287 4847 -21217
rect 4687 -21327 4737 -21287
rect 4707 -21347 4737 -21327
rect 4797 -21327 4847 -21287
rect 4797 -21347 4827 -21327
rect 4907 -21387 4967 -21127
rect 4567 -21397 4647 -21387
rect 4567 -21457 4577 -21397
rect 4637 -21407 4647 -21397
rect 4887 -21397 4967 -21387
rect 4887 -21407 4897 -21397
rect 4637 -21457 4897 -21407
rect 4957 -21457 4967 -21397
rect 4567 -21467 4967 -21457
rect 5023 -21047 5423 -21037
rect 5023 -21107 5033 -21047
rect 5093 -21097 5353 -21047
rect 5093 -21107 5103 -21097
rect 5023 -21117 5103 -21107
rect 5343 -21107 5353 -21097
rect 5413 -21107 5423 -21047
rect 5343 -21117 5423 -21107
rect 5023 -21387 5083 -21117
rect 5353 -21127 5423 -21117
rect 5163 -21177 5193 -21157
rect 5143 -21217 5193 -21177
rect 5253 -21177 5283 -21157
rect 5253 -21217 5303 -21177
rect 5143 -21287 5303 -21217
rect 5143 -21327 5193 -21287
rect 5163 -21347 5193 -21327
rect 5253 -21327 5303 -21287
rect 5253 -21347 5283 -21327
rect 5363 -21387 5423 -21127
rect 5023 -21397 5103 -21387
rect 5023 -21457 5033 -21397
rect 5093 -21407 5103 -21397
rect 5343 -21397 5423 -21387
rect 5343 -21407 5353 -21397
rect 5093 -21457 5353 -21407
rect 5413 -21457 5423 -21397
rect 5023 -21467 5423 -21457
rect 5481 -21047 5881 -21037
rect 5481 -21107 5491 -21047
rect 5551 -21097 5811 -21047
rect 5551 -21107 5561 -21097
rect 5481 -21117 5561 -21107
rect 5801 -21107 5811 -21097
rect 5871 -21107 5881 -21047
rect 5801 -21117 5881 -21107
rect 5481 -21387 5541 -21117
rect 5811 -21127 5881 -21117
rect 5621 -21177 5651 -21157
rect 5601 -21217 5651 -21177
rect 5711 -21177 5741 -21157
rect 5711 -21217 5761 -21177
rect 5601 -21287 5761 -21217
rect 5601 -21327 5651 -21287
rect 5621 -21347 5651 -21327
rect 5711 -21327 5761 -21287
rect 5711 -21347 5741 -21327
rect 5821 -21387 5881 -21127
rect 5481 -21397 5561 -21387
rect 5481 -21457 5491 -21397
rect 5551 -21407 5561 -21397
rect 5801 -21397 5881 -21387
rect 5801 -21407 5811 -21397
rect 5551 -21457 5811 -21407
rect 5871 -21457 5881 -21397
rect 5481 -21467 5881 -21457
rect 5937 -21047 6337 -21037
rect 5937 -21107 5947 -21047
rect 6007 -21097 6267 -21047
rect 6007 -21107 6017 -21097
rect 5937 -21117 6017 -21107
rect 6257 -21107 6267 -21097
rect 6327 -21107 6337 -21047
rect 6257 -21117 6337 -21107
rect 5937 -21387 5997 -21117
rect 6267 -21127 6337 -21117
rect 6077 -21177 6107 -21157
rect 6057 -21217 6107 -21177
rect 6167 -21177 6197 -21157
rect 6167 -21217 6217 -21177
rect 6057 -21287 6217 -21217
rect 6057 -21327 6107 -21287
rect 6077 -21347 6107 -21327
rect 6167 -21327 6217 -21287
rect 6167 -21347 6197 -21327
rect 6277 -21387 6337 -21127
rect 5937 -21397 6017 -21387
rect 5937 -21457 5947 -21397
rect 6007 -21407 6017 -21397
rect 6257 -21397 6337 -21387
rect 6257 -21407 6267 -21397
rect 6007 -21457 6267 -21407
rect 6327 -21457 6337 -21397
rect 5937 -21467 6337 -21457
rect 6393 -21047 6793 -21037
rect 6393 -21107 6403 -21047
rect 6463 -21097 6723 -21047
rect 6463 -21107 6473 -21097
rect 6393 -21117 6473 -21107
rect 6713 -21107 6723 -21097
rect 6783 -21107 6793 -21047
rect 6713 -21117 6793 -21107
rect 6393 -21387 6453 -21117
rect 6723 -21127 6793 -21117
rect 6533 -21177 6563 -21157
rect 6513 -21217 6563 -21177
rect 6623 -21177 6653 -21157
rect 6623 -21217 6673 -21177
rect 6513 -21287 6673 -21217
rect 6513 -21327 6563 -21287
rect 6533 -21347 6563 -21327
rect 6623 -21327 6673 -21287
rect 6623 -21347 6653 -21327
rect 6733 -21387 6793 -21127
rect 6393 -21397 6473 -21387
rect 6393 -21457 6403 -21397
rect 6463 -21407 6473 -21397
rect 6713 -21397 6793 -21387
rect 6713 -21407 6723 -21397
rect 6463 -21457 6723 -21407
rect 6783 -21457 6793 -21397
rect 6393 -21467 6793 -21457
rect 6851 -21047 7251 -21037
rect 6851 -21107 6861 -21047
rect 6921 -21097 7181 -21047
rect 6921 -21107 6931 -21097
rect 6851 -21117 6931 -21107
rect 7171 -21107 7181 -21097
rect 7241 -21107 7251 -21047
rect 7171 -21117 7251 -21107
rect 6851 -21387 6911 -21117
rect 7181 -21127 7251 -21117
rect 6991 -21177 7021 -21157
rect 6971 -21217 7021 -21177
rect 7081 -21177 7111 -21157
rect 7081 -21217 7131 -21177
rect 6971 -21287 7131 -21217
rect 6971 -21327 7021 -21287
rect 6991 -21347 7021 -21327
rect 7081 -21327 7131 -21287
rect 7081 -21347 7111 -21327
rect 7191 -21387 7251 -21127
rect 6851 -21397 6931 -21387
rect 6851 -21457 6861 -21397
rect 6921 -21407 6931 -21397
rect 7171 -21397 7251 -21387
rect 7171 -21407 7181 -21397
rect 6921 -21457 7181 -21407
rect 7241 -21457 7251 -21397
rect 6851 -21467 7251 -21457
rect 7307 -21047 7707 -21037
rect 7307 -21107 7317 -21047
rect 7377 -21097 7637 -21047
rect 7377 -21107 7387 -21097
rect 7307 -21117 7387 -21107
rect 7627 -21107 7637 -21097
rect 7697 -21107 7707 -21047
rect 7627 -21117 7707 -21107
rect 7307 -21387 7367 -21117
rect 7637 -21127 7707 -21117
rect 7447 -21177 7477 -21157
rect 7427 -21217 7477 -21177
rect 7537 -21177 7567 -21157
rect 7537 -21217 7587 -21177
rect 7427 -21287 7587 -21217
rect 7427 -21327 7477 -21287
rect 7447 -21347 7477 -21327
rect 7537 -21327 7587 -21287
rect 7537 -21347 7567 -21327
rect 7647 -21387 7707 -21127
rect 7307 -21397 7387 -21387
rect 7307 -21457 7317 -21397
rect 7377 -21407 7387 -21397
rect 7627 -21397 7707 -21387
rect 7627 -21407 7637 -21397
rect 7377 -21457 7637 -21407
rect 7697 -21457 7707 -21397
rect 7307 -21467 7707 -21457
rect 7763 -21047 8163 -21037
rect 7763 -21107 7773 -21047
rect 7833 -21097 8093 -21047
rect 7833 -21107 7843 -21097
rect 7763 -21117 7843 -21107
rect 8083 -21107 8093 -21097
rect 8153 -21107 8163 -21047
rect 8083 -21117 8163 -21107
rect 7763 -21387 7823 -21117
rect 8093 -21127 8163 -21117
rect 7903 -21177 7933 -21157
rect 7883 -21217 7933 -21177
rect 7993 -21177 8023 -21157
rect 7993 -21217 8043 -21177
rect 7883 -21287 8043 -21217
rect 7883 -21327 7933 -21287
rect 7903 -21347 7933 -21327
rect 7993 -21327 8043 -21287
rect 7993 -21347 8023 -21327
rect 8103 -21387 8163 -21127
rect 7763 -21397 7843 -21387
rect 7763 -21457 7773 -21397
rect 7833 -21407 7843 -21397
rect 8083 -21397 8163 -21387
rect 8083 -21407 8093 -21397
rect 7833 -21457 8093 -21407
rect 8153 -21457 8163 -21397
rect 7763 -21467 8163 -21457
rect 8237 -21047 8637 -21037
rect 8237 -21107 8247 -21047
rect 8307 -21097 8567 -21047
rect 8307 -21107 8317 -21097
rect 8237 -21117 8317 -21107
rect 8557 -21107 8567 -21097
rect 8627 -21107 8637 -21047
rect 8557 -21117 8637 -21107
rect 8237 -21387 8297 -21117
rect 8567 -21127 8637 -21117
rect 8377 -21177 8407 -21157
rect 8357 -21217 8407 -21177
rect 8467 -21177 8497 -21157
rect 8467 -21217 8517 -21177
rect 8357 -21287 8517 -21217
rect 8357 -21327 8407 -21287
rect 8377 -21347 8407 -21327
rect 8467 -21327 8517 -21287
rect 8467 -21347 8497 -21327
rect 8577 -21387 8637 -21127
rect 8237 -21397 8317 -21387
rect 8237 -21457 8247 -21397
rect 8307 -21407 8317 -21397
rect 8557 -21397 8637 -21387
rect 8557 -21407 8567 -21397
rect 8307 -21457 8567 -21407
rect 8627 -21457 8637 -21397
rect 8237 -21467 8637 -21457
rect 8693 -21047 9093 -21037
rect 8693 -21107 8703 -21047
rect 8763 -21097 9023 -21047
rect 8763 -21107 8773 -21097
rect 8693 -21117 8773 -21107
rect 9013 -21107 9023 -21097
rect 9083 -21107 9093 -21047
rect 9013 -21117 9093 -21107
rect 8693 -21387 8753 -21117
rect 9023 -21127 9093 -21117
rect 8833 -21177 8863 -21157
rect 8813 -21217 8863 -21177
rect 8923 -21177 8953 -21157
rect 8923 -21217 8973 -21177
rect 8813 -21287 8973 -21217
rect 8813 -21327 8863 -21287
rect 8833 -21347 8863 -21327
rect 8923 -21327 8973 -21287
rect 8923 -21347 8953 -21327
rect 9033 -21387 9093 -21127
rect 8693 -21397 8773 -21387
rect 8693 -21457 8703 -21397
rect 8763 -21407 8773 -21397
rect 9013 -21397 9093 -21387
rect 9013 -21407 9023 -21397
rect 8763 -21457 9023 -21407
rect 9083 -21457 9093 -21397
rect 8693 -21467 9093 -21457
rect 9151 -21047 9551 -21037
rect 9151 -21107 9161 -21047
rect 9221 -21097 9481 -21047
rect 9221 -21107 9231 -21097
rect 9151 -21117 9231 -21107
rect 9471 -21107 9481 -21097
rect 9541 -21107 9551 -21047
rect 9471 -21117 9551 -21107
rect 9151 -21387 9211 -21117
rect 9481 -21127 9551 -21117
rect 9291 -21177 9321 -21157
rect 9271 -21217 9321 -21177
rect 9381 -21177 9411 -21157
rect 9381 -21217 9431 -21177
rect 9271 -21287 9431 -21217
rect 9271 -21327 9321 -21287
rect 9291 -21347 9321 -21327
rect 9381 -21327 9431 -21287
rect 9381 -21347 9411 -21327
rect 9491 -21387 9551 -21127
rect 9151 -21397 9231 -21387
rect 9151 -21457 9161 -21397
rect 9221 -21407 9231 -21397
rect 9471 -21397 9551 -21387
rect 9471 -21407 9481 -21397
rect 9221 -21457 9481 -21407
rect 9541 -21457 9551 -21397
rect 9151 -21467 9551 -21457
rect 9607 -21047 10007 -21037
rect 9607 -21107 9617 -21047
rect 9677 -21097 9937 -21047
rect 9677 -21107 9687 -21097
rect 9607 -21117 9687 -21107
rect 9927 -21107 9937 -21097
rect 9997 -21107 10007 -21047
rect 9927 -21117 10007 -21107
rect 9607 -21387 9667 -21117
rect 9937 -21127 10007 -21117
rect 9747 -21177 9777 -21157
rect 9727 -21217 9777 -21177
rect 9837 -21177 9867 -21157
rect 9837 -21217 9887 -21177
rect 9727 -21287 9887 -21217
rect 9727 -21327 9777 -21287
rect 9747 -21347 9777 -21327
rect 9837 -21327 9887 -21287
rect 9837 -21347 9867 -21327
rect 9947 -21387 10007 -21127
rect 9607 -21397 9687 -21387
rect 9607 -21457 9617 -21397
rect 9677 -21407 9687 -21397
rect 9927 -21397 10007 -21387
rect 9927 -21407 9937 -21397
rect 9677 -21457 9937 -21407
rect 9997 -21457 10007 -21397
rect 9607 -21467 10007 -21457
rect 10063 -21047 10463 -21037
rect 10063 -21107 10073 -21047
rect 10133 -21097 10393 -21047
rect 10133 -21107 10143 -21097
rect 10063 -21117 10143 -21107
rect 10383 -21107 10393 -21097
rect 10453 -21107 10463 -21047
rect 10383 -21117 10463 -21107
rect 10063 -21387 10123 -21117
rect 10393 -21127 10463 -21117
rect 10203 -21177 10233 -21157
rect 10183 -21217 10233 -21177
rect 10293 -21177 10323 -21157
rect 10293 -21217 10343 -21177
rect 10183 -21287 10343 -21217
rect 10183 -21327 10233 -21287
rect 10203 -21347 10233 -21327
rect 10293 -21327 10343 -21287
rect 10293 -21347 10323 -21327
rect 10403 -21387 10463 -21127
rect 10063 -21397 10143 -21387
rect 10063 -21457 10073 -21397
rect 10133 -21407 10143 -21397
rect 10383 -21397 10463 -21387
rect 10383 -21407 10393 -21397
rect 10133 -21457 10393 -21407
rect 10453 -21457 10463 -21397
rect 10063 -21467 10463 -21457
rect 10521 -21047 10921 -21037
rect 10521 -21107 10531 -21047
rect 10591 -21097 10851 -21047
rect 10591 -21107 10601 -21097
rect 10521 -21117 10601 -21107
rect 10841 -21107 10851 -21097
rect 10911 -21107 10921 -21047
rect 10841 -21117 10921 -21107
rect 10521 -21387 10581 -21117
rect 10851 -21127 10921 -21117
rect 10661 -21177 10691 -21157
rect 10641 -21217 10691 -21177
rect 10751 -21177 10781 -21157
rect 10751 -21217 10801 -21177
rect 10641 -21287 10801 -21217
rect 10641 -21327 10691 -21287
rect 10661 -21347 10691 -21327
rect 10751 -21327 10801 -21287
rect 10751 -21347 10781 -21327
rect 10861 -21387 10921 -21127
rect 10521 -21397 10601 -21387
rect 10521 -21457 10531 -21397
rect 10591 -21407 10601 -21397
rect 10841 -21397 10921 -21387
rect 10841 -21407 10851 -21397
rect 10591 -21457 10851 -21407
rect 10911 -21457 10921 -21397
rect 10521 -21467 10921 -21457
rect 10977 -21047 11377 -21037
rect 10977 -21107 10987 -21047
rect 11047 -21097 11307 -21047
rect 11047 -21107 11057 -21097
rect 10977 -21117 11057 -21107
rect 11297 -21107 11307 -21097
rect 11367 -21107 11377 -21047
rect 11297 -21117 11377 -21107
rect 10977 -21387 11037 -21117
rect 11307 -21127 11377 -21117
rect 11117 -21177 11147 -21157
rect 11097 -21217 11147 -21177
rect 11207 -21177 11237 -21157
rect 11207 -21217 11257 -21177
rect 11097 -21287 11257 -21217
rect 11097 -21327 11147 -21287
rect 11117 -21347 11147 -21327
rect 11207 -21327 11257 -21287
rect 11207 -21347 11237 -21327
rect 11317 -21387 11377 -21127
rect 10977 -21397 11057 -21387
rect 10977 -21457 10987 -21397
rect 11047 -21407 11057 -21397
rect 11297 -21397 11377 -21387
rect 11297 -21407 11307 -21397
rect 11047 -21457 11307 -21407
rect 11367 -21457 11377 -21397
rect 10977 -21467 11377 -21457
rect 11433 -21047 11833 -21037
rect 11433 -21107 11443 -21047
rect 11503 -21097 11763 -21047
rect 11503 -21107 11513 -21097
rect 11433 -21117 11513 -21107
rect 11753 -21107 11763 -21097
rect 11823 -21107 11833 -21047
rect 11753 -21117 11833 -21107
rect 11433 -21387 11493 -21117
rect 11763 -21127 11833 -21117
rect 11573 -21177 11603 -21157
rect 11553 -21217 11603 -21177
rect 11663 -21177 11693 -21157
rect 11663 -21217 11713 -21177
rect 11553 -21287 11713 -21217
rect 11553 -21327 11603 -21287
rect 11573 -21347 11603 -21327
rect 11663 -21327 11713 -21287
rect 11663 -21347 11693 -21327
rect 11773 -21387 11833 -21127
rect 11433 -21397 11513 -21387
rect 11433 -21457 11443 -21397
rect 11503 -21407 11513 -21397
rect 11753 -21397 11833 -21387
rect 11753 -21407 11763 -21397
rect 11503 -21457 11763 -21407
rect 11823 -21457 11833 -21397
rect 11433 -21467 11833 -21457
rect 11891 -21047 12291 -21037
rect 11891 -21107 11901 -21047
rect 11961 -21097 12221 -21047
rect 11961 -21107 11971 -21097
rect 11891 -21117 11971 -21107
rect 12211 -21107 12221 -21097
rect 12281 -21107 12291 -21047
rect 12211 -21117 12291 -21107
rect 11891 -21387 11951 -21117
rect 12221 -21127 12291 -21117
rect 12031 -21177 12061 -21157
rect 12011 -21217 12061 -21177
rect 12121 -21177 12151 -21157
rect 12121 -21217 12171 -21177
rect 12011 -21287 12171 -21217
rect 12011 -21327 12061 -21287
rect 12031 -21347 12061 -21327
rect 12121 -21327 12171 -21287
rect 12121 -21347 12151 -21327
rect 12231 -21387 12291 -21127
rect 11891 -21397 11971 -21387
rect 11891 -21457 11901 -21397
rect 11961 -21407 11971 -21397
rect 12211 -21397 12291 -21387
rect 12211 -21407 12221 -21397
rect 11961 -21457 12221 -21407
rect 12281 -21457 12291 -21397
rect 11891 -21467 12291 -21457
rect 12347 -21047 12747 -21037
rect 12347 -21107 12357 -21047
rect 12417 -21097 12677 -21047
rect 12417 -21107 12427 -21097
rect 12347 -21117 12427 -21107
rect 12667 -21107 12677 -21097
rect 12737 -21107 12747 -21047
rect 12667 -21117 12747 -21107
rect 12347 -21387 12407 -21117
rect 12677 -21127 12747 -21117
rect 12487 -21177 12517 -21157
rect 12467 -21217 12517 -21177
rect 12577 -21177 12607 -21157
rect 12577 -21217 12627 -21177
rect 12467 -21287 12627 -21217
rect 12467 -21327 12517 -21287
rect 12487 -21347 12517 -21327
rect 12577 -21327 12627 -21287
rect 12577 -21347 12607 -21327
rect 12687 -21387 12747 -21127
rect 12347 -21397 12427 -21387
rect 12347 -21457 12357 -21397
rect 12417 -21407 12427 -21397
rect 12667 -21397 12747 -21387
rect 12667 -21407 12677 -21397
rect 12417 -21457 12677 -21407
rect 12737 -21457 12747 -21397
rect 12347 -21467 12747 -21457
rect 12803 -21047 13203 -21037
rect 12803 -21107 12813 -21047
rect 12873 -21097 13133 -21047
rect 12873 -21107 12883 -21097
rect 12803 -21117 12883 -21107
rect 13123 -21107 13133 -21097
rect 13193 -21107 13203 -21047
rect 13123 -21117 13203 -21107
rect 12803 -21387 12863 -21117
rect 13133 -21127 13203 -21117
rect 12943 -21177 12973 -21157
rect 12923 -21217 12973 -21177
rect 13033 -21177 13063 -21157
rect 13033 -21217 13083 -21177
rect 12923 -21287 13083 -21217
rect 12923 -21327 12973 -21287
rect 12943 -21347 12973 -21327
rect 13033 -21327 13083 -21287
rect 13033 -21347 13063 -21327
rect 13143 -21387 13203 -21127
rect 12803 -21397 12883 -21387
rect 12803 -21457 12813 -21397
rect 12873 -21407 12883 -21397
rect 13123 -21397 13203 -21387
rect 13123 -21407 13133 -21397
rect 12873 -21457 13133 -21407
rect 13193 -21457 13203 -21397
rect 12803 -21467 13203 -21457
rect 13261 -21047 13661 -21037
rect 13261 -21107 13271 -21047
rect 13331 -21097 13591 -21047
rect 13331 -21107 13341 -21097
rect 13261 -21117 13341 -21107
rect 13581 -21107 13591 -21097
rect 13651 -21107 13661 -21047
rect 13581 -21117 13661 -21107
rect 13261 -21387 13321 -21117
rect 13591 -21127 13661 -21117
rect 13401 -21177 13431 -21157
rect 13381 -21217 13431 -21177
rect 13491 -21177 13521 -21157
rect 13491 -21217 13541 -21177
rect 13381 -21287 13541 -21217
rect 13381 -21327 13431 -21287
rect 13401 -21347 13431 -21327
rect 13491 -21327 13541 -21287
rect 13491 -21347 13521 -21327
rect 13601 -21387 13661 -21127
rect 13261 -21397 13341 -21387
rect 13261 -21457 13271 -21397
rect 13331 -21407 13341 -21397
rect 13581 -21397 13661 -21387
rect 13581 -21407 13591 -21397
rect 13331 -21457 13591 -21407
rect 13651 -21457 13661 -21397
rect 13261 -21467 13661 -21457
rect 13717 -21047 14117 -21037
rect 13717 -21107 13727 -21047
rect 13787 -21097 14047 -21047
rect 13787 -21107 13797 -21097
rect 13717 -21117 13797 -21107
rect 14037 -21107 14047 -21097
rect 14107 -21107 14117 -21047
rect 14037 -21117 14117 -21107
rect 13717 -21387 13777 -21117
rect 14047 -21127 14117 -21117
rect 13857 -21177 13887 -21157
rect 13837 -21217 13887 -21177
rect 13947 -21177 13977 -21157
rect 13947 -21217 13997 -21177
rect 13837 -21287 13997 -21217
rect 13837 -21327 13887 -21287
rect 13857 -21347 13887 -21327
rect 13947 -21327 13997 -21287
rect 13947 -21347 13977 -21327
rect 14057 -21387 14117 -21127
rect 13717 -21397 13797 -21387
rect 13717 -21457 13727 -21397
rect 13787 -21407 13797 -21397
rect 14037 -21397 14117 -21387
rect 14037 -21407 14047 -21397
rect 13787 -21457 14047 -21407
rect 14107 -21457 14117 -21397
rect 13717 -21467 14117 -21457
rect 14173 -21047 14573 -21037
rect 14173 -21107 14183 -21047
rect 14243 -21097 14503 -21047
rect 14243 -21107 14253 -21097
rect 14173 -21117 14253 -21107
rect 14493 -21107 14503 -21097
rect 14563 -21107 14573 -21047
rect 14493 -21117 14573 -21107
rect 14173 -21387 14233 -21117
rect 14503 -21127 14573 -21117
rect 14313 -21177 14343 -21157
rect 14293 -21217 14343 -21177
rect 14403 -21177 14433 -21157
rect 14403 -21217 14453 -21177
rect 14293 -21287 14453 -21217
rect 14293 -21327 14343 -21287
rect 14313 -21347 14343 -21327
rect 14403 -21327 14453 -21287
rect 14403 -21347 14433 -21327
rect 14513 -21387 14573 -21127
rect 14173 -21397 14253 -21387
rect 14173 -21457 14183 -21397
rect 14243 -21407 14253 -21397
rect 14493 -21397 14573 -21387
rect 14493 -21407 14503 -21397
rect 14243 -21457 14503 -21407
rect 14563 -21457 14573 -21397
rect 14173 -21467 14573 -21457
rect 14631 -21047 15031 -21037
rect 14631 -21107 14641 -21047
rect 14701 -21097 14961 -21047
rect 14701 -21107 14711 -21097
rect 14631 -21117 14711 -21107
rect 14951 -21107 14961 -21097
rect 15021 -21107 15031 -21047
rect 14951 -21117 15031 -21107
rect 14631 -21387 14691 -21117
rect 14961 -21127 15031 -21117
rect 14771 -21177 14801 -21157
rect 14751 -21217 14801 -21177
rect 14861 -21177 14891 -21157
rect 14861 -21217 14911 -21177
rect 14751 -21287 14911 -21217
rect 14751 -21327 14801 -21287
rect 14771 -21347 14801 -21327
rect 14861 -21327 14911 -21287
rect 14861 -21347 14891 -21327
rect 14971 -21387 15031 -21127
rect 14631 -21397 14711 -21387
rect 14631 -21457 14641 -21397
rect 14701 -21407 14711 -21397
rect 14951 -21397 15031 -21387
rect 14951 -21407 14961 -21397
rect 14701 -21457 14961 -21407
rect 15021 -21457 15031 -21397
rect 14631 -21467 15031 -21457
rect 15087 -21047 15487 -21037
rect 15087 -21107 15097 -21047
rect 15157 -21097 15417 -21047
rect 15157 -21107 15167 -21097
rect 15087 -21117 15167 -21107
rect 15407 -21107 15417 -21097
rect 15477 -21107 15487 -21047
rect 15407 -21117 15487 -21107
rect 15087 -21387 15147 -21117
rect 15417 -21127 15487 -21117
rect 15227 -21177 15257 -21157
rect 15207 -21217 15257 -21177
rect 15317 -21177 15347 -21157
rect 15317 -21217 15367 -21177
rect 15207 -21287 15367 -21217
rect 15207 -21327 15257 -21287
rect 15227 -21347 15257 -21327
rect 15317 -21327 15367 -21287
rect 15317 -21347 15347 -21327
rect 15427 -21387 15487 -21127
rect 15087 -21397 15167 -21387
rect 15087 -21457 15097 -21397
rect 15157 -21407 15167 -21397
rect 15407 -21397 15487 -21387
rect 15407 -21407 15417 -21397
rect 15157 -21457 15417 -21407
rect 15477 -21457 15487 -21397
rect 15087 -21467 15487 -21457
rect 1 -21549 401 -21539
rect 1 -21609 11 -21549
rect 71 -21599 331 -21549
rect 71 -21609 81 -21599
rect 1 -21619 81 -21609
rect 321 -21609 331 -21599
rect 391 -21609 401 -21549
rect 321 -21619 401 -21609
rect 1 -21889 61 -21619
rect 331 -21629 401 -21619
rect 141 -21679 171 -21659
rect 121 -21719 171 -21679
rect 231 -21679 261 -21659
rect 231 -21719 281 -21679
rect 121 -21789 281 -21719
rect 121 -21829 171 -21789
rect 141 -21849 171 -21829
rect 231 -21829 281 -21789
rect 231 -21849 261 -21829
rect 341 -21889 401 -21629
rect 1 -21899 81 -21889
rect 1 -21959 11 -21899
rect 71 -21909 81 -21899
rect 321 -21899 401 -21889
rect 321 -21909 331 -21899
rect 71 -21959 331 -21909
rect 391 -21959 401 -21899
rect 1 -21969 401 -21959
rect 457 -21549 857 -21539
rect 457 -21609 467 -21549
rect 527 -21599 787 -21549
rect 527 -21609 537 -21599
rect 457 -21619 537 -21609
rect 777 -21609 787 -21599
rect 847 -21609 857 -21549
rect 777 -21619 857 -21609
rect 457 -21889 517 -21619
rect 787 -21629 857 -21619
rect 597 -21679 627 -21659
rect 577 -21719 627 -21679
rect 687 -21679 717 -21659
rect 687 -21719 737 -21679
rect 577 -21789 737 -21719
rect 577 -21829 627 -21789
rect 597 -21849 627 -21829
rect 687 -21829 737 -21789
rect 687 -21849 717 -21829
rect 797 -21889 857 -21629
rect 457 -21899 537 -21889
rect 457 -21959 467 -21899
rect 527 -21909 537 -21899
rect 777 -21899 857 -21889
rect 777 -21909 787 -21899
rect 527 -21959 787 -21909
rect 847 -21959 857 -21899
rect 457 -21969 857 -21959
rect 913 -21549 1313 -21539
rect 913 -21609 923 -21549
rect 983 -21599 1243 -21549
rect 983 -21609 993 -21599
rect 913 -21619 993 -21609
rect 1233 -21609 1243 -21599
rect 1303 -21609 1313 -21549
rect 1233 -21619 1313 -21609
rect 913 -21889 973 -21619
rect 1243 -21629 1313 -21619
rect 1053 -21679 1083 -21659
rect 1033 -21719 1083 -21679
rect 1143 -21679 1173 -21659
rect 1143 -21719 1193 -21679
rect 1033 -21789 1193 -21719
rect 1033 -21829 1083 -21789
rect 1053 -21849 1083 -21829
rect 1143 -21829 1193 -21789
rect 1143 -21849 1173 -21829
rect 1253 -21889 1313 -21629
rect 913 -21899 993 -21889
rect 913 -21959 923 -21899
rect 983 -21909 993 -21899
rect 1233 -21899 1313 -21889
rect 1233 -21909 1243 -21899
rect 983 -21959 1243 -21909
rect 1303 -21959 1313 -21899
rect 913 -21969 1313 -21959
rect 1371 -21549 1771 -21539
rect 1371 -21609 1381 -21549
rect 1441 -21599 1701 -21549
rect 1441 -21609 1451 -21599
rect 1371 -21619 1451 -21609
rect 1691 -21609 1701 -21599
rect 1761 -21609 1771 -21549
rect 1691 -21619 1771 -21609
rect 1371 -21889 1431 -21619
rect 1701 -21629 1771 -21619
rect 1511 -21679 1541 -21659
rect 1491 -21719 1541 -21679
rect 1601 -21679 1631 -21659
rect 1601 -21719 1651 -21679
rect 1491 -21789 1651 -21719
rect 1491 -21829 1541 -21789
rect 1511 -21849 1541 -21829
rect 1601 -21829 1651 -21789
rect 1601 -21849 1631 -21829
rect 1711 -21889 1771 -21629
rect 1371 -21899 1451 -21889
rect 1371 -21959 1381 -21899
rect 1441 -21909 1451 -21899
rect 1691 -21899 1771 -21889
rect 1691 -21909 1701 -21899
rect 1441 -21959 1701 -21909
rect 1761 -21959 1771 -21899
rect 1371 -21969 1771 -21959
rect 1827 -21549 2227 -21539
rect 1827 -21609 1837 -21549
rect 1897 -21599 2157 -21549
rect 1897 -21609 1907 -21599
rect 1827 -21619 1907 -21609
rect 2147 -21609 2157 -21599
rect 2217 -21609 2227 -21549
rect 2147 -21619 2227 -21609
rect 1827 -21889 1887 -21619
rect 2157 -21629 2227 -21619
rect 1967 -21679 1997 -21659
rect 1947 -21719 1997 -21679
rect 2057 -21679 2087 -21659
rect 2057 -21719 2107 -21679
rect 1947 -21789 2107 -21719
rect 1947 -21829 1997 -21789
rect 1967 -21849 1997 -21829
rect 2057 -21829 2107 -21789
rect 2057 -21849 2087 -21829
rect 2167 -21889 2227 -21629
rect 1827 -21899 1907 -21889
rect 1827 -21959 1837 -21899
rect 1897 -21909 1907 -21899
rect 2147 -21899 2227 -21889
rect 2147 -21909 2157 -21899
rect 1897 -21959 2157 -21909
rect 2217 -21959 2227 -21899
rect 1827 -21969 2227 -21959
rect 2283 -21549 2683 -21539
rect 2283 -21609 2293 -21549
rect 2353 -21599 2613 -21549
rect 2353 -21609 2363 -21599
rect 2283 -21619 2363 -21609
rect 2603 -21609 2613 -21599
rect 2673 -21609 2683 -21549
rect 2603 -21619 2683 -21609
rect 2283 -21889 2343 -21619
rect 2613 -21629 2683 -21619
rect 2423 -21679 2453 -21659
rect 2403 -21719 2453 -21679
rect 2513 -21679 2543 -21659
rect 2513 -21719 2563 -21679
rect 2403 -21789 2563 -21719
rect 2403 -21829 2453 -21789
rect 2423 -21849 2453 -21829
rect 2513 -21829 2563 -21789
rect 2513 -21849 2543 -21829
rect 2623 -21889 2683 -21629
rect 2283 -21899 2363 -21889
rect 2283 -21959 2293 -21899
rect 2353 -21909 2363 -21899
rect 2603 -21899 2683 -21889
rect 2603 -21909 2613 -21899
rect 2353 -21959 2613 -21909
rect 2673 -21959 2683 -21899
rect 2283 -21969 2683 -21959
rect 2741 -21549 3141 -21539
rect 2741 -21609 2751 -21549
rect 2811 -21599 3071 -21549
rect 2811 -21609 2821 -21599
rect 2741 -21619 2821 -21609
rect 3061 -21609 3071 -21599
rect 3131 -21609 3141 -21549
rect 3061 -21619 3141 -21609
rect 2741 -21889 2801 -21619
rect 3071 -21629 3141 -21619
rect 2881 -21679 2911 -21659
rect 2861 -21719 2911 -21679
rect 2971 -21679 3001 -21659
rect 2971 -21719 3021 -21679
rect 2861 -21789 3021 -21719
rect 2861 -21829 2911 -21789
rect 2881 -21849 2911 -21829
rect 2971 -21829 3021 -21789
rect 2971 -21849 3001 -21829
rect 3081 -21889 3141 -21629
rect 2741 -21899 2821 -21889
rect 2741 -21959 2751 -21899
rect 2811 -21909 2821 -21899
rect 3061 -21899 3141 -21889
rect 3061 -21909 3071 -21899
rect 2811 -21959 3071 -21909
rect 3131 -21959 3141 -21899
rect 2741 -21969 3141 -21959
rect 3197 -21549 3597 -21539
rect 3197 -21609 3207 -21549
rect 3267 -21599 3527 -21549
rect 3267 -21609 3277 -21599
rect 3197 -21619 3277 -21609
rect 3517 -21609 3527 -21599
rect 3587 -21609 3597 -21549
rect 3517 -21619 3597 -21609
rect 3197 -21889 3257 -21619
rect 3527 -21629 3597 -21619
rect 3337 -21679 3367 -21659
rect 3317 -21719 3367 -21679
rect 3427 -21679 3457 -21659
rect 3427 -21719 3477 -21679
rect 3317 -21789 3477 -21719
rect 3317 -21829 3367 -21789
rect 3337 -21849 3367 -21829
rect 3427 -21829 3477 -21789
rect 3427 -21849 3457 -21829
rect 3537 -21889 3597 -21629
rect 3197 -21899 3277 -21889
rect 3197 -21959 3207 -21899
rect 3267 -21909 3277 -21899
rect 3517 -21899 3597 -21889
rect 3517 -21909 3527 -21899
rect 3267 -21959 3527 -21909
rect 3587 -21959 3597 -21899
rect 3197 -21969 3597 -21959
rect 3653 -21549 4053 -21539
rect 3653 -21609 3663 -21549
rect 3723 -21599 3983 -21549
rect 3723 -21609 3733 -21599
rect 3653 -21619 3733 -21609
rect 3973 -21609 3983 -21599
rect 4043 -21609 4053 -21549
rect 3973 -21619 4053 -21609
rect 3653 -21889 3713 -21619
rect 3983 -21629 4053 -21619
rect 3793 -21679 3823 -21659
rect 3773 -21719 3823 -21679
rect 3883 -21679 3913 -21659
rect 3883 -21719 3933 -21679
rect 3773 -21789 3933 -21719
rect 3773 -21829 3823 -21789
rect 3793 -21849 3823 -21829
rect 3883 -21829 3933 -21789
rect 3883 -21849 3913 -21829
rect 3993 -21889 4053 -21629
rect 3653 -21899 3733 -21889
rect 3653 -21959 3663 -21899
rect 3723 -21909 3733 -21899
rect 3973 -21899 4053 -21889
rect 3973 -21909 3983 -21899
rect 3723 -21959 3983 -21909
rect 4043 -21959 4053 -21899
rect 3653 -21969 4053 -21959
rect 4111 -21549 4511 -21539
rect 4111 -21609 4121 -21549
rect 4181 -21599 4441 -21549
rect 4181 -21609 4191 -21599
rect 4111 -21619 4191 -21609
rect 4431 -21609 4441 -21599
rect 4501 -21609 4511 -21549
rect 4431 -21619 4511 -21609
rect 4111 -21889 4171 -21619
rect 4441 -21629 4511 -21619
rect 4251 -21679 4281 -21659
rect 4231 -21719 4281 -21679
rect 4341 -21679 4371 -21659
rect 4341 -21719 4391 -21679
rect 4231 -21789 4391 -21719
rect 4231 -21829 4281 -21789
rect 4251 -21849 4281 -21829
rect 4341 -21829 4391 -21789
rect 4341 -21849 4371 -21829
rect 4451 -21889 4511 -21629
rect 4111 -21899 4191 -21889
rect 4111 -21959 4121 -21899
rect 4181 -21909 4191 -21899
rect 4431 -21899 4511 -21889
rect 4431 -21909 4441 -21899
rect 4181 -21959 4441 -21909
rect 4501 -21959 4511 -21899
rect 4111 -21969 4511 -21959
rect 4567 -21549 4967 -21539
rect 4567 -21609 4577 -21549
rect 4637 -21599 4897 -21549
rect 4637 -21609 4647 -21599
rect 4567 -21619 4647 -21609
rect 4887 -21609 4897 -21599
rect 4957 -21609 4967 -21549
rect 4887 -21619 4967 -21609
rect 4567 -21889 4627 -21619
rect 4897 -21629 4967 -21619
rect 4707 -21679 4737 -21659
rect 4687 -21719 4737 -21679
rect 4797 -21679 4827 -21659
rect 4797 -21719 4847 -21679
rect 4687 -21789 4847 -21719
rect 4687 -21829 4737 -21789
rect 4707 -21849 4737 -21829
rect 4797 -21829 4847 -21789
rect 4797 -21849 4827 -21829
rect 4907 -21889 4967 -21629
rect 4567 -21899 4647 -21889
rect 4567 -21959 4577 -21899
rect 4637 -21909 4647 -21899
rect 4887 -21899 4967 -21889
rect 4887 -21909 4897 -21899
rect 4637 -21959 4897 -21909
rect 4957 -21959 4967 -21899
rect 4567 -21969 4967 -21959
rect 5023 -21549 5423 -21539
rect 5023 -21609 5033 -21549
rect 5093 -21599 5353 -21549
rect 5093 -21609 5103 -21599
rect 5023 -21619 5103 -21609
rect 5343 -21609 5353 -21599
rect 5413 -21609 5423 -21549
rect 5343 -21619 5423 -21609
rect 5023 -21889 5083 -21619
rect 5353 -21629 5423 -21619
rect 5163 -21679 5193 -21659
rect 5143 -21719 5193 -21679
rect 5253 -21679 5283 -21659
rect 5253 -21719 5303 -21679
rect 5143 -21789 5303 -21719
rect 5143 -21829 5193 -21789
rect 5163 -21849 5193 -21829
rect 5253 -21829 5303 -21789
rect 5253 -21849 5283 -21829
rect 5363 -21889 5423 -21629
rect 5023 -21899 5103 -21889
rect 5023 -21959 5033 -21899
rect 5093 -21909 5103 -21899
rect 5343 -21899 5423 -21889
rect 5343 -21909 5353 -21899
rect 5093 -21959 5353 -21909
rect 5413 -21959 5423 -21899
rect 5023 -21969 5423 -21959
rect 5481 -21549 5881 -21539
rect 5481 -21609 5491 -21549
rect 5551 -21599 5811 -21549
rect 5551 -21609 5561 -21599
rect 5481 -21619 5561 -21609
rect 5801 -21609 5811 -21599
rect 5871 -21609 5881 -21549
rect 5801 -21619 5881 -21609
rect 5481 -21889 5541 -21619
rect 5811 -21629 5881 -21619
rect 5621 -21679 5651 -21659
rect 5601 -21719 5651 -21679
rect 5711 -21679 5741 -21659
rect 5711 -21719 5761 -21679
rect 5601 -21789 5761 -21719
rect 5601 -21829 5651 -21789
rect 5621 -21849 5651 -21829
rect 5711 -21829 5761 -21789
rect 5711 -21849 5741 -21829
rect 5821 -21889 5881 -21629
rect 5481 -21899 5561 -21889
rect 5481 -21959 5491 -21899
rect 5551 -21909 5561 -21899
rect 5801 -21899 5881 -21889
rect 5801 -21909 5811 -21899
rect 5551 -21959 5811 -21909
rect 5871 -21959 5881 -21899
rect 5481 -21969 5881 -21959
rect 5937 -21549 6337 -21539
rect 5937 -21609 5947 -21549
rect 6007 -21599 6267 -21549
rect 6007 -21609 6017 -21599
rect 5937 -21619 6017 -21609
rect 6257 -21609 6267 -21599
rect 6327 -21609 6337 -21549
rect 6257 -21619 6337 -21609
rect 5937 -21889 5997 -21619
rect 6267 -21629 6337 -21619
rect 6077 -21679 6107 -21659
rect 6057 -21719 6107 -21679
rect 6167 -21679 6197 -21659
rect 6167 -21719 6217 -21679
rect 6057 -21789 6217 -21719
rect 6057 -21829 6107 -21789
rect 6077 -21849 6107 -21829
rect 6167 -21829 6217 -21789
rect 6167 -21849 6197 -21829
rect 6277 -21889 6337 -21629
rect 5937 -21899 6017 -21889
rect 5937 -21959 5947 -21899
rect 6007 -21909 6017 -21899
rect 6257 -21899 6337 -21889
rect 6257 -21909 6267 -21899
rect 6007 -21959 6267 -21909
rect 6327 -21959 6337 -21899
rect 5937 -21969 6337 -21959
rect 6393 -21549 6793 -21539
rect 6393 -21609 6403 -21549
rect 6463 -21599 6723 -21549
rect 6463 -21609 6473 -21599
rect 6393 -21619 6473 -21609
rect 6713 -21609 6723 -21599
rect 6783 -21609 6793 -21549
rect 6713 -21619 6793 -21609
rect 6393 -21889 6453 -21619
rect 6723 -21629 6793 -21619
rect 6533 -21679 6563 -21659
rect 6513 -21719 6563 -21679
rect 6623 -21679 6653 -21659
rect 6623 -21719 6673 -21679
rect 6513 -21789 6673 -21719
rect 6513 -21829 6563 -21789
rect 6533 -21849 6563 -21829
rect 6623 -21829 6673 -21789
rect 6623 -21849 6653 -21829
rect 6733 -21889 6793 -21629
rect 6393 -21899 6473 -21889
rect 6393 -21959 6403 -21899
rect 6463 -21909 6473 -21899
rect 6713 -21899 6793 -21889
rect 6713 -21909 6723 -21899
rect 6463 -21959 6723 -21909
rect 6783 -21959 6793 -21899
rect 6393 -21969 6793 -21959
rect 6851 -21549 7251 -21539
rect 6851 -21609 6861 -21549
rect 6921 -21599 7181 -21549
rect 6921 -21609 6931 -21599
rect 6851 -21619 6931 -21609
rect 7171 -21609 7181 -21599
rect 7241 -21609 7251 -21549
rect 7171 -21619 7251 -21609
rect 6851 -21889 6911 -21619
rect 7181 -21629 7251 -21619
rect 6991 -21679 7021 -21659
rect 6971 -21719 7021 -21679
rect 7081 -21679 7111 -21659
rect 7081 -21719 7131 -21679
rect 6971 -21789 7131 -21719
rect 6971 -21829 7021 -21789
rect 6991 -21849 7021 -21829
rect 7081 -21829 7131 -21789
rect 7081 -21849 7111 -21829
rect 7191 -21889 7251 -21629
rect 6851 -21899 6931 -21889
rect 6851 -21959 6861 -21899
rect 6921 -21909 6931 -21899
rect 7171 -21899 7251 -21889
rect 7171 -21909 7181 -21899
rect 6921 -21959 7181 -21909
rect 7241 -21959 7251 -21899
rect 6851 -21969 7251 -21959
rect 7307 -21549 7707 -21539
rect 7307 -21609 7317 -21549
rect 7377 -21599 7637 -21549
rect 7377 -21609 7387 -21599
rect 7307 -21619 7387 -21609
rect 7627 -21609 7637 -21599
rect 7697 -21609 7707 -21549
rect 7627 -21619 7707 -21609
rect 7307 -21889 7367 -21619
rect 7637 -21629 7707 -21619
rect 7447 -21679 7477 -21659
rect 7427 -21719 7477 -21679
rect 7537 -21679 7567 -21659
rect 7537 -21719 7587 -21679
rect 7427 -21789 7587 -21719
rect 7427 -21829 7477 -21789
rect 7447 -21849 7477 -21829
rect 7537 -21829 7587 -21789
rect 7537 -21849 7567 -21829
rect 7647 -21889 7707 -21629
rect 7307 -21899 7387 -21889
rect 7307 -21959 7317 -21899
rect 7377 -21909 7387 -21899
rect 7627 -21899 7707 -21889
rect 7627 -21909 7637 -21899
rect 7377 -21959 7637 -21909
rect 7697 -21959 7707 -21899
rect 7307 -21969 7707 -21959
rect 7763 -21549 8163 -21539
rect 7763 -21609 7773 -21549
rect 7833 -21599 8093 -21549
rect 7833 -21609 7843 -21599
rect 7763 -21619 7843 -21609
rect 8083 -21609 8093 -21599
rect 8153 -21609 8163 -21549
rect 8083 -21619 8163 -21609
rect 7763 -21889 7823 -21619
rect 8093 -21629 8163 -21619
rect 7903 -21679 7933 -21659
rect 7883 -21719 7933 -21679
rect 7993 -21679 8023 -21659
rect 7993 -21719 8043 -21679
rect 7883 -21789 8043 -21719
rect 7883 -21829 7933 -21789
rect 7903 -21849 7933 -21829
rect 7993 -21829 8043 -21789
rect 7993 -21849 8023 -21829
rect 8103 -21889 8163 -21629
rect 7763 -21899 7843 -21889
rect 7763 -21959 7773 -21899
rect 7833 -21909 7843 -21899
rect 8083 -21899 8163 -21889
rect 8083 -21909 8093 -21899
rect 7833 -21959 8093 -21909
rect 8153 -21959 8163 -21899
rect 7763 -21969 8163 -21959
rect 8237 -21549 8637 -21539
rect 8237 -21609 8247 -21549
rect 8307 -21599 8567 -21549
rect 8307 -21609 8317 -21599
rect 8237 -21619 8317 -21609
rect 8557 -21609 8567 -21599
rect 8627 -21609 8637 -21549
rect 8557 -21619 8637 -21609
rect 8237 -21889 8297 -21619
rect 8567 -21629 8637 -21619
rect 8377 -21679 8407 -21659
rect 8357 -21719 8407 -21679
rect 8467 -21679 8497 -21659
rect 8467 -21719 8517 -21679
rect 8357 -21789 8517 -21719
rect 8357 -21829 8407 -21789
rect 8377 -21849 8407 -21829
rect 8467 -21829 8517 -21789
rect 8467 -21849 8497 -21829
rect 8577 -21889 8637 -21629
rect 8237 -21899 8317 -21889
rect 8237 -21959 8247 -21899
rect 8307 -21909 8317 -21899
rect 8557 -21899 8637 -21889
rect 8557 -21909 8567 -21899
rect 8307 -21959 8567 -21909
rect 8627 -21959 8637 -21899
rect 8237 -21969 8637 -21959
rect 8693 -21549 9093 -21539
rect 8693 -21609 8703 -21549
rect 8763 -21599 9023 -21549
rect 8763 -21609 8773 -21599
rect 8693 -21619 8773 -21609
rect 9013 -21609 9023 -21599
rect 9083 -21609 9093 -21549
rect 9013 -21619 9093 -21609
rect 8693 -21889 8753 -21619
rect 9023 -21629 9093 -21619
rect 8833 -21679 8863 -21659
rect 8813 -21719 8863 -21679
rect 8923 -21679 8953 -21659
rect 8923 -21719 8973 -21679
rect 8813 -21789 8973 -21719
rect 8813 -21829 8863 -21789
rect 8833 -21849 8863 -21829
rect 8923 -21829 8973 -21789
rect 8923 -21849 8953 -21829
rect 9033 -21889 9093 -21629
rect 8693 -21899 8773 -21889
rect 8693 -21959 8703 -21899
rect 8763 -21909 8773 -21899
rect 9013 -21899 9093 -21889
rect 9013 -21909 9023 -21899
rect 8763 -21959 9023 -21909
rect 9083 -21959 9093 -21899
rect 8693 -21969 9093 -21959
rect 9151 -21549 9551 -21539
rect 9151 -21609 9161 -21549
rect 9221 -21599 9481 -21549
rect 9221 -21609 9231 -21599
rect 9151 -21619 9231 -21609
rect 9471 -21609 9481 -21599
rect 9541 -21609 9551 -21549
rect 9471 -21619 9551 -21609
rect 9151 -21889 9211 -21619
rect 9481 -21629 9551 -21619
rect 9291 -21679 9321 -21659
rect 9271 -21719 9321 -21679
rect 9381 -21679 9411 -21659
rect 9381 -21719 9431 -21679
rect 9271 -21789 9431 -21719
rect 9271 -21829 9321 -21789
rect 9291 -21849 9321 -21829
rect 9381 -21829 9431 -21789
rect 9381 -21849 9411 -21829
rect 9491 -21889 9551 -21629
rect 9151 -21899 9231 -21889
rect 9151 -21959 9161 -21899
rect 9221 -21909 9231 -21899
rect 9471 -21899 9551 -21889
rect 9471 -21909 9481 -21899
rect 9221 -21959 9481 -21909
rect 9541 -21959 9551 -21899
rect 9151 -21969 9551 -21959
rect 9607 -21549 10007 -21539
rect 9607 -21609 9617 -21549
rect 9677 -21599 9937 -21549
rect 9677 -21609 9687 -21599
rect 9607 -21619 9687 -21609
rect 9927 -21609 9937 -21599
rect 9997 -21609 10007 -21549
rect 9927 -21619 10007 -21609
rect 9607 -21889 9667 -21619
rect 9937 -21629 10007 -21619
rect 9747 -21679 9777 -21659
rect 9727 -21719 9777 -21679
rect 9837 -21679 9867 -21659
rect 9837 -21719 9887 -21679
rect 9727 -21789 9887 -21719
rect 9727 -21829 9777 -21789
rect 9747 -21849 9777 -21829
rect 9837 -21829 9887 -21789
rect 9837 -21849 9867 -21829
rect 9947 -21889 10007 -21629
rect 9607 -21899 9687 -21889
rect 9607 -21959 9617 -21899
rect 9677 -21909 9687 -21899
rect 9927 -21899 10007 -21889
rect 9927 -21909 9937 -21899
rect 9677 -21959 9937 -21909
rect 9997 -21959 10007 -21899
rect 9607 -21969 10007 -21959
rect 10063 -21549 10463 -21539
rect 10063 -21609 10073 -21549
rect 10133 -21599 10393 -21549
rect 10133 -21609 10143 -21599
rect 10063 -21619 10143 -21609
rect 10383 -21609 10393 -21599
rect 10453 -21609 10463 -21549
rect 10383 -21619 10463 -21609
rect 10063 -21889 10123 -21619
rect 10393 -21629 10463 -21619
rect 10203 -21679 10233 -21659
rect 10183 -21719 10233 -21679
rect 10293 -21679 10323 -21659
rect 10293 -21719 10343 -21679
rect 10183 -21789 10343 -21719
rect 10183 -21829 10233 -21789
rect 10203 -21849 10233 -21829
rect 10293 -21829 10343 -21789
rect 10293 -21849 10323 -21829
rect 10403 -21889 10463 -21629
rect 10063 -21899 10143 -21889
rect 10063 -21959 10073 -21899
rect 10133 -21909 10143 -21899
rect 10383 -21899 10463 -21889
rect 10383 -21909 10393 -21899
rect 10133 -21959 10393 -21909
rect 10453 -21959 10463 -21899
rect 10063 -21969 10463 -21959
rect 10521 -21549 10921 -21539
rect 10521 -21609 10531 -21549
rect 10591 -21599 10851 -21549
rect 10591 -21609 10601 -21599
rect 10521 -21619 10601 -21609
rect 10841 -21609 10851 -21599
rect 10911 -21609 10921 -21549
rect 10841 -21619 10921 -21609
rect 10521 -21889 10581 -21619
rect 10851 -21629 10921 -21619
rect 10661 -21679 10691 -21659
rect 10641 -21719 10691 -21679
rect 10751 -21679 10781 -21659
rect 10751 -21719 10801 -21679
rect 10641 -21789 10801 -21719
rect 10641 -21829 10691 -21789
rect 10661 -21849 10691 -21829
rect 10751 -21829 10801 -21789
rect 10751 -21849 10781 -21829
rect 10861 -21889 10921 -21629
rect 10521 -21899 10601 -21889
rect 10521 -21959 10531 -21899
rect 10591 -21909 10601 -21899
rect 10841 -21899 10921 -21889
rect 10841 -21909 10851 -21899
rect 10591 -21959 10851 -21909
rect 10911 -21959 10921 -21899
rect 10521 -21969 10921 -21959
rect 10977 -21549 11377 -21539
rect 10977 -21609 10987 -21549
rect 11047 -21599 11307 -21549
rect 11047 -21609 11057 -21599
rect 10977 -21619 11057 -21609
rect 11297 -21609 11307 -21599
rect 11367 -21609 11377 -21549
rect 11297 -21619 11377 -21609
rect 10977 -21889 11037 -21619
rect 11307 -21629 11377 -21619
rect 11117 -21679 11147 -21659
rect 11097 -21719 11147 -21679
rect 11207 -21679 11237 -21659
rect 11207 -21719 11257 -21679
rect 11097 -21789 11257 -21719
rect 11097 -21829 11147 -21789
rect 11117 -21849 11147 -21829
rect 11207 -21829 11257 -21789
rect 11207 -21849 11237 -21829
rect 11317 -21889 11377 -21629
rect 10977 -21899 11057 -21889
rect 10977 -21959 10987 -21899
rect 11047 -21909 11057 -21899
rect 11297 -21899 11377 -21889
rect 11297 -21909 11307 -21899
rect 11047 -21959 11307 -21909
rect 11367 -21959 11377 -21899
rect 10977 -21969 11377 -21959
rect 11433 -21549 11833 -21539
rect 11433 -21609 11443 -21549
rect 11503 -21599 11763 -21549
rect 11503 -21609 11513 -21599
rect 11433 -21619 11513 -21609
rect 11753 -21609 11763 -21599
rect 11823 -21609 11833 -21549
rect 11753 -21619 11833 -21609
rect 11433 -21889 11493 -21619
rect 11763 -21629 11833 -21619
rect 11573 -21679 11603 -21659
rect 11553 -21719 11603 -21679
rect 11663 -21679 11693 -21659
rect 11663 -21719 11713 -21679
rect 11553 -21789 11713 -21719
rect 11553 -21829 11603 -21789
rect 11573 -21849 11603 -21829
rect 11663 -21829 11713 -21789
rect 11663 -21849 11693 -21829
rect 11773 -21889 11833 -21629
rect 11433 -21899 11513 -21889
rect 11433 -21959 11443 -21899
rect 11503 -21909 11513 -21899
rect 11753 -21899 11833 -21889
rect 11753 -21909 11763 -21899
rect 11503 -21959 11763 -21909
rect 11823 -21959 11833 -21899
rect 11433 -21969 11833 -21959
rect 11891 -21549 12291 -21539
rect 11891 -21609 11901 -21549
rect 11961 -21599 12221 -21549
rect 11961 -21609 11971 -21599
rect 11891 -21619 11971 -21609
rect 12211 -21609 12221 -21599
rect 12281 -21609 12291 -21549
rect 12211 -21619 12291 -21609
rect 11891 -21889 11951 -21619
rect 12221 -21629 12291 -21619
rect 12031 -21679 12061 -21659
rect 12011 -21719 12061 -21679
rect 12121 -21679 12151 -21659
rect 12121 -21719 12171 -21679
rect 12011 -21789 12171 -21719
rect 12011 -21829 12061 -21789
rect 12031 -21849 12061 -21829
rect 12121 -21829 12171 -21789
rect 12121 -21849 12151 -21829
rect 12231 -21889 12291 -21629
rect 11891 -21899 11971 -21889
rect 11891 -21959 11901 -21899
rect 11961 -21909 11971 -21899
rect 12211 -21899 12291 -21889
rect 12211 -21909 12221 -21899
rect 11961 -21959 12221 -21909
rect 12281 -21959 12291 -21899
rect 11891 -21969 12291 -21959
rect 12347 -21549 12747 -21539
rect 12347 -21609 12357 -21549
rect 12417 -21599 12677 -21549
rect 12417 -21609 12427 -21599
rect 12347 -21619 12427 -21609
rect 12667 -21609 12677 -21599
rect 12737 -21609 12747 -21549
rect 12667 -21619 12747 -21609
rect 12347 -21889 12407 -21619
rect 12677 -21629 12747 -21619
rect 12487 -21679 12517 -21659
rect 12467 -21719 12517 -21679
rect 12577 -21679 12607 -21659
rect 12577 -21719 12627 -21679
rect 12467 -21789 12627 -21719
rect 12467 -21829 12517 -21789
rect 12487 -21849 12517 -21829
rect 12577 -21829 12627 -21789
rect 12577 -21849 12607 -21829
rect 12687 -21889 12747 -21629
rect 12347 -21899 12427 -21889
rect 12347 -21959 12357 -21899
rect 12417 -21909 12427 -21899
rect 12667 -21899 12747 -21889
rect 12667 -21909 12677 -21899
rect 12417 -21959 12677 -21909
rect 12737 -21959 12747 -21899
rect 12347 -21969 12747 -21959
rect 12803 -21549 13203 -21539
rect 12803 -21609 12813 -21549
rect 12873 -21599 13133 -21549
rect 12873 -21609 12883 -21599
rect 12803 -21619 12883 -21609
rect 13123 -21609 13133 -21599
rect 13193 -21609 13203 -21549
rect 13123 -21619 13203 -21609
rect 12803 -21889 12863 -21619
rect 13133 -21629 13203 -21619
rect 12943 -21679 12973 -21659
rect 12923 -21719 12973 -21679
rect 13033 -21679 13063 -21659
rect 13033 -21719 13083 -21679
rect 12923 -21789 13083 -21719
rect 12923 -21829 12973 -21789
rect 12943 -21849 12973 -21829
rect 13033 -21829 13083 -21789
rect 13033 -21849 13063 -21829
rect 13143 -21889 13203 -21629
rect 12803 -21899 12883 -21889
rect 12803 -21959 12813 -21899
rect 12873 -21909 12883 -21899
rect 13123 -21899 13203 -21889
rect 13123 -21909 13133 -21899
rect 12873 -21959 13133 -21909
rect 13193 -21959 13203 -21899
rect 12803 -21969 13203 -21959
rect 13261 -21549 13661 -21539
rect 13261 -21609 13271 -21549
rect 13331 -21599 13591 -21549
rect 13331 -21609 13341 -21599
rect 13261 -21619 13341 -21609
rect 13581 -21609 13591 -21599
rect 13651 -21609 13661 -21549
rect 13581 -21619 13661 -21609
rect 13261 -21889 13321 -21619
rect 13591 -21629 13661 -21619
rect 13401 -21679 13431 -21659
rect 13381 -21719 13431 -21679
rect 13491 -21679 13521 -21659
rect 13491 -21719 13541 -21679
rect 13381 -21789 13541 -21719
rect 13381 -21829 13431 -21789
rect 13401 -21849 13431 -21829
rect 13491 -21829 13541 -21789
rect 13491 -21849 13521 -21829
rect 13601 -21889 13661 -21629
rect 13261 -21899 13341 -21889
rect 13261 -21959 13271 -21899
rect 13331 -21909 13341 -21899
rect 13581 -21899 13661 -21889
rect 13581 -21909 13591 -21899
rect 13331 -21959 13591 -21909
rect 13651 -21959 13661 -21899
rect 13261 -21969 13661 -21959
rect 13717 -21549 14117 -21539
rect 13717 -21609 13727 -21549
rect 13787 -21599 14047 -21549
rect 13787 -21609 13797 -21599
rect 13717 -21619 13797 -21609
rect 14037 -21609 14047 -21599
rect 14107 -21609 14117 -21549
rect 14037 -21619 14117 -21609
rect 13717 -21889 13777 -21619
rect 14047 -21629 14117 -21619
rect 13857 -21679 13887 -21659
rect 13837 -21719 13887 -21679
rect 13947 -21679 13977 -21659
rect 13947 -21719 13997 -21679
rect 13837 -21789 13997 -21719
rect 13837 -21829 13887 -21789
rect 13857 -21849 13887 -21829
rect 13947 -21829 13997 -21789
rect 13947 -21849 13977 -21829
rect 14057 -21889 14117 -21629
rect 13717 -21899 13797 -21889
rect 13717 -21959 13727 -21899
rect 13787 -21909 13797 -21899
rect 14037 -21899 14117 -21889
rect 14037 -21909 14047 -21899
rect 13787 -21959 14047 -21909
rect 14107 -21959 14117 -21899
rect 13717 -21969 14117 -21959
rect 14173 -21549 14573 -21539
rect 14173 -21609 14183 -21549
rect 14243 -21599 14503 -21549
rect 14243 -21609 14253 -21599
rect 14173 -21619 14253 -21609
rect 14493 -21609 14503 -21599
rect 14563 -21609 14573 -21549
rect 14493 -21619 14573 -21609
rect 14173 -21889 14233 -21619
rect 14503 -21629 14573 -21619
rect 14313 -21679 14343 -21659
rect 14293 -21719 14343 -21679
rect 14403 -21679 14433 -21659
rect 14403 -21719 14453 -21679
rect 14293 -21789 14453 -21719
rect 14293 -21829 14343 -21789
rect 14313 -21849 14343 -21829
rect 14403 -21829 14453 -21789
rect 14403 -21849 14433 -21829
rect 14513 -21889 14573 -21629
rect 14173 -21899 14253 -21889
rect 14173 -21959 14183 -21899
rect 14243 -21909 14253 -21899
rect 14493 -21899 14573 -21889
rect 14493 -21909 14503 -21899
rect 14243 -21959 14503 -21909
rect 14563 -21959 14573 -21899
rect 14173 -21969 14573 -21959
rect 14631 -21549 15031 -21539
rect 14631 -21609 14641 -21549
rect 14701 -21599 14961 -21549
rect 14701 -21609 14711 -21599
rect 14631 -21619 14711 -21609
rect 14951 -21609 14961 -21599
rect 15021 -21609 15031 -21549
rect 14951 -21619 15031 -21609
rect 14631 -21889 14691 -21619
rect 14961 -21629 15031 -21619
rect 14771 -21679 14801 -21659
rect 14751 -21719 14801 -21679
rect 14861 -21679 14891 -21659
rect 14861 -21719 14911 -21679
rect 14751 -21789 14911 -21719
rect 14751 -21829 14801 -21789
rect 14771 -21849 14801 -21829
rect 14861 -21829 14911 -21789
rect 14861 -21849 14891 -21829
rect 14971 -21889 15031 -21629
rect 14631 -21899 14711 -21889
rect 14631 -21959 14641 -21899
rect 14701 -21909 14711 -21899
rect 14951 -21899 15031 -21889
rect 14951 -21909 14961 -21899
rect 14701 -21959 14961 -21909
rect 15021 -21959 15031 -21899
rect 14631 -21969 15031 -21959
rect 15087 -21549 15487 -21539
rect 15087 -21609 15097 -21549
rect 15157 -21599 15417 -21549
rect 15157 -21609 15167 -21599
rect 15087 -21619 15167 -21609
rect 15407 -21609 15417 -21599
rect 15477 -21609 15487 -21549
rect 15407 -21619 15487 -21609
rect 15087 -21889 15147 -21619
rect 15417 -21629 15487 -21619
rect 15227 -21679 15257 -21659
rect 15207 -21719 15257 -21679
rect 15317 -21679 15347 -21659
rect 15317 -21719 15367 -21679
rect 15207 -21789 15367 -21719
rect 15207 -21829 15257 -21789
rect 15227 -21849 15257 -21829
rect 15317 -21829 15367 -21789
rect 15317 -21849 15347 -21829
rect 15427 -21889 15487 -21629
rect 15087 -21899 15167 -21889
rect 15087 -21959 15097 -21899
rect 15157 -21909 15167 -21899
rect 15407 -21899 15487 -21889
rect 15407 -21909 15417 -21899
rect 15157 -21959 15417 -21909
rect 15477 -21959 15487 -21899
rect 15087 -21969 15487 -21959
rect 1 -22041 401 -22031
rect 1 -22101 11 -22041
rect 71 -22091 331 -22041
rect 71 -22101 81 -22091
rect 1 -22111 81 -22101
rect 321 -22101 331 -22091
rect 391 -22101 401 -22041
rect 321 -22111 401 -22101
rect 1 -22381 61 -22111
rect 331 -22121 401 -22111
rect 141 -22171 171 -22151
rect 121 -22211 171 -22171
rect 231 -22171 261 -22151
rect 231 -22211 281 -22171
rect 121 -22281 281 -22211
rect 121 -22321 171 -22281
rect 141 -22341 171 -22321
rect 231 -22321 281 -22281
rect 231 -22341 261 -22321
rect 341 -22381 401 -22121
rect 1 -22391 81 -22381
rect 1 -22451 11 -22391
rect 71 -22401 81 -22391
rect 321 -22391 401 -22381
rect 321 -22401 331 -22391
rect 71 -22451 331 -22401
rect 391 -22451 401 -22391
rect 1 -22461 401 -22451
rect 457 -22041 857 -22031
rect 457 -22101 467 -22041
rect 527 -22091 787 -22041
rect 527 -22101 537 -22091
rect 457 -22111 537 -22101
rect 777 -22101 787 -22091
rect 847 -22101 857 -22041
rect 777 -22111 857 -22101
rect 457 -22381 517 -22111
rect 787 -22121 857 -22111
rect 597 -22171 627 -22151
rect 577 -22211 627 -22171
rect 687 -22171 717 -22151
rect 687 -22211 737 -22171
rect 577 -22281 737 -22211
rect 577 -22321 627 -22281
rect 597 -22341 627 -22321
rect 687 -22321 737 -22281
rect 687 -22341 717 -22321
rect 797 -22381 857 -22121
rect 457 -22391 537 -22381
rect 457 -22451 467 -22391
rect 527 -22401 537 -22391
rect 777 -22391 857 -22381
rect 777 -22401 787 -22391
rect 527 -22451 787 -22401
rect 847 -22451 857 -22391
rect 457 -22461 857 -22451
rect 913 -22041 1313 -22031
rect 913 -22101 923 -22041
rect 983 -22091 1243 -22041
rect 983 -22101 993 -22091
rect 913 -22111 993 -22101
rect 1233 -22101 1243 -22091
rect 1303 -22101 1313 -22041
rect 1233 -22111 1313 -22101
rect 913 -22381 973 -22111
rect 1243 -22121 1313 -22111
rect 1053 -22171 1083 -22151
rect 1033 -22211 1083 -22171
rect 1143 -22171 1173 -22151
rect 1143 -22211 1193 -22171
rect 1033 -22281 1193 -22211
rect 1033 -22321 1083 -22281
rect 1053 -22341 1083 -22321
rect 1143 -22321 1193 -22281
rect 1143 -22341 1173 -22321
rect 1253 -22381 1313 -22121
rect 913 -22391 993 -22381
rect 913 -22451 923 -22391
rect 983 -22401 993 -22391
rect 1233 -22391 1313 -22381
rect 1233 -22401 1243 -22391
rect 983 -22451 1243 -22401
rect 1303 -22451 1313 -22391
rect 913 -22461 1313 -22451
rect 1371 -22041 1771 -22031
rect 1371 -22101 1381 -22041
rect 1441 -22091 1701 -22041
rect 1441 -22101 1451 -22091
rect 1371 -22111 1451 -22101
rect 1691 -22101 1701 -22091
rect 1761 -22101 1771 -22041
rect 1691 -22111 1771 -22101
rect 1371 -22381 1431 -22111
rect 1701 -22121 1771 -22111
rect 1511 -22171 1541 -22151
rect 1491 -22211 1541 -22171
rect 1601 -22171 1631 -22151
rect 1601 -22211 1651 -22171
rect 1491 -22281 1651 -22211
rect 1491 -22321 1541 -22281
rect 1511 -22341 1541 -22321
rect 1601 -22321 1651 -22281
rect 1601 -22341 1631 -22321
rect 1711 -22381 1771 -22121
rect 1371 -22391 1451 -22381
rect 1371 -22451 1381 -22391
rect 1441 -22401 1451 -22391
rect 1691 -22391 1771 -22381
rect 1691 -22401 1701 -22391
rect 1441 -22451 1701 -22401
rect 1761 -22451 1771 -22391
rect 1371 -22461 1771 -22451
rect 1827 -22041 2227 -22031
rect 1827 -22101 1837 -22041
rect 1897 -22091 2157 -22041
rect 1897 -22101 1907 -22091
rect 1827 -22111 1907 -22101
rect 2147 -22101 2157 -22091
rect 2217 -22101 2227 -22041
rect 2147 -22111 2227 -22101
rect 1827 -22381 1887 -22111
rect 2157 -22121 2227 -22111
rect 1967 -22171 1997 -22151
rect 1947 -22211 1997 -22171
rect 2057 -22171 2087 -22151
rect 2057 -22211 2107 -22171
rect 1947 -22281 2107 -22211
rect 1947 -22321 1997 -22281
rect 1967 -22341 1997 -22321
rect 2057 -22321 2107 -22281
rect 2057 -22341 2087 -22321
rect 2167 -22381 2227 -22121
rect 1827 -22391 1907 -22381
rect 1827 -22451 1837 -22391
rect 1897 -22401 1907 -22391
rect 2147 -22391 2227 -22381
rect 2147 -22401 2157 -22391
rect 1897 -22451 2157 -22401
rect 2217 -22451 2227 -22391
rect 1827 -22461 2227 -22451
rect 2283 -22041 2683 -22031
rect 2283 -22101 2293 -22041
rect 2353 -22091 2613 -22041
rect 2353 -22101 2363 -22091
rect 2283 -22111 2363 -22101
rect 2603 -22101 2613 -22091
rect 2673 -22101 2683 -22041
rect 2603 -22111 2683 -22101
rect 2283 -22381 2343 -22111
rect 2613 -22121 2683 -22111
rect 2423 -22171 2453 -22151
rect 2403 -22211 2453 -22171
rect 2513 -22171 2543 -22151
rect 2513 -22211 2563 -22171
rect 2403 -22281 2563 -22211
rect 2403 -22321 2453 -22281
rect 2423 -22341 2453 -22321
rect 2513 -22321 2563 -22281
rect 2513 -22341 2543 -22321
rect 2623 -22381 2683 -22121
rect 2283 -22391 2363 -22381
rect 2283 -22451 2293 -22391
rect 2353 -22401 2363 -22391
rect 2603 -22391 2683 -22381
rect 2603 -22401 2613 -22391
rect 2353 -22451 2613 -22401
rect 2673 -22451 2683 -22391
rect 2283 -22461 2683 -22451
rect 2741 -22041 3141 -22031
rect 2741 -22101 2751 -22041
rect 2811 -22091 3071 -22041
rect 2811 -22101 2821 -22091
rect 2741 -22111 2821 -22101
rect 3061 -22101 3071 -22091
rect 3131 -22101 3141 -22041
rect 3061 -22111 3141 -22101
rect 2741 -22381 2801 -22111
rect 3071 -22121 3141 -22111
rect 2881 -22171 2911 -22151
rect 2861 -22211 2911 -22171
rect 2971 -22171 3001 -22151
rect 2971 -22211 3021 -22171
rect 2861 -22281 3021 -22211
rect 2861 -22321 2911 -22281
rect 2881 -22341 2911 -22321
rect 2971 -22321 3021 -22281
rect 2971 -22341 3001 -22321
rect 3081 -22381 3141 -22121
rect 2741 -22391 2821 -22381
rect 2741 -22451 2751 -22391
rect 2811 -22401 2821 -22391
rect 3061 -22391 3141 -22381
rect 3061 -22401 3071 -22391
rect 2811 -22451 3071 -22401
rect 3131 -22451 3141 -22391
rect 2741 -22461 3141 -22451
rect 3197 -22041 3597 -22031
rect 3197 -22101 3207 -22041
rect 3267 -22091 3527 -22041
rect 3267 -22101 3277 -22091
rect 3197 -22111 3277 -22101
rect 3517 -22101 3527 -22091
rect 3587 -22101 3597 -22041
rect 3517 -22111 3597 -22101
rect 3197 -22381 3257 -22111
rect 3527 -22121 3597 -22111
rect 3337 -22171 3367 -22151
rect 3317 -22211 3367 -22171
rect 3427 -22171 3457 -22151
rect 3427 -22211 3477 -22171
rect 3317 -22281 3477 -22211
rect 3317 -22321 3367 -22281
rect 3337 -22341 3367 -22321
rect 3427 -22321 3477 -22281
rect 3427 -22341 3457 -22321
rect 3537 -22381 3597 -22121
rect 3197 -22391 3277 -22381
rect 3197 -22451 3207 -22391
rect 3267 -22401 3277 -22391
rect 3517 -22391 3597 -22381
rect 3517 -22401 3527 -22391
rect 3267 -22451 3527 -22401
rect 3587 -22451 3597 -22391
rect 3197 -22461 3597 -22451
rect 3653 -22041 4053 -22031
rect 3653 -22101 3663 -22041
rect 3723 -22091 3983 -22041
rect 3723 -22101 3733 -22091
rect 3653 -22111 3733 -22101
rect 3973 -22101 3983 -22091
rect 4043 -22101 4053 -22041
rect 3973 -22111 4053 -22101
rect 3653 -22381 3713 -22111
rect 3983 -22121 4053 -22111
rect 3793 -22171 3823 -22151
rect 3773 -22211 3823 -22171
rect 3883 -22171 3913 -22151
rect 3883 -22211 3933 -22171
rect 3773 -22281 3933 -22211
rect 3773 -22321 3823 -22281
rect 3793 -22341 3823 -22321
rect 3883 -22321 3933 -22281
rect 3883 -22341 3913 -22321
rect 3993 -22381 4053 -22121
rect 3653 -22391 3733 -22381
rect 3653 -22451 3663 -22391
rect 3723 -22401 3733 -22391
rect 3973 -22391 4053 -22381
rect 3973 -22401 3983 -22391
rect 3723 -22451 3983 -22401
rect 4043 -22451 4053 -22391
rect 3653 -22461 4053 -22451
rect 4111 -22041 4511 -22031
rect 4111 -22101 4121 -22041
rect 4181 -22091 4441 -22041
rect 4181 -22101 4191 -22091
rect 4111 -22111 4191 -22101
rect 4431 -22101 4441 -22091
rect 4501 -22101 4511 -22041
rect 4431 -22111 4511 -22101
rect 4111 -22381 4171 -22111
rect 4441 -22121 4511 -22111
rect 4251 -22171 4281 -22151
rect 4231 -22211 4281 -22171
rect 4341 -22171 4371 -22151
rect 4341 -22211 4391 -22171
rect 4231 -22281 4391 -22211
rect 4231 -22321 4281 -22281
rect 4251 -22341 4281 -22321
rect 4341 -22321 4391 -22281
rect 4341 -22341 4371 -22321
rect 4451 -22381 4511 -22121
rect 4111 -22391 4191 -22381
rect 4111 -22451 4121 -22391
rect 4181 -22401 4191 -22391
rect 4431 -22391 4511 -22381
rect 4431 -22401 4441 -22391
rect 4181 -22451 4441 -22401
rect 4501 -22451 4511 -22391
rect 4111 -22461 4511 -22451
rect 4567 -22041 4967 -22031
rect 4567 -22101 4577 -22041
rect 4637 -22091 4897 -22041
rect 4637 -22101 4647 -22091
rect 4567 -22111 4647 -22101
rect 4887 -22101 4897 -22091
rect 4957 -22101 4967 -22041
rect 4887 -22111 4967 -22101
rect 4567 -22381 4627 -22111
rect 4897 -22121 4967 -22111
rect 4707 -22171 4737 -22151
rect 4687 -22211 4737 -22171
rect 4797 -22171 4827 -22151
rect 4797 -22211 4847 -22171
rect 4687 -22281 4847 -22211
rect 4687 -22321 4737 -22281
rect 4707 -22341 4737 -22321
rect 4797 -22321 4847 -22281
rect 4797 -22341 4827 -22321
rect 4907 -22381 4967 -22121
rect 4567 -22391 4647 -22381
rect 4567 -22451 4577 -22391
rect 4637 -22401 4647 -22391
rect 4887 -22391 4967 -22381
rect 4887 -22401 4897 -22391
rect 4637 -22451 4897 -22401
rect 4957 -22451 4967 -22391
rect 4567 -22461 4967 -22451
rect 5023 -22041 5423 -22031
rect 5023 -22101 5033 -22041
rect 5093 -22091 5353 -22041
rect 5093 -22101 5103 -22091
rect 5023 -22111 5103 -22101
rect 5343 -22101 5353 -22091
rect 5413 -22101 5423 -22041
rect 5343 -22111 5423 -22101
rect 5023 -22381 5083 -22111
rect 5353 -22121 5423 -22111
rect 5163 -22171 5193 -22151
rect 5143 -22211 5193 -22171
rect 5253 -22171 5283 -22151
rect 5253 -22211 5303 -22171
rect 5143 -22281 5303 -22211
rect 5143 -22321 5193 -22281
rect 5163 -22341 5193 -22321
rect 5253 -22321 5303 -22281
rect 5253 -22341 5283 -22321
rect 5363 -22381 5423 -22121
rect 5023 -22391 5103 -22381
rect 5023 -22451 5033 -22391
rect 5093 -22401 5103 -22391
rect 5343 -22391 5423 -22381
rect 5343 -22401 5353 -22391
rect 5093 -22451 5353 -22401
rect 5413 -22451 5423 -22391
rect 5023 -22461 5423 -22451
rect 5481 -22041 5881 -22031
rect 5481 -22101 5491 -22041
rect 5551 -22091 5811 -22041
rect 5551 -22101 5561 -22091
rect 5481 -22111 5561 -22101
rect 5801 -22101 5811 -22091
rect 5871 -22101 5881 -22041
rect 5801 -22111 5881 -22101
rect 5481 -22381 5541 -22111
rect 5811 -22121 5881 -22111
rect 5621 -22171 5651 -22151
rect 5601 -22211 5651 -22171
rect 5711 -22171 5741 -22151
rect 5711 -22211 5761 -22171
rect 5601 -22281 5761 -22211
rect 5601 -22321 5651 -22281
rect 5621 -22341 5651 -22321
rect 5711 -22321 5761 -22281
rect 5711 -22341 5741 -22321
rect 5821 -22381 5881 -22121
rect 5481 -22391 5561 -22381
rect 5481 -22451 5491 -22391
rect 5551 -22401 5561 -22391
rect 5801 -22391 5881 -22381
rect 5801 -22401 5811 -22391
rect 5551 -22451 5811 -22401
rect 5871 -22451 5881 -22391
rect 5481 -22461 5881 -22451
rect 5937 -22041 6337 -22031
rect 5937 -22101 5947 -22041
rect 6007 -22091 6267 -22041
rect 6007 -22101 6017 -22091
rect 5937 -22111 6017 -22101
rect 6257 -22101 6267 -22091
rect 6327 -22101 6337 -22041
rect 6257 -22111 6337 -22101
rect 5937 -22381 5997 -22111
rect 6267 -22121 6337 -22111
rect 6077 -22171 6107 -22151
rect 6057 -22211 6107 -22171
rect 6167 -22171 6197 -22151
rect 6167 -22211 6217 -22171
rect 6057 -22281 6217 -22211
rect 6057 -22321 6107 -22281
rect 6077 -22341 6107 -22321
rect 6167 -22321 6217 -22281
rect 6167 -22341 6197 -22321
rect 6277 -22381 6337 -22121
rect 5937 -22391 6017 -22381
rect 5937 -22451 5947 -22391
rect 6007 -22401 6017 -22391
rect 6257 -22391 6337 -22381
rect 6257 -22401 6267 -22391
rect 6007 -22451 6267 -22401
rect 6327 -22451 6337 -22391
rect 5937 -22461 6337 -22451
rect 6393 -22041 6793 -22031
rect 6393 -22101 6403 -22041
rect 6463 -22091 6723 -22041
rect 6463 -22101 6473 -22091
rect 6393 -22111 6473 -22101
rect 6713 -22101 6723 -22091
rect 6783 -22101 6793 -22041
rect 6713 -22111 6793 -22101
rect 6393 -22381 6453 -22111
rect 6723 -22121 6793 -22111
rect 6533 -22171 6563 -22151
rect 6513 -22211 6563 -22171
rect 6623 -22171 6653 -22151
rect 6623 -22211 6673 -22171
rect 6513 -22281 6673 -22211
rect 6513 -22321 6563 -22281
rect 6533 -22341 6563 -22321
rect 6623 -22321 6673 -22281
rect 6623 -22341 6653 -22321
rect 6733 -22381 6793 -22121
rect 6393 -22391 6473 -22381
rect 6393 -22451 6403 -22391
rect 6463 -22401 6473 -22391
rect 6713 -22391 6793 -22381
rect 6713 -22401 6723 -22391
rect 6463 -22451 6723 -22401
rect 6783 -22451 6793 -22391
rect 6393 -22461 6793 -22451
rect 6851 -22041 7251 -22031
rect 6851 -22101 6861 -22041
rect 6921 -22091 7181 -22041
rect 6921 -22101 6931 -22091
rect 6851 -22111 6931 -22101
rect 7171 -22101 7181 -22091
rect 7241 -22101 7251 -22041
rect 7171 -22111 7251 -22101
rect 6851 -22381 6911 -22111
rect 7181 -22121 7251 -22111
rect 6991 -22171 7021 -22151
rect 6971 -22211 7021 -22171
rect 7081 -22171 7111 -22151
rect 7081 -22211 7131 -22171
rect 6971 -22281 7131 -22211
rect 6971 -22321 7021 -22281
rect 6991 -22341 7021 -22321
rect 7081 -22321 7131 -22281
rect 7081 -22341 7111 -22321
rect 7191 -22381 7251 -22121
rect 6851 -22391 6931 -22381
rect 6851 -22451 6861 -22391
rect 6921 -22401 6931 -22391
rect 7171 -22391 7251 -22381
rect 7171 -22401 7181 -22391
rect 6921 -22451 7181 -22401
rect 7241 -22451 7251 -22391
rect 6851 -22461 7251 -22451
rect 7307 -22041 7707 -22031
rect 7307 -22101 7317 -22041
rect 7377 -22091 7637 -22041
rect 7377 -22101 7387 -22091
rect 7307 -22111 7387 -22101
rect 7627 -22101 7637 -22091
rect 7697 -22101 7707 -22041
rect 7627 -22111 7707 -22101
rect 7307 -22381 7367 -22111
rect 7637 -22121 7707 -22111
rect 7447 -22171 7477 -22151
rect 7427 -22211 7477 -22171
rect 7537 -22171 7567 -22151
rect 7537 -22211 7587 -22171
rect 7427 -22281 7587 -22211
rect 7427 -22321 7477 -22281
rect 7447 -22341 7477 -22321
rect 7537 -22321 7587 -22281
rect 7537 -22341 7567 -22321
rect 7647 -22381 7707 -22121
rect 7307 -22391 7387 -22381
rect 7307 -22451 7317 -22391
rect 7377 -22401 7387 -22391
rect 7627 -22391 7707 -22381
rect 7627 -22401 7637 -22391
rect 7377 -22451 7637 -22401
rect 7697 -22451 7707 -22391
rect 7307 -22461 7707 -22451
rect 7763 -22041 8163 -22031
rect 7763 -22101 7773 -22041
rect 7833 -22091 8093 -22041
rect 7833 -22101 7843 -22091
rect 7763 -22111 7843 -22101
rect 8083 -22101 8093 -22091
rect 8153 -22101 8163 -22041
rect 8083 -22111 8163 -22101
rect 7763 -22381 7823 -22111
rect 8093 -22121 8163 -22111
rect 7903 -22171 7933 -22151
rect 7883 -22211 7933 -22171
rect 7993 -22171 8023 -22151
rect 7993 -22211 8043 -22171
rect 7883 -22281 8043 -22211
rect 7883 -22321 7933 -22281
rect 7903 -22341 7933 -22321
rect 7993 -22321 8043 -22281
rect 7993 -22341 8023 -22321
rect 8103 -22381 8163 -22121
rect 7763 -22391 7843 -22381
rect 7763 -22451 7773 -22391
rect 7833 -22401 7843 -22391
rect 8083 -22391 8163 -22381
rect 8083 -22401 8093 -22391
rect 7833 -22451 8093 -22401
rect 8153 -22451 8163 -22391
rect 7763 -22461 8163 -22451
rect 8237 -22041 8637 -22031
rect 8237 -22101 8247 -22041
rect 8307 -22091 8567 -22041
rect 8307 -22101 8317 -22091
rect 8237 -22111 8317 -22101
rect 8557 -22101 8567 -22091
rect 8627 -22101 8637 -22041
rect 8557 -22111 8637 -22101
rect 8237 -22381 8297 -22111
rect 8567 -22121 8637 -22111
rect 8377 -22171 8407 -22151
rect 8357 -22211 8407 -22171
rect 8467 -22171 8497 -22151
rect 8467 -22211 8517 -22171
rect 8357 -22281 8517 -22211
rect 8357 -22321 8407 -22281
rect 8377 -22341 8407 -22321
rect 8467 -22321 8517 -22281
rect 8467 -22341 8497 -22321
rect 8577 -22381 8637 -22121
rect 8237 -22391 8317 -22381
rect 8237 -22451 8247 -22391
rect 8307 -22401 8317 -22391
rect 8557 -22391 8637 -22381
rect 8557 -22401 8567 -22391
rect 8307 -22451 8567 -22401
rect 8627 -22451 8637 -22391
rect 8237 -22461 8637 -22451
rect 8693 -22041 9093 -22031
rect 8693 -22101 8703 -22041
rect 8763 -22091 9023 -22041
rect 8763 -22101 8773 -22091
rect 8693 -22111 8773 -22101
rect 9013 -22101 9023 -22091
rect 9083 -22101 9093 -22041
rect 9013 -22111 9093 -22101
rect 8693 -22381 8753 -22111
rect 9023 -22121 9093 -22111
rect 8833 -22171 8863 -22151
rect 8813 -22211 8863 -22171
rect 8923 -22171 8953 -22151
rect 8923 -22211 8973 -22171
rect 8813 -22281 8973 -22211
rect 8813 -22321 8863 -22281
rect 8833 -22341 8863 -22321
rect 8923 -22321 8973 -22281
rect 8923 -22341 8953 -22321
rect 9033 -22381 9093 -22121
rect 8693 -22391 8773 -22381
rect 8693 -22451 8703 -22391
rect 8763 -22401 8773 -22391
rect 9013 -22391 9093 -22381
rect 9013 -22401 9023 -22391
rect 8763 -22451 9023 -22401
rect 9083 -22451 9093 -22391
rect 8693 -22461 9093 -22451
rect 9151 -22041 9551 -22031
rect 9151 -22101 9161 -22041
rect 9221 -22091 9481 -22041
rect 9221 -22101 9231 -22091
rect 9151 -22111 9231 -22101
rect 9471 -22101 9481 -22091
rect 9541 -22101 9551 -22041
rect 9471 -22111 9551 -22101
rect 9151 -22381 9211 -22111
rect 9481 -22121 9551 -22111
rect 9291 -22171 9321 -22151
rect 9271 -22211 9321 -22171
rect 9381 -22171 9411 -22151
rect 9381 -22211 9431 -22171
rect 9271 -22281 9431 -22211
rect 9271 -22321 9321 -22281
rect 9291 -22341 9321 -22321
rect 9381 -22321 9431 -22281
rect 9381 -22341 9411 -22321
rect 9491 -22381 9551 -22121
rect 9151 -22391 9231 -22381
rect 9151 -22451 9161 -22391
rect 9221 -22401 9231 -22391
rect 9471 -22391 9551 -22381
rect 9471 -22401 9481 -22391
rect 9221 -22451 9481 -22401
rect 9541 -22451 9551 -22391
rect 9151 -22461 9551 -22451
rect 9607 -22041 10007 -22031
rect 9607 -22101 9617 -22041
rect 9677 -22091 9937 -22041
rect 9677 -22101 9687 -22091
rect 9607 -22111 9687 -22101
rect 9927 -22101 9937 -22091
rect 9997 -22101 10007 -22041
rect 9927 -22111 10007 -22101
rect 9607 -22381 9667 -22111
rect 9937 -22121 10007 -22111
rect 9747 -22171 9777 -22151
rect 9727 -22211 9777 -22171
rect 9837 -22171 9867 -22151
rect 9837 -22211 9887 -22171
rect 9727 -22281 9887 -22211
rect 9727 -22321 9777 -22281
rect 9747 -22341 9777 -22321
rect 9837 -22321 9887 -22281
rect 9837 -22341 9867 -22321
rect 9947 -22381 10007 -22121
rect 9607 -22391 9687 -22381
rect 9607 -22451 9617 -22391
rect 9677 -22401 9687 -22391
rect 9927 -22391 10007 -22381
rect 9927 -22401 9937 -22391
rect 9677 -22451 9937 -22401
rect 9997 -22451 10007 -22391
rect 9607 -22461 10007 -22451
rect 10063 -22041 10463 -22031
rect 10063 -22101 10073 -22041
rect 10133 -22091 10393 -22041
rect 10133 -22101 10143 -22091
rect 10063 -22111 10143 -22101
rect 10383 -22101 10393 -22091
rect 10453 -22101 10463 -22041
rect 10383 -22111 10463 -22101
rect 10063 -22381 10123 -22111
rect 10393 -22121 10463 -22111
rect 10203 -22171 10233 -22151
rect 10183 -22211 10233 -22171
rect 10293 -22171 10323 -22151
rect 10293 -22211 10343 -22171
rect 10183 -22281 10343 -22211
rect 10183 -22321 10233 -22281
rect 10203 -22341 10233 -22321
rect 10293 -22321 10343 -22281
rect 10293 -22341 10323 -22321
rect 10403 -22381 10463 -22121
rect 10063 -22391 10143 -22381
rect 10063 -22451 10073 -22391
rect 10133 -22401 10143 -22391
rect 10383 -22391 10463 -22381
rect 10383 -22401 10393 -22391
rect 10133 -22451 10393 -22401
rect 10453 -22451 10463 -22391
rect 10063 -22461 10463 -22451
rect 10521 -22041 10921 -22031
rect 10521 -22101 10531 -22041
rect 10591 -22091 10851 -22041
rect 10591 -22101 10601 -22091
rect 10521 -22111 10601 -22101
rect 10841 -22101 10851 -22091
rect 10911 -22101 10921 -22041
rect 10841 -22111 10921 -22101
rect 10521 -22381 10581 -22111
rect 10851 -22121 10921 -22111
rect 10661 -22171 10691 -22151
rect 10641 -22211 10691 -22171
rect 10751 -22171 10781 -22151
rect 10751 -22211 10801 -22171
rect 10641 -22281 10801 -22211
rect 10641 -22321 10691 -22281
rect 10661 -22341 10691 -22321
rect 10751 -22321 10801 -22281
rect 10751 -22341 10781 -22321
rect 10861 -22381 10921 -22121
rect 10521 -22391 10601 -22381
rect 10521 -22451 10531 -22391
rect 10591 -22401 10601 -22391
rect 10841 -22391 10921 -22381
rect 10841 -22401 10851 -22391
rect 10591 -22451 10851 -22401
rect 10911 -22451 10921 -22391
rect 10521 -22461 10921 -22451
rect 10977 -22041 11377 -22031
rect 10977 -22101 10987 -22041
rect 11047 -22091 11307 -22041
rect 11047 -22101 11057 -22091
rect 10977 -22111 11057 -22101
rect 11297 -22101 11307 -22091
rect 11367 -22101 11377 -22041
rect 11297 -22111 11377 -22101
rect 10977 -22381 11037 -22111
rect 11307 -22121 11377 -22111
rect 11117 -22171 11147 -22151
rect 11097 -22211 11147 -22171
rect 11207 -22171 11237 -22151
rect 11207 -22211 11257 -22171
rect 11097 -22281 11257 -22211
rect 11097 -22321 11147 -22281
rect 11117 -22341 11147 -22321
rect 11207 -22321 11257 -22281
rect 11207 -22341 11237 -22321
rect 11317 -22381 11377 -22121
rect 10977 -22391 11057 -22381
rect 10977 -22451 10987 -22391
rect 11047 -22401 11057 -22391
rect 11297 -22391 11377 -22381
rect 11297 -22401 11307 -22391
rect 11047 -22451 11307 -22401
rect 11367 -22451 11377 -22391
rect 10977 -22461 11377 -22451
rect 11433 -22041 11833 -22031
rect 11433 -22101 11443 -22041
rect 11503 -22091 11763 -22041
rect 11503 -22101 11513 -22091
rect 11433 -22111 11513 -22101
rect 11753 -22101 11763 -22091
rect 11823 -22101 11833 -22041
rect 11753 -22111 11833 -22101
rect 11433 -22381 11493 -22111
rect 11763 -22121 11833 -22111
rect 11573 -22171 11603 -22151
rect 11553 -22211 11603 -22171
rect 11663 -22171 11693 -22151
rect 11663 -22211 11713 -22171
rect 11553 -22281 11713 -22211
rect 11553 -22321 11603 -22281
rect 11573 -22341 11603 -22321
rect 11663 -22321 11713 -22281
rect 11663 -22341 11693 -22321
rect 11773 -22381 11833 -22121
rect 11433 -22391 11513 -22381
rect 11433 -22451 11443 -22391
rect 11503 -22401 11513 -22391
rect 11753 -22391 11833 -22381
rect 11753 -22401 11763 -22391
rect 11503 -22451 11763 -22401
rect 11823 -22451 11833 -22391
rect 11433 -22461 11833 -22451
rect 11891 -22041 12291 -22031
rect 11891 -22101 11901 -22041
rect 11961 -22091 12221 -22041
rect 11961 -22101 11971 -22091
rect 11891 -22111 11971 -22101
rect 12211 -22101 12221 -22091
rect 12281 -22101 12291 -22041
rect 12211 -22111 12291 -22101
rect 11891 -22381 11951 -22111
rect 12221 -22121 12291 -22111
rect 12031 -22171 12061 -22151
rect 12011 -22211 12061 -22171
rect 12121 -22171 12151 -22151
rect 12121 -22211 12171 -22171
rect 12011 -22281 12171 -22211
rect 12011 -22321 12061 -22281
rect 12031 -22341 12061 -22321
rect 12121 -22321 12171 -22281
rect 12121 -22341 12151 -22321
rect 12231 -22381 12291 -22121
rect 11891 -22391 11971 -22381
rect 11891 -22451 11901 -22391
rect 11961 -22401 11971 -22391
rect 12211 -22391 12291 -22381
rect 12211 -22401 12221 -22391
rect 11961 -22451 12221 -22401
rect 12281 -22451 12291 -22391
rect 11891 -22461 12291 -22451
rect 12347 -22041 12747 -22031
rect 12347 -22101 12357 -22041
rect 12417 -22091 12677 -22041
rect 12417 -22101 12427 -22091
rect 12347 -22111 12427 -22101
rect 12667 -22101 12677 -22091
rect 12737 -22101 12747 -22041
rect 12667 -22111 12747 -22101
rect 12347 -22381 12407 -22111
rect 12677 -22121 12747 -22111
rect 12487 -22171 12517 -22151
rect 12467 -22211 12517 -22171
rect 12577 -22171 12607 -22151
rect 12577 -22211 12627 -22171
rect 12467 -22281 12627 -22211
rect 12467 -22321 12517 -22281
rect 12487 -22341 12517 -22321
rect 12577 -22321 12627 -22281
rect 12577 -22341 12607 -22321
rect 12687 -22381 12747 -22121
rect 12347 -22391 12427 -22381
rect 12347 -22451 12357 -22391
rect 12417 -22401 12427 -22391
rect 12667 -22391 12747 -22381
rect 12667 -22401 12677 -22391
rect 12417 -22451 12677 -22401
rect 12737 -22451 12747 -22391
rect 12347 -22461 12747 -22451
rect 12803 -22041 13203 -22031
rect 12803 -22101 12813 -22041
rect 12873 -22091 13133 -22041
rect 12873 -22101 12883 -22091
rect 12803 -22111 12883 -22101
rect 13123 -22101 13133 -22091
rect 13193 -22101 13203 -22041
rect 13123 -22111 13203 -22101
rect 12803 -22381 12863 -22111
rect 13133 -22121 13203 -22111
rect 12943 -22171 12973 -22151
rect 12923 -22211 12973 -22171
rect 13033 -22171 13063 -22151
rect 13033 -22211 13083 -22171
rect 12923 -22281 13083 -22211
rect 12923 -22321 12973 -22281
rect 12943 -22341 12973 -22321
rect 13033 -22321 13083 -22281
rect 13033 -22341 13063 -22321
rect 13143 -22381 13203 -22121
rect 12803 -22391 12883 -22381
rect 12803 -22451 12813 -22391
rect 12873 -22401 12883 -22391
rect 13123 -22391 13203 -22381
rect 13123 -22401 13133 -22391
rect 12873 -22451 13133 -22401
rect 13193 -22451 13203 -22391
rect 12803 -22461 13203 -22451
rect 13261 -22041 13661 -22031
rect 13261 -22101 13271 -22041
rect 13331 -22091 13591 -22041
rect 13331 -22101 13341 -22091
rect 13261 -22111 13341 -22101
rect 13581 -22101 13591 -22091
rect 13651 -22101 13661 -22041
rect 13581 -22111 13661 -22101
rect 13261 -22381 13321 -22111
rect 13591 -22121 13661 -22111
rect 13401 -22171 13431 -22151
rect 13381 -22211 13431 -22171
rect 13491 -22171 13521 -22151
rect 13491 -22211 13541 -22171
rect 13381 -22281 13541 -22211
rect 13381 -22321 13431 -22281
rect 13401 -22341 13431 -22321
rect 13491 -22321 13541 -22281
rect 13491 -22341 13521 -22321
rect 13601 -22381 13661 -22121
rect 13261 -22391 13341 -22381
rect 13261 -22451 13271 -22391
rect 13331 -22401 13341 -22391
rect 13581 -22391 13661 -22381
rect 13581 -22401 13591 -22391
rect 13331 -22451 13591 -22401
rect 13651 -22451 13661 -22391
rect 13261 -22461 13661 -22451
rect 13717 -22041 14117 -22031
rect 13717 -22101 13727 -22041
rect 13787 -22091 14047 -22041
rect 13787 -22101 13797 -22091
rect 13717 -22111 13797 -22101
rect 14037 -22101 14047 -22091
rect 14107 -22101 14117 -22041
rect 14037 -22111 14117 -22101
rect 13717 -22381 13777 -22111
rect 14047 -22121 14117 -22111
rect 13857 -22171 13887 -22151
rect 13837 -22211 13887 -22171
rect 13947 -22171 13977 -22151
rect 13947 -22211 13997 -22171
rect 13837 -22281 13997 -22211
rect 13837 -22321 13887 -22281
rect 13857 -22341 13887 -22321
rect 13947 -22321 13997 -22281
rect 13947 -22341 13977 -22321
rect 14057 -22381 14117 -22121
rect 13717 -22391 13797 -22381
rect 13717 -22451 13727 -22391
rect 13787 -22401 13797 -22391
rect 14037 -22391 14117 -22381
rect 14037 -22401 14047 -22391
rect 13787 -22451 14047 -22401
rect 14107 -22451 14117 -22391
rect 13717 -22461 14117 -22451
rect 14173 -22041 14573 -22031
rect 14173 -22101 14183 -22041
rect 14243 -22091 14503 -22041
rect 14243 -22101 14253 -22091
rect 14173 -22111 14253 -22101
rect 14493 -22101 14503 -22091
rect 14563 -22101 14573 -22041
rect 14493 -22111 14573 -22101
rect 14173 -22381 14233 -22111
rect 14503 -22121 14573 -22111
rect 14313 -22171 14343 -22151
rect 14293 -22211 14343 -22171
rect 14403 -22171 14433 -22151
rect 14403 -22211 14453 -22171
rect 14293 -22281 14453 -22211
rect 14293 -22321 14343 -22281
rect 14313 -22341 14343 -22321
rect 14403 -22321 14453 -22281
rect 14403 -22341 14433 -22321
rect 14513 -22381 14573 -22121
rect 14173 -22391 14253 -22381
rect 14173 -22451 14183 -22391
rect 14243 -22401 14253 -22391
rect 14493 -22391 14573 -22381
rect 14493 -22401 14503 -22391
rect 14243 -22451 14503 -22401
rect 14563 -22451 14573 -22391
rect 14173 -22461 14573 -22451
rect 14631 -22041 15031 -22031
rect 14631 -22101 14641 -22041
rect 14701 -22091 14961 -22041
rect 14701 -22101 14711 -22091
rect 14631 -22111 14711 -22101
rect 14951 -22101 14961 -22091
rect 15021 -22101 15031 -22041
rect 14951 -22111 15031 -22101
rect 14631 -22381 14691 -22111
rect 14961 -22121 15031 -22111
rect 14771 -22171 14801 -22151
rect 14751 -22211 14801 -22171
rect 14861 -22171 14891 -22151
rect 14861 -22211 14911 -22171
rect 14751 -22281 14911 -22211
rect 14751 -22321 14801 -22281
rect 14771 -22341 14801 -22321
rect 14861 -22321 14911 -22281
rect 14861 -22341 14891 -22321
rect 14971 -22381 15031 -22121
rect 14631 -22391 14711 -22381
rect 14631 -22451 14641 -22391
rect 14701 -22401 14711 -22391
rect 14951 -22391 15031 -22381
rect 14951 -22401 14961 -22391
rect 14701 -22451 14961 -22401
rect 15021 -22451 15031 -22391
rect 14631 -22461 15031 -22451
rect 15087 -22041 15487 -22031
rect 15087 -22101 15097 -22041
rect 15157 -22091 15417 -22041
rect 15157 -22101 15167 -22091
rect 15087 -22111 15167 -22101
rect 15407 -22101 15417 -22091
rect 15477 -22101 15487 -22041
rect 15407 -22111 15487 -22101
rect 15087 -22381 15147 -22111
rect 15417 -22121 15487 -22111
rect 15227 -22171 15257 -22151
rect 15207 -22211 15257 -22171
rect 15317 -22171 15347 -22151
rect 15317 -22211 15367 -22171
rect 15207 -22281 15367 -22211
rect 15207 -22321 15257 -22281
rect 15227 -22341 15257 -22321
rect 15317 -22321 15367 -22281
rect 15317 -22341 15347 -22321
rect 15427 -22381 15487 -22121
rect 15087 -22391 15167 -22381
rect 15087 -22451 15097 -22391
rect 15157 -22401 15167 -22391
rect 15407 -22391 15487 -22381
rect 15407 -22401 15417 -22391
rect 15157 -22451 15417 -22401
rect 15477 -22451 15487 -22391
rect 15087 -22461 15487 -22451
rect 1 -22528 401 -22518
rect 1 -22588 11 -22528
rect 71 -22578 331 -22528
rect 71 -22588 81 -22578
rect 1 -22598 81 -22588
rect 321 -22588 331 -22578
rect 391 -22588 401 -22528
rect 321 -22598 401 -22588
rect 1 -22868 61 -22598
rect 141 -22658 171 -22638
rect 121 -22698 171 -22658
rect 231 -22658 261 -22638
rect 231 -22698 281 -22658
rect 121 -22768 281 -22698
rect 121 -22808 171 -22768
rect 141 -22828 171 -22808
rect 231 -22808 281 -22768
rect 231 -22828 261 -22808
rect 341 -22858 401 -22598
rect 331 -22868 401 -22858
rect 1 -22878 81 -22868
rect 1 -22938 11 -22878
rect 71 -22888 81 -22878
rect 321 -22878 401 -22868
rect 321 -22888 331 -22878
rect 71 -22938 331 -22888
rect 391 -22938 401 -22878
rect 1 -22948 401 -22938
rect 457 -22528 857 -22518
rect 457 -22588 467 -22528
rect 527 -22578 787 -22528
rect 527 -22588 537 -22578
rect 457 -22598 537 -22588
rect 777 -22588 787 -22578
rect 847 -22588 857 -22528
rect 777 -22598 857 -22588
rect 457 -22868 517 -22598
rect 597 -22658 627 -22638
rect 577 -22698 627 -22658
rect 687 -22658 717 -22638
rect 687 -22698 737 -22658
rect 577 -22768 737 -22698
rect 577 -22808 627 -22768
rect 597 -22828 627 -22808
rect 687 -22808 737 -22768
rect 687 -22828 717 -22808
rect 797 -22858 857 -22598
rect 787 -22868 857 -22858
rect 457 -22878 537 -22868
rect 457 -22938 467 -22878
rect 527 -22888 537 -22878
rect 777 -22878 857 -22868
rect 777 -22888 787 -22878
rect 527 -22938 787 -22888
rect 847 -22938 857 -22878
rect 457 -22948 857 -22938
rect 913 -22528 1313 -22518
rect 913 -22588 923 -22528
rect 983 -22578 1243 -22528
rect 983 -22588 993 -22578
rect 913 -22598 993 -22588
rect 1233 -22588 1243 -22578
rect 1303 -22588 1313 -22528
rect 1233 -22598 1313 -22588
rect 913 -22868 973 -22598
rect 1053 -22658 1083 -22638
rect 1033 -22698 1083 -22658
rect 1143 -22658 1173 -22638
rect 1143 -22698 1193 -22658
rect 1033 -22768 1193 -22698
rect 1033 -22808 1083 -22768
rect 1053 -22828 1083 -22808
rect 1143 -22808 1193 -22768
rect 1143 -22828 1173 -22808
rect 1253 -22858 1313 -22598
rect 1243 -22868 1313 -22858
rect 913 -22878 993 -22868
rect 913 -22938 923 -22878
rect 983 -22888 993 -22878
rect 1233 -22878 1313 -22868
rect 1233 -22888 1243 -22878
rect 983 -22938 1243 -22888
rect 1303 -22938 1313 -22878
rect 913 -22948 1313 -22938
rect 1371 -22528 1771 -22518
rect 1371 -22588 1381 -22528
rect 1441 -22578 1701 -22528
rect 1441 -22588 1451 -22578
rect 1371 -22598 1451 -22588
rect 1691 -22588 1701 -22578
rect 1761 -22588 1771 -22528
rect 1691 -22598 1771 -22588
rect 1371 -22868 1431 -22598
rect 1511 -22658 1541 -22638
rect 1491 -22698 1541 -22658
rect 1601 -22658 1631 -22638
rect 1601 -22698 1651 -22658
rect 1491 -22768 1651 -22698
rect 1491 -22808 1541 -22768
rect 1511 -22828 1541 -22808
rect 1601 -22808 1651 -22768
rect 1601 -22828 1631 -22808
rect 1711 -22858 1771 -22598
rect 1701 -22868 1771 -22858
rect 1371 -22878 1451 -22868
rect 1371 -22938 1381 -22878
rect 1441 -22888 1451 -22878
rect 1691 -22878 1771 -22868
rect 1691 -22888 1701 -22878
rect 1441 -22938 1701 -22888
rect 1761 -22938 1771 -22878
rect 1371 -22948 1771 -22938
rect 1827 -22528 2227 -22518
rect 1827 -22588 1837 -22528
rect 1897 -22578 2157 -22528
rect 1897 -22588 1907 -22578
rect 1827 -22598 1907 -22588
rect 2147 -22588 2157 -22578
rect 2217 -22588 2227 -22528
rect 2147 -22598 2227 -22588
rect 1827 -22868 1887 -22598
rect 1967 -22658 1997 -22638
rect 1947 -22698 1997 -22658
rect 2057 -22658 2087 -22638
rect 2057 -22698 2107 -22658
rect 1947 -22768 2107 -22698
rect 1947 -22808 1997 -22768
rect 1967 -22828 1997 -22808
rect 2057 -22808 2107 -22768
rect 2057 -22828 2087 -22808
rect 2167 -22858 2227 -22598
rect 2157 -22868 2227 -22858
rect 1827 -22878 1907 -22868
rect 1827 -22938 1837 -22878
rect 1897 -22888 1907 -22878
rect 2147 -22878 2227 -22868
rect 2147 -22888 2157 -22878
rect 1897 -22938 2157 -22888
rect 2217 -22938 2227 -22878
rect 1827 -22948 2227 -22938
rect 2283 -22528 2683 -22518
rect 2283 -22588 2293 -22528
rect 2353 -22578 2613 -22528
rect 2353 -22588 2363 -22578
rect 2283 -22598 2363 -22588
rect 2603 -22588 2613 -22578
rect 2673 -22588 2683 -22528
rect 2603 -22598 2683 -22588
rect 2283 -22868 2343 -22598
rect 2423 -22658 2453 -22638
rect 2403 -22698 2453 -22658
rect 2513 -22658 2543 -22638
rect 2513 -22698 2563 -22658
rect 2403 -22768 2563 -22698
rect 2403 -22808 2453 -22768
rect 2423 -22828 2453 -22808
rect 2513 -22808 2563 -22768
rect 2513 -22828 2543 -22808
rect 2623 -22858 2683 -22598
rect 2613 -22868 2683 -22858
rect 2283 -22878 2363 -22868
rect 2283 -22938 2293 -22878
rect 2353 -22888 2363 -22878
rect 2603 -22878 2683 -22868
rect 2603 -22888 2613 -22878
rect 2353 -22938 2613 -22888
rect 2673 -22938 2683 -22878
rect 2283 -22948 2683 -22938
rect 2741 -22528 3141 -22518
rect 2741 -22588 2751 -22528
rect 2811 -22578 3071 -22528
rect 2811 -22588 2821 -22578
rect 2741 -22598 2821 -22588
rect 3061 -22588 3071 -22578
rect 3131 -22588 3141 -22528
rect 3061 -22598 3141 -22588
rect 2741 -22868 2801 -22598
rect 2881 -22658 2911 -22638
rect 2861 -22698 2911 -22658
rect 2971 -22658 3001 -22638
rect 2971 -22698 3021 -22658
rect 2861 -22768 3021 -22698
rect 2861 -22808 2911 -22768
rect 2881 -22828 2911 -22808
rect 2971 -22808 3021 -22768
rect 2971 -22828 3001 -22808
rect 3081 -22858 3141 -22598
rect 3071 -22868 3141 -22858
rect 2741 -22878 2821 -22868
rect 2741 -22938 2751 -22878
rect 2811 -22888 2821 -22878
rect 3061 -22878 3141 -22868
rect 3061 -22888 3071 -22878
rect 2811 -22938 3071 -22888
rect 3131 -22938 3141 -22878
rect 2741 -22948 3141 -22938
rect 3197 -22528 3597 -22518
rect 3197 -22588 3207 -22528
rect 3267 -22578 3527 -22528
rect 3267 -22588 3277 -22578
rect 3197 -22598 3277 -22588
rect 3517 -22588 3527 -22578
rect 3587 -22588 3597 -22528
rect 3517 -22598 3597 -22588
rect 3197 -22868 3257 -22598
rect 3337 -22658 3367 -22638
rect 3317 -22698 3367 -22658
rect 3427 -22658 3457 -22638
rect 3427 -22698 3477 -22658
rect 3317 -22768 3477 -22698
rect 3317 -22808 3367 -22768
rect 3337 -22828 3367 -22808
rect 3427 -22808 3477 -22768
rect 3427 -22828 3457 -22808
rect 3537 -22858 3597 -22598
rect 3527 -22868 3597 -22858
rect 3197 -22878 3277 -22868
rect 3197 -22938 3207 -22878
rect 3267 -22888 3277 -22878
rect 3517 -22878 3597 -22868
rect 3517 -22888 3527 -22878
rect 3267 -22938 3527 -22888
rect 3587 -22938 3597 -22878
rect 3197 -22948 3597 -22938
rect 3653 -22528 4053 -22518
rect 3653 -22588 3663 -22528
rect 3723 -22578 3983 -22528
rect 3723 -22588 3733 -22578
rect 3653 -22598 3733 -22588
rect 3973 -22588 3983 -22578
rect 4043 -22588 4053 -22528
rect 3973 -22598 4053 -22588
rect 3653 -22868 3713 -22598
rect 3793 -22658 3823 -22638
rect 3773 -22698 3823 -22658
rect 3883 -22658 3913 -22638
rect 3883 -22698 3933 -22658
rect 3773 -22768 3933 -22698
rect 3773 -22808 3823 -22768
rect 3793 -22828 3823 -22808
rect 3883 -22808 3933 -22768
rect 3883 -22828 3913 -22808
rect 3993 -22858 4053 -22598
rect 3983 -22868 4053 -22858
rect 3653 -22878 3733 -22868
rect 3653 -22938 3663 -22878
rect 3723 -22888 3733 -22878
rect 3973 -22878 4053 -22868
rect 3973 -22888 3983 -22878
rect 3723 -22938 3983 -22888
rect 4043 -22938 4053 -22878
rect 3653 -22948 4053 -22938
rect 4111 -22528 4511 -22518
rect 4111 -22588 4121 -22528
rect 4181 -22578 4441 -22528
rect 4181 -22588 4191 -22578
rect 4111 -22598 4191 -22588
rect 4431 -22588 4441 -22578
rect 4501 -22588 4511 -22528
rect 4431 -22598 4511 -22588
rect 4111 -22868 4171 -22598
rect 4251 -22658 4281 -22638
rect 4231 -22698 4281 -22658
rect 4341 -22658 4371 -22638
rect 4341 -22698 4391 -22658
rect 4231 -22768 4391 -22698
rect 4231 -22808 4281 -22768
rect 4251 -22828 4281 -22808
rect 4341 -22808 4391 -22768
rect 4341 -22828 4371 -22808
rect 4451 -22858 4511 -22598
rect 4441 -22868 4511 -22858
rect 4111 -22878 4191 -22868
rect 4111 -22938 4121 -22878
rect 4181 -22888 4191 -22878
rect 4431 -22878 4511 -22868
rect 4431 -22888 4441 -22878
rect 4181 -22938 4441 -22888
rect 4501 -22938 4511 -22878
rect 4111 -22948 4511 -22938
rect 4567 -22528 4967 -22518
rect 4567 -22588 4577 -22528
rect 4637 -22578 4897 -22528
rect 4637 -22588 4647 -22578
rect 4567 -22598 4647 -22588
rect 4887 -22588 4897 -22578
rect 4957 -22588 4967 -22528
rect 4887 -22598 4967 -22588
rect 4567 -22868 4627 -22598
rect 4707 -22658 4737 -22638
rect 4687 -22698 4737 -22658
rect 4797 -22658 4827 -22638
rect 4797 -22698 4847 -22658
rect 4687 -22768 4847 -22698
rect 4687 -22808 4737 -22768
rect 4707 -22828 4737 -22808
rect 4797 -22808 4847 -22768
rect 4797 -22828 4827 -22808
rect 4907 -22858 4967 -22598
rect 4897 -22868 4967 -22858
rect 4567 -22878 4647 -22868
rect 4567 -22938 4577 -22878
rect 4637 -22888 4647 -22878
rect 4887 -22878 4967 -22868
rect 4887 -22888 4897 -22878
rect 4637 -22938 4897 -22888
rect 4957 -22938 4967 -22878
rect 4567 -22948 4967 -22938
rect 5023 -22528 5423 -22518
rect 5023 -22588 5033 -22528
rect 5093 -22578 5353 -22528
rect 5093 -22588 5103 -22578
rect 5023 -22598 5103 -22588
rect 5343 -22588 5353 -22578
rect 5413 -22588 5423 -22528
rect 5343 -22598 5423 -22588
rect 5023 -22868 5083 -22598
rect 5163 -22658 5193 -22638
rect 5143 -22698 5193 -22658
rect 5253 -22658 5283 -22638
rect 5253 -22698 5303 -22658
rect 5143 -22768 5303 -22698
rect 5143 -22808 5193 -22768
rect 5163 -22828 5193 -22808
rect 5253 -22808 5303 -22768
rect 5253 -22828 5283 -22808
rect 5363 -22858 5423 -22598
rect 5353 -22868 5423 -22858
rect 5023 -22878 5103 -22868
rect 5023 -22938 5033 -22878
rect 5093 -22888 5103 -22878
rect 5343 -22878 5423 -22868
rect 5343 -22888 5353 -22878
rect 5093 -22938 5353 -22888
rect 5413 -22938 5423 -22878
rect 5023 -22948 5423 -22938
rect 5481 -22528 5881 -22518
rect 5481 -22588 5491 -22528
rect 5551 -22578 5811 -22528
rect 5551 -22588 5561 -22578
rect 5481 -22598 5561 -22588
rect 5801 -22588 5811 -22578
rect 5871 -22588 5881 -22528
rect 5801 -22598 5881 -22588
rect 5481 -22868 5541 -22598
rect 5621 -22658 5651 -22638
rect 5601 -22698 5651 -22658
rect 5711 -22658 5741 -22638
rect 5711 -22698 5761 -22658
rect 5601 -22768 5761 -22698
rect 5601 -22808 5651 -22768
rect 5621 -22828 5651 -22808
rect 5711 -22808 5761 -22768
rect 5711 -22828 5741 -22808
rect 5821 -22858 5881 -22598
rect 5811 -22868 5881 -22858
rect 5481 -22878 5561 -22868
rect 5481 -22938 5491 -22878
rect 5551 -22888 5561 -22878
rect 5801 -22878 5881 -22868
rect 5801 -22888 5811 -22878
rect 5551 -22938 5811 -22888
rect 5871 -22938 5881 -22878
rect 5481 -22948 5881 -22938
rect 5937 -22528 6337 -22518
rect 5937 -22588 5947 -22528
rect 6007 -22578 6267 -22528
rect 6007 -22588 6017 -22578
rect 5937 -22598 6017 -22588
rect 6257 -22588 6267 -22578
rect 6327 -22588 6337 -22528
rect 6257 -22598 6337 -22588
rect 5937 -22868 5997 -22598
rect 6077 -22658 6107 -22638
rect 6057 -22698 6107 -22658
rect 6167 -22658 6197 -22638
rect 6167 -22698 6217 -22658
rect 6057 -22768 6217 -22698
rect 6057 -22808 6107 -22768
rect 6077 -22828 6107 -22808
rect 6167 -22808 6217 -22768
rect 6167 -22828 6197 -22808
rect 6277 -22858 6337 -22598
rect 6267 -22868 6337 -22858
rect 5937 -22878 6017 -22868
rect 5937 -22938 5947 -22878
rect 6007 -22888 6017 -22878
rect 6257 -22878 6337 -22868
rect 6257 -22888 6267 -22878
rect 6007 -22938 6267 -22888
rect 6327 -22938 6337 -22878
rect 5937 -22948 6337 -22938
rect 6393 -22528 6793 -22518
rect 6393 -22588 6403 -22528
rect 6463 -22578 6723 -22528
rect 6463 -22588 6473 -22578
rect 6393 -22598 6473 -22588
rect 6713 -22588 6723 -22578
rect 6783 -22588 6793 -22528
rect 6713 -22598 6793 -22588
rect 6393 -22868 6453 -22598
rect 6533 -22658 6563 -22638
rect 6513 -22698 6563 -22658
rect 6623 -22658 6653 -22638
rect 6623 -22698 6673 -22658
rect 6513 -22768 6673 -22698
rect 6513 -22808 6563 -22768
rect 6533 -22828 6563 -22808
rect 6623 -22808 6673 -22768
rect 6623 -22828 6653 -22808
rect 6733 -22858 6793 -22598
rect 6723 -22868 6793 -22858
rect 6393 -22878 6473 -22868
rect 6393 -22938 6403 -22878
rect 6463 -22888 6473 -22878
rect 6713 -22878 6793 -22868
rect 6713 -22888 6723 -22878
rect 6463 -22938 6723 -22888
rect 6783 -22938 6793 -22878
rect 6393 -22948 6793 -22938
rect 6851 -22528 7251 -22518
rect 6851 -22588 6861 -22528
rect 6921 -22578 7181 -22528
rect 6921 -22588 6931 -22578
rect 6851 -22598 6931 -22588
rect 7171 -22588 7181 -22578
rect 7241 -22588 7251 -22528
rect 7171 -22598 7251 -22588
rect 6851 -22868 6911 -22598
rect 6991 -22658 7021 -22638
rect 6971 -22698 7021 -22658
rect 7081 -22658 7111 -22638
rect 7081 -22698 7131 -22658
rect 6971 -22768 7131 -22698
rect 6971 -22808 7021 -22768
rect 6991 -22828 7021 -22808
rect 7081 -22808 7131 -22768
rect 7081 -22828 7111 -22808
rect 7191 -22858 7251 -22598
rect 7181 -22868 7251 -22858
rect 6851 -22878 6931 -22868
rect 6851 -22938 6861 -22878
rect 6921 -22888 6931 -22878
rect 7171 -22878 7251 -22868
rect 7171 -22888 7181 -22878
rect 6921 -22938 7181 -22888
rect 7241 -22938 7251 -22878
rect 6851 -22948 7251 -22938
rect 7307 -22528 7707 -22518
rect 7307 -22588 7317 -22528
rect 7377 -22578 7637 -22528
rect 7377 -22588 7387 -22578
rect 7307 -22598 7387 -22588
rect 7627 -22588 7637 -22578
rect 7697 -22588 7707 -22528
rect 7627 -22598 7707 -22588
rect 7307 -22868 7367 -22598
rect 7447 -22658 7477 -22638
rect 7427 -22698 7477 -22658
rect 7537 -22658 7567 -22638
rect 7537 -22698 7587 -22658
rect 7427 -22768 7587 -22698
rect 7427 -22808 7477 -22768
rect 7447 -22828 7477 -22808
rect 7537 -22808 7587 -22768
rect 7537 -22828 7567 -22808
rect 7647 -22858 7707 -22598
rect 7637 -22868 7707 -22858
rect 7307 -22878 7387 -22868
rect 7307 -22938 7317 -22878
rect 7377 -22888 7387 -22878
rect 7627 -22878 7707 -22868
rect 7627 -22888 7637 -22878
rect 7377 -22938 7637 -22888
rect 7697 -22938 7707 -22878
rect 7307 -22948 7707 -22938
rect 7763 -22528 8163 -22518
rect 7763 -22588 7773 -22528
rect 7833 -22578 8093 -22528
rect 7833 -22588 7843 -22578
rect 7763 -22598 7843 -22588
rect 8083 -22588 8093 -22578
rect 8153 -22588 8163 -22528
rect 8083 -22598 8163 -22588
rect 7763 -22868 7823 -22598
rect 7903 -22658 7933 -22638
rect 7883 -22698 7933 -22658
rect 7993 -22658 8023 -22638
rect 7993 -22698 8043 -22658
rect 7883 -22768 8043 -22698
rect 7883 -22808 7933 -22768
rect 7903 -22828 7933 -22808
rect 7993 -22808 8043 -22768
rect 7993 -22828 8023 -22808
rect 8103 -22858 8163 -22598
rect 8093 -22868 8163 -22858
rect 7763 -22878 7843 -22868
rect 7763 -22938 7773 -22878
rect 7833 -22888 7843 -22878
rect 8083 -22878 8163 -22868
rect 8083 -22888 8093 -22878
rect 7833 -22938 8093 -22888
rect 8153 -22938 8163 -22878
rect 7763 -22948 8163 -22938
rect 8237 -22528 8637 -22518
rect 8237 -22588 8247 -22528
rect 8307 -22578 8567 -22528
rect 8307 -22588 8317 -22578
rect 8237 -22598 8317 -22588
rect 8557 -22588 8567 -22578
rect 8627 -22588 8637 -22528
rect 8557 -22598 8637 -22588
rect 8237 -22868 8297 -22598
rect 8377 -22658 8407 -22638
rect 8357 -22698 8407 -22658
rect 8467 -22658 8497 -22638
rect 8467 -22698 8517 -22658
rect 8357 -22768 8517 -22698
rect 8357 -22808 8407 -22768
rect 8377 -22828 8407 -22808
rect 8467 -22808 8517 -22768
rect 8467 -22828 8497 -22808
rect 8577 -22858 8637 -22598
rect 8567 -22868 8637 -22858
rect 8237 -22878 8317 -22868
rect 8237 -22938 8247 -22878
rect 8307 -22888 8317 -22878
rect 8557 -22878 8637 -22868
rect 8557 -22888 8567 -22878
rect 8307 -22938 8567 -22888
rect 8627 -22938 8637 -22878
rect 8237 -22948 8637 -22938
rect 8693 -22528 9093 -22518
rect 8693 -22588 8703 -22528
rect 8763 -22578 9023 -22528
rect 8763 -22588 8773 -22578
rect 8693 -22598 8773 -22588
rect 9013 -22588 9023 -22578
rect 9083 -22588 9093 -22528
rect 9013 -22598 9093 -22588
rect 8693 -22868 8753 -22598
rect 8833 -22658 8863 -22638
rect 8813 -22698 8863 -22658
rect 8923 -22658 8953 -22638
rect 8923 -22698 8973 -22658
rect 8813 -22768 8973 -22698
rect 8813 -22808 8863 -22768
rect 8833 -22828 8863 -22808
rect 8923 -22808 8973 -22768
rect 8923 -22828 8953 -22808
rect 9033 -22858 9093 -22598
rect 9023 -22868 9093 -22858
rect 8693 -22878 8773 -22868
rect 8693 -22938 8703 -22878
rect 8763 -22888 8773 -22878
rect 9013 -22878 9093 -22868
rect 9013 -22888 9023 -22878
rect 8763 -22938 9023 -22888
rect 9083 -22938 9093 -22878
rect 8693 -22948 9093 -22938
rect 9151 -22528 9551 -22518
rect 9151 -22588 9161 -22528
rect 9221 -22578 9481 -22528
rect 9221 -22588 9231 -22578
rect 9151 -22598 9231 -22588
rect 9471 -22588 9481 -22578
rect 9541 -22588 9551 -22528
rect 9471 -22598 9551 -22588
rect 9151 -22868 9211 -22598
rect 9291 -22658 9321 -22638
rect 9271 -22698 9321 -22658
rect 9381 -22658 9411 -22638
rect 9381 -22698 9431 -22658
rect 9271 -22768 9431 -22698
rect 9271 -22808 9321 -22768
rect 9291 -22828 9321 -22808
rect 9381 -22808 9431 -22768
rect 9381 -22828 9411 -22808
rect 9491 -22858 9551 -22598
rect 9481 -22868 9551 -22858
rect 9151 -22878 9231 -22868
rect 9151 -22938 9161 -22878
rect 9221 -22888 9231 -22878
rect 9471 -22878 9551 -22868
rect 9471 -22888 9481 -22878
rect 9221 -22938 9481 -22888
rect 9541 -22938 9551 -22878
rect 9151 -22948 9551 -22938
rect 9607 -22528 10007 -22518
rect 9607 -22588 9617 -22528
rect 9677 -22578 9937 -22528
rect 9677 -22588 9687 -22578
rect 9607 -22598 9687 -22588
rect 9927 -22588 9937 -22578
rect 9997 -22588 10007 -22528
rect 9927 -22598 10007 -22588
rect 9607 -22868 9667 -22598
rect 9747 -22658 9777 -22638
rect 9727 -22698 9777 -22658
rect 9837 -22658 9867 -22638
rect 9837 -22698 9887 -22658
rect 9727 -22768 9887 -22698
rect 9727 -22808 9777 -22768
rect 9747 -22828 9777 -22808
rect 9837 -22808 9887 -22768
rect 9837 -22828 9867 -22808
rect 9947 -22858 10007 -22598
rect 9937 -22868 10007 -22858
rect 9607 -22878 9687 -22868
rect 9607 -22938 9617 -22878
rect 9677 -22888 9687 -22878
rect 9927 -22878 10007 -22868
rect 9927 -22888 9937 -22878
rect 9677 -22938 9937 -22888
rect 9997 -22938 10007 -22878
rect 9607 -22948 10007 -22938
rect 10063 -22528 10463 -22518
rect 10063 -22588 10073 -22528
rect 10133 -22578 10393 -22528
rect 10133 -22588 10143 -22578
rect 10063 -22598 10143 -22588
rect 10383 -22588 10393 -22578
rect 10453 -22588 10463 -22528
rect 10383 -22598 10463 -22588
rect 10063 -22868 10123 -22598
rect 10203 -22658 10233 -22638
rect 10183 -22698 10233 -22658
rect 10293 -22658 10323 -22638
rect 10293 -22698 10343 -22658
rect 10183 -22768 10343 -22698
rect 10183 -22808 10233 -22768
rect 10203 -22828 10233 -22808
rect 10293 -22808 10343 -22768
rect 10293 -22828 10323 -22808
rect 10403 -22858 10463 -22598
rect 10393 -22868 10463 -22858
rect 10063 -22878 10143 -22868
rect 10063 -22938 10073 -22878
rect 10133 -22888 10143 -22878
rect 10383 -22878 10463 -22868
rect 10383 -22888 10393 -22878
rect 10133 -22938 10393 -22888
rect 10453 -22938 10463 -22878
rect 10063 -22948 10463 -22938
rect 10521 -22528 10921 -22518
rect 10521 -22588 10531 -22528
rect 10591 -22578 10851 -22528
rect 10591 -22588 10601 -22578
rect 10521 -22598 10601 -22588
rect 10841 -22588 10851 -22578
rect 10911 -22588 10921 -22528
rect 10841 -22598 10921 -22588
rect 10521 -22868 10581 -22598
rect 10661 -22658 10691 -22638
rect 10641 -22698 10691 -22658
rect 10751 -22658 10781 -22638
rect 10751 -22698 10801 -22658
rect 10641 -22768 10801 -22698
rect 10641 -22808 10691 -22768
rect 10661 -22828 10691 -22808
rect 10751 -22808 10801 -22768
rect 10751 -22828 10781 -22808
rect 10861 -22858 10921 -22598
rect 10851 -22868 10921 -22858
rect 10521 -22878 10601 -22868
rect 10521 -22938 10531 -22878
rect 10591 -22888 10601 -22878
rect 10841 -22878 10921 -22868
rect 10841 -22888 10851 -22878
rect 10591 -22938 10851 -22888
rect 10911 -22938 10921 -22878
rect 10521 -22948 10921 -22938
rect 10977 -22528 11377 -22518
rect 10977 -22588 10987 -22528
rect 11047 -22578 11307 -22528
rect 11047 -22588 11057 -22578
rect 10977 -22598 11057 -22588
rect 11297 -22588 11307 -22578
rect 11367 -22588 11377 -22528
rect 11297 -22598 11377 -22588
rect 10977 -22868 11037 -22598
rect 11117 -22658 11147 -22638
rect 11097 -22698 11147 -22658
rect 11207 -22658 11237 -22638
rect 11207 -22698 11257 -22658
rect 11097 -22768 11257 -22698
rect 11097 -22808 11147 -22768
rect 11117 -22828 11147 -22808
rect 11207 -22808 11257 -22768
rect 11207 -22828 11237 -22808
rect 11317 -22858 11377 -22598
rect 11307 -22868 11377 -22858
rect 10977 -22878 11057 -22868
rect 10977 -22938 10987 -22878
rect 11047 -22888 11057 -22878
rect 11297 -22878 11377 -22868
rect 11297 -22888 11307 -22878
rect 11047 -22938 11307 -22888
rect 11367 -22938 11377 -22878
rect 10977 -22948 11377 -22938
rect 11433 -22528 11833 -22518
rect 11433 -22588 11443 -22528
rect 11503 -22578 11763 -22528
rect 11503 -22588 11513 -22578
rect 11433 -22598 11513 -22588
rect 11753 -22588 11763 -22578
rect 11823 -22588 11833 -22528
rect 11753 -22598 11833 -22588
rect 11433 -22868 11493 -22598
rect 11573 -22658 11603 -22638
rect 11553 -22698 11603 -22658
rect 11663 -22658 11693 -22638
rect 11663 -22698 11713 -22658
rect 11553 -22768 11713 -22698
rect 11553 -22808 11603 -22768
rect 11573 -22828 11603 -22808
rect 11663 -22808 11713 -22768
rect 11663 -22828 11693 -22808
rect 11773 -22858 11833 -22598
rect 11763 -22868 11833 -22858
rect 11433 -22878 11513 -22868
rect 11433 -22938 11443 -22878
rect 11503 -22888 11513 -22878
rect 11753 -22878 11833 -22868
rect 11753 -22888 11763 -22878
rect 11503 -22938 11763 -22888
rect 11823 -22938 11833 -22878
rect 11433 -22948 11833 -22938
rect 11891 -22528 12291 -22518
rect 11891 -22588 11901 -22528
rect 11961 -22578 12221 -22528
rect 11961 -22588 11971 -22578
rect 11891 -22598 11971 -22588
rect 12211 -22588 12221 -22578
rect 12281 -22588 12291 -22528
rect 12211 -22598 12291 -22588
rect 11891 -22868 11951 -22598
rect 12031 -22658 12061 -22638
rect 12011 -22698 12061 -22658
rect 12121 -22658 12151 -22638
rect 12121 -22698 12171 -22658
rect 12011 -22768 12171 -22698
rect 12011 -22808 12061 -22768
rect 12031 -22828 12061 -22808
rect 12121 -22808 12171 -22768
rect 12121 -22828 12151 -22808
rect 12231 -22858 12291 -22598
rect 12221 -22868 12291 -22858
rect 11891 -22878 11971 -22868
rect 11891 -22938 11901 -22878
rect 11961 -22888 11971 -22878
rect 12211 -22878 12291 -22868
rect 12211 -22888 12221 -22878
rect 11961 -22938 12221 -22888
rect 12281 -22938 12291 -22878
rect 11891 -22948 12291 -22938
rect 12347 -22528 12747 -22518
rect 12347 -22588 12357 -22528
rect 12417 -22578 12677 -22528
rect 12417 -22588 12427 -22578
rect 12347 -22598 12427 -22588
rect 12667 -22588 12677 -22578
rect 12737 -22588 12747 -22528
rect 12667 -22598 12747 -22588
rect 12347 -22868 12407 -22598
rect 12487 -22658 12517 -22638
rect 12467 -22698 12517 -22658
rect 12577 -22658 12607 -22638
rect 12577 -22698 12627 -22658
rect 12467 -22768 12627 -22698
rect 12467 -22808 12517 -22768
rect 12487 -22828 12517 -22808
rect 12577 -22808 12627 -22768
rect 12577 -22828 12607 -22808
rect 12687 -22858 12747 -22598
rect 12677 -22868 12747 -22858
rect 12347 -22878 12427 -22868
rect 12347 -22938 12357 -22878
rect 12417 -22888 12427 -22878
rect 12667 -22878 12747 -22868
rect 12667 -22888 12677 -22878
rect 12417 -22938 12677 -22888
rect 12737 -22938 12747 -22878
rect 12347 -22948 12747 -22938
rect 12803 -22528 13203 -22518
rect 12803 -22588 12813 -22528
rect 12873 -22578 13133 -22528
rect 12873 -22588 12883 -22578
rect 12803 -22598 12883 -22588
rect 13123 -22588 13133 -22578
rect 13193 -22588 13203 -22528
rect 13123 -22598 13203 -22588
rect 12803 -22868 12863 -22598
rect 12943 -22658 12973 -22638
rect 12923 -22698 12973 -22658
rect 13033 -22658 13063 -22638
rect 13033 -22698 13083 -22658
rect 12923 -22768 13083 -22698
rect 12923 -22808 12973 -22768
rect 12943 -22828 12973 -22808
rect 13033 -22808 13083 -22768
rect 13033 -22828 13063 -22808
rect 13143 -22858 13203 -22598
rect 13133 -22868 13203 -22858
rect 12803 -22878 12883 -22868
rect 12803 -22938 12813 -22878
rect 12873 -22888 12883 -22878
rect 13123 -22878 13203 -22868
rect 13123 -22888 13133 -22878
rect 12873 -22938 13133 -22888
rect 13193 -22938 13203 -22878
rect 12803 -22948 13203 -22938
rect 13261 -22528 13661 -22518
rect 13261 -22588 13271 -22528
rect 13331 -22578 13591 -22528
rect 13331 -22588 13341 -22578
rect 13261 -22598 13341 -22588
rect 13581 -22588 13591 -22578
rect 13651 -22588 13661 -22528
rect 13581 -22598 13661 -22588
rect 13261 -22868 13321 -22598
rect 13401 -22658 13431 -22638
rect 13381 -22698 13431 -22658
rect 13491 -22658 13521 -22638
rect 13491 -22698 13541 -22658
rect 13381 -22768 13541 -22698
rect 13381 -22808 13431 -22768
rect 13401 -22828 13431 -22808
rect 13491 -22808 13541 -22768
rect 13491 -22828 13521 -22808
rect 13601 -22858 13661 -22598
rect 13591 -22868 13661 -22858
rect 13261 -22878 13341 -22868
rect 13261 -22938 13271 -22878
rect 13331 -22888 13341 -22878
rect 13581 -22878 13661 -22868
rect 13581 -22888 13591 -22878
rect 13331 -22938 13591 -22888
rect 13651 -22938 13661 -22878
rect 13261 -22948 13661 -22938
rect 13717 -22528 14117 -22518
rect 13717 -22588 13727 -22528
rect 13787 -22578 14047 -22528
rect 13787 -22588 13797 -22578
rect 13717 -22598 13797 -22588
rect 14037 -22588 14047 -22578
rect 14107 -22588 14117 -22528
rect 14037 -22598 14117 -22588
rect 13717 -22868 13777 -22598
rect 13857 -22658 13887 -22638
rect 13837 -22698 13887 -22658
rect 13947 -22658 13977 -22638
rect 13947 -22698 13997 -22658
rect 13837 -22768 13997 -22698
rect 13837 -22808 13887 -22768
rect 13857 -22828 13887 -22808
rect 13947 -22808 13997 -22768
rect 13947 -22828 13977 -22808
rect 14057 -22858 14117 -22598
rect 14047 -22868 14117 -22858
rect 13717 -22878 13797 -22868
rect 13717 -22938 13727 -22878
rect 13787 -22888 13797 -22878
rect 14037 -22878 14117 -22868
rect 14037 -22888 14047 -22878
rect 13787 -22938 14047 -22888
rect 14107 -22938 14117 -22878
rect 13717 -22948 14117 -22938
rect 14173 -22528 14573 -22518
rect 14173 -22588 14183 -22528
rect 14243 -22578 14503 -22528
rect 14243 -22588 14253 -22578
rect 14173 -22598 14253 -22588
rect 14493 -22588 14503 -22578
rect 14563 -22588 14573 -22528
rect 14493 -22598 14573 -22588
rect 14173 -22868 14233 -22598
rect 14313 -22658 14343 -22638
rect 14293 -22698 14343 -22658
rect 14403 -22658 14433 -22638
rect 14403 -22698 14453 -22658
rect 14293 -22768 14453 -22698
rect 14293 -22808 14343 -22768
rect 14313 -22828 14343 -22808
rect 14403 -22808 14453 -22768
rect 14403 -22828 14433 -22808
rect 14513 -22858 14573 -22598
rect 14503 -22868 14573 -22858
rect 14173 -22878 14253 -22868
rect 14173 -22938 14183 -22878
rect 14243 -22888 14253 -22878
rect 14493 -22878 14573 -22868
rect 14493 -22888 14503 -22878
rect 14243 -22938 14503 -22888
rect 14563 -22938 14573 -22878
rect 14173 -22948 14573 -22938
rect 14631 -22528 15031 -22518
rect 14631 -22588 14641 -22528
rect 14701 -22578 14961 -22528
rect 14701 -22588 14711 -22578
rect 14631 -22598 14711 -22588
rect 14951 -22588 14961 -22578
rect 15021 -22588 15031 -22528
rect 14951 -22598 15031 -22588
rect 14631 -22868 14691 -22598
rect 14771 -22658 14801 -22638
rect 14751 -22698 14801 -22658
rect 14861 -22658 14891 -22638
rect 14861 -22698 14911 -22658
rect 14751 -22768 14911 -22698
rect 14751 -22808 14801 -22768
rect 14771 -22828 14801 -22808
rect 14861 -22808 14911 -22768
rect 14861 -22828 14891 -22808
rect 14971 -22858 15031 -22598
rect 14961 -22868 15031 -22858
rect 14631 -22878 14711 -22868
rect 14631 -22938 14641 -22878
rect 14701 -22888 14711 -22878
rect 14951 -22878 15031 -22868
rect 14951 -22888 14961 -22878
rect 14701 -22938 14961 -22888
rect 15021 -22938 15031 -22878
rect 14631 -22948 15031 -22938
rect 15087 -22528 15487 -22518
rect 15087 -22588 15097 -22528
rect 15157 -22578 15417 -22528
rect 15157 -22588 15167 -22578
rect 15087 -22598 15167 -22588
rect 15407 -22588 15417 -22578
rect 15477 -22588 15487 -22528
rect 15407 -22598 15487 -22588
rect 15087 -22868 15147 -22598
rect 15227 -22658 15257 -22638
rect 15207 -22698 15257 -22658
rect 15317 -22658 15347 -22638
rect 15317 -22698 15367 -22658
rect 15207 -22768 15367 -22698
rect 15207 -22808 15257 -22768
rect 15227 -22828 15257 -22808
rect 15317 -22808 15367 -22768
rect 15317 -22828 15347 -22808
rect 15427 -22858 15487 -22598
rect 15417 -22868 15487 -22858
rect 15087 -22878 15167 -22868
rect 15087 -22938 15097 -22878
rect 15157 -22888 15167 -22878
rect 15407 -22878 15487 -22868
rect 15407 -22888 15417 -22878
rect 15157 -22938 15417 -22888
rect 15477 -22938 15487 -22878
rect 15087 -22948 15487 -22938
rect 1 -23030 401 -23020
rect 1 -23090 11 -23030
rect 71 -23080 331 -23030
rect 71 -23090 81 -23080
rect 1 -23100 81 -23090
rect 321 -23090 331 -23080
rect 391 -23090 401 -23030
rect 321 -23100 401 -23090
rect 1 -23370 61 -23100
rect 141 -23160 171 -23140
rect 121 -23200 171 -23160
rect 231 -23160 261 -23140
rect 231 -23200 281 -23160
rect 121 -23270 281 -23200
rect 121 -23310 171 -23270
rect 141 -23330 171 -23310
rect 231 -23310 281 -23270
rect 231 -23330 261 -23310
rect 341 -23360 401 -23100
rect 331 -23370 401 -23360
rect 1 -23380 81 -23370
rect 1 -23440 11 -23380
rect 71 -23390 81 -23380
rect 321 -23380 401 -23370
rect 321 -23390 331 -23380
rect 71 -23440 331 -23390
rect 391 -23440 401 -23380
rect 1 -23450 401 -23440
rect 457 -23030 857 -23020
rect 457 -23090 467 -23030
rect 527 -23080 787 -23030
rect 527 -23090 537 -23080
rect 457 -23100 537 -23090
rect 777 -23090 787 -23080
rect 847 -23090 857 -23030
rect 777 -23100 857 -23090
rect 457 -23370 517 -23100
rect 597 -23160 627 -23140
rect 577 -23200 627 -23160
rect 687 -23160 717 -23140
rect 687 -23200 737 -23160
rect 577 -23270 737 -23200
rect 577 -23310 627 -23270
rect 597 -23330 627 -23310
rect 687 -23310 737 -23270
rect 687 -23330 717 -23310
rect 797 -23360 857 -23100
rect 787 -23370 857 -23360
rect 457 -23380 537 -23370
rect 457 -23440 467 -23380
rect 527 -23390 537 -23380
rect 777 -23380 857 -23370
rect 777 -23390 787 -23380
rect 527 -23440 787 -23390
rect 847 -23440 857 -23380
rect 457 -23450 857 -23440
rect 913 -23030 1313 -23020
rect 913 -23090 923 -23030
rect 983 -23080 1243 -23030
rect 983 -23090 993 -23080
rect 913 -23100 993 -23090
rect 1233 -23090 1243 -23080
rect 1303 -23090 1313 -23030
rect 1233 -23100 1313 -23090
rect 913 -23370 973 -23100
rect 1053 -23160 1083 -23140
rect 1033 -23200 1083 -23160
rect 1143 -23160 1173 -23140
rect 1143 -23200 1193 -23160
rect 1033 -23270 1193 -23200
rect 1033 -23310 1083 -23270
rect 1053 -23330 1083 -23310
rect 1143 -23310 1193 -23270
rect 1143 -23330 1173 -23310
rect 1253 -23360 1313 -23100
rect 1243 -23370 1313 -23360
rect 913 -23380 993 -23370
rect 913 -23440 923 -23380
rect 983 -23390 993 -23380
rect 1233 -23380 1313 -23370
rect 1233 -23390 1243 -23380
rect 983 -23440 1243 -23390
rect 1303 -23440 1313 -23380
rect 913 -23450 1313 -23440
rect 1371 -23030 1771 -23020
rect 1371 -23090 1381 -23030
rect 1441 -23080 1701 -23030
rect 1441 -23090 1451 -23080
rect 1371 -23100 1451 -23090
rect 1691 -23090 1701 -23080
rect 1761 -23090 1771 -23030
rect 1691 -23100 1771 -23090
rect 1371 -23370 1431 -23100
rect 1511 -23160 1541 -23140
rect 1491 -23200 1541 -23160
rect 1601 -23160 1631 -23140
rect 1601 -23200 1651 -23160
rect 1491 -23270 1651 -23200
rect 1491 -23310 1541 -23270
rect 1511 -23330 1541 -23310
rect 1601 -23310 1651 -23270
rect 1601 -23330 1631 -23310
rect 1711 -23360 1771 -23100
rect 1701 -23370 1771 -23360
rect 1371 -23380 1451 -23370
rect 1371 -23440 1381 -23380
rect 1441 -23390 1451 -23380
rect 1691 -23380 1771 -23370
rect 1691 -23390 1701 -23380
rect 1441 -23440 1701 -23390
rect 1761 -23440 1771 -23380
rect 1371 -23450 1771 -23440
rect 1827 -23030 2227 -23020
rect 1827 -23090 1837 -23030
rect 1897 -23080 2157 -23030
rect 1897 -23090 1907 -23080
rect 1827 -23100 1907 -23090
rect 2147 -23090 2157 -23080
rect 2217 -23090 2227 -23030
rect 2147 -23100 2227 -23090
rect 1827 -23370 1887 -23100
rect 1967 -23160 1997 -23140
rect 1947 -23200 1997 -23160
rect 2057 -23160 2087 -23140
rect 2057 -23200 2107 -23160
rect 1947 -23270 2107 -23200
rect 1947 -23310 1997 -23270
rect 1967 -23330 1997 -23310
rect 2057 -23310 2107 -23270
rect 2057 -23330 2087 -23310
rect 2167 -23360 2227 -23100
rect 2157 -23370 2227 -23360
rect 1827 -23380 1907 -23370
rect 1827 -23440 1837 -23380
rect 1897 -23390 1907 -23380
rect 2147 -23380 2227 -23370
rect 2147 -23390 2157 -23380
rect 1897 -23440 2157 -23390
rect 2217 -23440 2227 -23380
rect 1827 -23450 2227 -23440
rect 2283 -23030 2683 -23020
rect 2283 -23090 2293 -23030
rect 2353 -23080 2613 -23030
rect 2353 -23090 2363 -23080
rect 2283 -23100 2363 -23090
rect 2603 -23090 2613 -23080
rect 2673 -23090 2683 -23030
rect 2603 -23100 2683 -23090
rect 2283 -23370 2343 -23100
rect 2423 -23160 2453 -23140
rect 2403 -23200 2453 -23160
rect 2513 -23160 2543 -23140
rect 2513 -23200 2563 -23160
rect 2403 -23270 2563 -23200
rect 2403 -23310 2453 -23270
rect 2423 -23330 2453 -23310
rect 2513 -23310 2563 -23270
rect 2513 -23330 2543 -23310
rect 2623 -23360 2683 -23100
rect 2613 -23370 2683 -23360
rect 2283 -23380 2363 -23370
rect 2283 -23440 2293 -23380
rect 2353 -23390 2363 -23380
rect 2603 -23380 2683 -23370
rect 2603 -23390 2613 -23380
rect 2353 -23440 2613 -23390
rect 2673 -23440 2683 -23380
rect 2283 -23450 2683 -23440
rect 2741 -23030 3141 -23020
rect 2741 -23090 2751 -23030
rect 2811 -23080 3071 -23030
rect 2811 -23090 2821 -23080
rect 2741 -23100 2821 -23090
rect 3061 -23090 3071 -23080
rect 3131 -23090 3141 -23030
rect 3061 -23100 3141 -23090
rect 2741 -23370 2801 -23100
rect 2881 -23160 2911 -23140
rect 2861 -23200 2911 -23160
rect 2971 -23160 3001 -23140
rect 2971 -23200 3021 -23160
rect 2861 -23270 3021 -23200
rect 2861 -23310 2911 -23270
rect 2881 -23330 2911 -23310
rect 2971 -23310 3021 -23270
rect 2971 -23330 3001 -23310
rect 3081 -23360 3141 -23100
rect 3071 -23370 3141 -23360
rect 2741 -23380 2821 -23370
rect 2741 -23440 2751 -23380
rect 2811 -23390 2821 -23380
rect 3061 -23380 3141 -23370
rect 3061 -23390 3071 -23380
rect 2811 -23440 3071 -23390
rect 3131 -23440 3141 -23380
rect 2741 -23450 3141 -23440
rect 3197 -23030 3597 -23020
rect 3197 -23090 3207 -23030
rect 3267 -23080 3527 -23030
rect 3267 -23090 3277 -23080
rect 3197 -23100 3277 -23090
rect 3517 -23090 3527 -23080
rect 3587 -23090 3597 -23030
rect 3517 -23100 3597 -23090
rect 3197 -23370 3257 -23100
rect 3337 -23160 3367 -23140
rect 3317 -23200 3367 -23160
rect 3427 -23160 3457 -23140
rect 3427 -23200 3477 -23160
rect 3317 -23270 3477 -23200
rect 3317 -23310 3367 -23270
rect 3337 -23330 3367 -23310
rect 3427 -23310 3477 -23270
rect 3427 -23330 3457 -23310
rect 3537 -23360 3597 -23100
rect 3527 -23370 3597 -23360
rect 3197 -23380 3277 -23370
rect 3197 -23440 3207 -23380
rect 3267 -23390 3277 -23380
rect 3517 -23380 3597 -23370
rect 3517 -23390 3527 -23380
rect 3267 -23440 3527 -23390
rect 3587 -23440 3597 -23380
rect 3197 -23450 3597 -23440
rect 3653 -23030 4053 -23020
rect 3653 -23090 3663 -23030
rect 3723 -23080 3983 -23030
rect 3723 -23090 3733 -23080
rect 3653 -23100 3733 -23090
rect 3973 -23090 3983 -23080
rect 4043 -23090 4053 -23030
rect 3973 -23100 4053 -23090
rect 3653 -23370 3713 -23100
rect 3793 -23160 3823 -23140
rect 3773 -23200 3823 -23160
rect 3883 -23160 3913 -23140
rect 3883 -23200 3933 -23160
rect 3773 -23270 3933 -23200
rect 3773 -23310 3823 -23270
rect 3793 -23330 3823 -23310
rect 3883 -23310 3933 -23270
rect 3883 -23330 3913 -23310
rect 3993 -23360 4053 -23100
rect 3983 -23370 4053 -23360
rect 3653 -23380 3733 -23370
rect 3653 -23440 3663 -23380
rect 3723 -23390 3733 -23380
rect 3973 -23380 4053 -23370
rect 3973 -23390 3983 -23380
rect 3723 -23440 3983 -23390
rect 4043 -23440 4053 -23380
rect 3653 -23450 4053 -23440
rect 4111 -23030 4511 -23020
rect 4111 -23090 4121 -23030
rect 4181 -23080 4441 -23030
rect 4181 -23090 4191 -23080
rect 4111 -23100 4191 -23090
rect 4431 -23090 4441 -23080
rect 4501 -23090 4511 -23030
rect 4431 -23100 4511 -23090
rect 4111 -23370 4171 -23100
rect 4251 -23160 4281 -23140
rect 4231 -23200 4281 -23160
rect 4341 -23160 4371 -23140
rect 4341 -23200 4391 -23160
rect 4231 -23270 4391 -23200
rect 4231 -23310 4281 -23270
rect 4251 -23330 4281 -23310
rect 4341 -23310 4391 -23270
rect 4341 -23330 4371 -23310
rect 4451 -23360 4511 -23100
rect 4441 -23370 4511 -23360
rect 4111 -23380 4191 -23370
rect 4111 -23440 4121 -23380
rect 4181 -23390 4191 -23380
rect 4431 -23380 4511 -23370
rect 4431 -23390 4441 -23380
rect 4181 -23440 4441 -23390
rect 4501 -23440 4511 -23380
rect 4111 -23450 4511 -23440
rect 4567 -23030 4967 -23020
rect 4567 -23090 4577 -23030
rect 4637 -23080 4897 -23030
rect 4637 -23090 4647 -23080
rect 4567 -23100 4647 -23090
rect 4887 -23090 4897 -23080
rect 4957 -23090 4967 -23030
rect 4887 -23100 4967 -23090
rect 4567 -23370 4627 -23100
rect 4707 -23160 4737 -23140
rect 4687 -23200 4737 -23160
rect 4797 -23160 4827 -23140
rect 4797 -23200 4847 -23160
rect 4687 -23270 4847 -23200
rect 4687 -23310 4737 -23270
rect 4707 -23330 4737 -23310
rect 4797 -23310 4847 -23270
rect 4797 -23330 4827 -23310
rect 4907 -23360 4967 -23100
rect 4897 -23370 4967 -23360
rect 4567 -23380 4647 -23370
rect 4567 -23440 4577 -23380
rect 4637 -23390 4647 -23380
rect 4887 -23380 4967 -23370
rect 4887 -23390 4897 -23380
rect 4637 -23440 4897 -23390
rect 4957 -23440 4967 -23380
rect 4567 -23450 4967 -23440
rect 5023 -23030 5423 -23020
rect 5023 -23090 5033 -23030
rect 5093 -23080 5353 -23030
rect 5093 -23090 5103 -23080
rect 5023 -23100 5103 -23090
rect 5343 -23090 5353 -23080
rect 5413 -23090 5423 -23030
rect 5343 -23100 5423 -23090
rect 5023 -23370 5083 -23100
rect 5163 -23160 5193 -23140
rect 5143 -23200 5193 -23160
rect 5253 -23160 5283 -23140
rect 5253 -23200 5303 -23160
rect 5143 -23270 5303 -23200
rect 5143 -23310 5193 -23270
rect 5163 -23330 5193 -23310
rect 5253 -23310 5303 -23270
rect 5253 -23330 5283 -23310
rect 5363 -23360 5423 -23100
rect 5353 -23370 5423 -23360
rect 5023 -23380 5103 -23370
rect 5023 -23440 5033 -23380
rect 5093 -23390 5103 -23380
rect 5343 -23380 5423 -23370
rect 5343 -23390 5353 -23380
rect 5093 -23440 5353 -23390
rect 5413 -23440 5423 -23380
rect 5023 -23450 5423 -23440
rect 5481 -23030 5881 -23020
rect 5481 -23090 5491 -23030
rect 5551 -23080 5811 -23030
rect 5551 -23090 5561 -23080
rect 5481 -23100 5561 -23090
rect 5801 -23090 5811 -23080
rect 5871 -23090 5881 -23030
rect 5801 -23100 5881 -23090
rect 5481 -23370 5541 -23100
rect 5621 -23160 5651 -23140
rect 5601 -23200 5651 -23160
rect 5711 -23160 5741 -23140
rect 5711 -23200 5761 -23160
rect 5601 -23270 5761 -23200
rect 5601 -23310 5651 -23270
rect 5621 -23330 5651 -23310
rect 5711 -23310 5761 -23270
rect 5711 -23330 5741 -23310
rect 5821 -23360 5881 -23100
rect 5811 -23370 5881 -23360
rect 5481 -23380 5561 -23370
rect 5481 -23440 5491 -23380
rect 5551 -23390 5561 -23380
rect 5801 -23380 5881 -23370
rect 5801 -23390 5811 -23380
rect 5551 -23440 5811 -23390
rect 5871 -23440 5881 -23380
rect 5481 -23450 5881 -23440
rect 5937 -23030 6337 -23020
rect 5937 -23090 5947 -23030
rect 6007 -23080 6267 -23030
rect 6007 -23090 6017 -23080
rect 5937 -23100 6017 -23090
rect 6257 -23090 6267 -23080
rect 6327 -23090 6337 -23030
rect 6257 -23100 6337 -23090
rect 5937 -23370 5997 -23100
rect 6077 -23160 6107 -23140
rect 6057 -23200 6107 -23160
rect 6167 -23160 6197 -23140
rect 6167 -23200 6217 -23160
rect 6057 -23270 6217 -23200
rect 6057 -23310 6107 -23270
rect 6077 -23330 6107 -23310
rect 6167 -23310 6217 -23270
rect 6167 -23330 6197 -23310
rect 6277 -23360 6337 -23100
rect 6267 -23370 6337 -23360
rect 5937 -23380 6017 -23370
rect 5937 -23440 5947 -23380
rect 6007 -23390 6017 -23380
rect 6257 -23380 6337 -23370
rect 6257 -23390 6267 -23380
rect 6007 -23440 6267 -23390
rect 6327 -23440 6337 -23380
rect 5937 -23450 6337 -23440
rect 6393 -23030 6793 -23020
rect 6393 -23090 6403 -23030
rect 6463 -23080 6723 -23030
rect 6463 -23090 6473 -23080
rect 6393 -23100 6473 -23090
rect 6713 -23090 6723 -23080
rect 6783 -23090 6793 -23030
rect 6713 -23100 6793 -23090
rect 6393 -23370 6453 -23100
rect 6533 -23160 6563 -23140
rect 6513 -23200 6563 -23160
rect 6623 -23160 6653 -23140
rect 6623 -23200 6673 -23160
rect 6513 -23270 6673 -23200
rect 6513 -23310 6563 -23270
rect 6533 -23330 6563 -23310
rect 6623 -23310 6673 -23270
rect 6623 -23330 6653 -23310
rect 6733 -23360 6793 -23100
rect 6723 -23370 6793 -23360
rect 6393 -23380 6473 -23370
rect 6393 -23440 6403 -23380
rect 6463 -23390 6473 -23380
rect 6713 -23380 6793 -23370
rect 6713 -23390 6723 -23380
rect 6463 -23440 6723 -23390
rect 6783 -23440 6793 -23380
rect 6393 -23450 6793 -23440
rect 6851 -23030 7251 -23020
rect 6851 -23090 6861 -23030
rect 6921 -23080 7181 -23030
rect 6921 -23090 6931 -23080
rect 6851 -23100 6931 -23090
rect 7171 -23090 7181 -23080
rect 7241 -23090 7251 -23030
rect 7171 -23100 7251 -23090
rect 6851 -23370 6911 -23100
rect 6991 -23160 7021 -23140
rect 6971 -23200 7021 -23160
rect 7081 -23160 7111 -23140
rect 7081 -23200 7131 -23160
rect 6971 -23270 7131 -23200
rect 6971 -23310 7021 -23270
rect 6991 -23330 7021 -23310
rect 7081 -23310 7131 -23270
rect 7081 -23330 7111 -23310
rect 7191 -23360 7251 -23100
rect 7181 -23370 7251 -23360
rect 6851 -23380 6931 -23370
rect 6851 -23440 6861 -23380
rect 6921 -23390 6931 -23380
rect 7171 -23380 7251 -23370
rect 7171 -23390 7181 -23380
rect 6921 -23440 7181 -23390
rect 7241 -23440 7251 -23380
rect 6851 -23450 7251 -23440
rect 7307 -23030 7707 -23020
rect 7307 -23090 7317 -23030
rect 7377 -23080 7637 -23030
rect 7377 -23090 7387 -23080
rect 7307 -23100 7387 -23090
rect 7627 -23090 7637 -23080
rect 7697 -23090 7707 -23030
rect 7627 -23100 7707 -23090
rect 7307 -23370 7367 -23100
rect 7447 -23160 7477 -23140
rect 7427 -23200 7477 -23160
rect 7537 -23160 7567 -23140
rect 7537 -23200 7587 -23160
rect 7427 -23270 7587 -23200
rect 7427 -23310 7477 -23270
rect 7447 -23330 7477 -23310
rect 7537 -23310 7587 -23270
rect 7537 -23330 7567 -23310
rect 7647 -23360 7707 -23100
rect 7637 -23370 7707 -23360
rect 7307 -23380 7387 -23370
rect 7307 -23440 7317 -23380
rect 7377 -23390 7387 -23380
rect 7627 -23380 7707 -23370
rect 7627 -23390 7637 -23380
rect 7377 -23440 7637 -23390
rect 7697 -23440 7707 -23380
rect 7307 -23450 7707 -23440
rect 7763 -23030 8163 -23020
rect 7763 -23090 7773 -23030
rect 7833 -23080 8093 -23030
rect 7833 -23090 7843 -23080
rect 7763 -23100 7843 -23090
rect 8083 -23090 8093 -23080
rect 8153 -23090 8163 -23030
rect 8083 -23100 8163 -23090
rect 7763 -23370 7823 -23100
rect 7903 -23160 7933 -23140
rect 7883 -23200 7933 -23160
rect 7993 -23160 8023 -23140
rect 7993 -23200 8043 -23160
rect 7883 -23270 8043 -23200
rect 7883 -23310 7933 -23270
rect 7903 -23330 7933 -23310
rect 7993 -23310 8043 -23270
rect 7993 -23330 8023 -23310
rect 8103 -23360 8163 -23100
rect 8093 -23370 8163 -23360
rect 7763 -23380 7843 -23370
rect 7763 -23440 7773 -23380
rect 7833 -23390 7843 -23380
rect 8083 -23380 8163 -23370
rect 8083 -23390 8093 -23380
rect 7833 -23440 8093 -23390
rect 8153 -23440 8163 -23380
rect 7763 -23450 8163 -23440
rect 8237 -23030 8637 -23020
rect 8237 -23090 8247 -23030
rect 8307 -23080 8567 -23030
rect 8307 -23090 8317 -23080
rect 8237 -23100 8317 -23090
rect 8557 -23090 8567 -23080
rect 8627 -23090 8637 -23030
rect 8557 -23100 8637 -23090
rect 8237 -23370 8297 -23100
rect 8377 -23160 8407 -23140
rect 8357 -23200 8407 -23160
rect 8467 -23160 8497 -23140
rect 8467 -23200 8517 -23160
rect 8357 -23270 8517 -23200
rect 8357 -23310 8407 -23270
rect 8377 -23330 8407 -23310
rect 8467 -23310 8517 -23270
rect 8467 -23330 8497 -23310
rect 8577 -23360 8637 -23100
rect 8567 -23370 8637 -23360
rect 8237 -23380 8317 -23370
rect 8237 -23440 8247 -23380
rect 8307 -23390 8317 -23380
rect 8557 -23380 8637 -23370
rect 8557 -23390 8567 -23380
rect 8307 -23440 8567 -23390
rect 8627 -23440 8637 -23380
rect 8237 -23450 8637 -23440
rect 8693 -23030 9093 -23020
rect 8693 -23090 8703 -23030
rect 8763 -23080 9023 -23030
rect 8763 -23090 8773 -23080
rect 8693 -23100 8773 -23090
rect 9013 -23090 9023 -23080
rect 9083 -23090 9093 -23030
rect 9013 -23100 9093 -23090
rect 8693 -23370 8753 -23100
rect 8833 -23160 8863 -23140
rect 8813 -23200 8863 -23160
rect 8923 -23160 8953 -23140
rect 8923 -23200 8973 -23160
rect 8813 -23270 8973 -23200
rect 8813 -23310 8863 -23270
rect 8833 -23330 8863 -23310
rect 8923 -23310 8973 -23270
rect 8923 -23330 8953 -23310
rect 9033 -23360 9093 -23100
rect 9023 -23370 9093 -23360
rect 8693 -23380 8773 -23370
rect 8693 -23440 8703 -23380
rect 8763 -23390 8773 -23380
rect 9013 -23380 9093 -23370
rect 9013 -23390 9023 -23380
rect 8763 -23440 9023 -23390
rect 9083 -23440 9093 -23380
rect 8693 -23450 9093 -23440
rect 9151 -23030 9551 -23020
rect 9151 -23090 9161 -23030
rect 9221 -23080 9481 -23030
rect 9221 -23090 9231 -23080
rect 9151 -23100 9231 -23090
rect 9471 -23090 9481 -23080
rect 9541 -23090 9551 -23030
rect 9471 -23100 9551 -23090
rect 9151 -23370 9211 -23100
rect 9291 -23160 9321 -23140
rect 9271 -23200 9321 -23160
rect 9381 -23160 9411 -23140
rect 9381 -23200 9431 -23160
rect 9271 -23270 9431 -23200
rect 9271 -23310 9321 -23270
rect 9291 -23330 9321 -23310
rect 9381 -23310 9431 -23270
rect 9381 -23330 9411 -23310
rect 9491 -23360 9551 -23100
rect 9481 -23370 9551 -23360
rect 9151 -23380 9231 -23370
rect 9151 -23440 9161 -23380
rect 9221 -23390 9231 -23380
rect 9471 -23380 9551 -23370
rect 9471 -23390 9481 -23380
rect 9221 -23440 9481 -23390
rect 9541 -23440 9551 -23380
rect 9151 -23450 9551 -23440
rect 9607 -23030 10007 -23020
rect 9607 -23090 9617 -23030
rect 9677 -23080 9937 -23030
rect 9677 -23090 9687 -23080
rect 9607 -23100 9687 -23090
rect 9927 -23090 9937 -23080
rect 9997 -23090 10007 -23030
rect 9927 -23100 10007 -23090
rect 9607 -23370 9667 -23100
rect 9747 -23160 9777 -23140
rect 9727 -23200 9777 -23160
rect 9837 -23160 9867 -23140
rect 9837 -23200 9887 -23160
rect 9727 -23270 9887 -23200
rect 9727 -23310 9777 -23270
rect 9747 -23330 9777 -23310
rect 9837 -23310 9887 -23270
rect 9837 -23330 9867 -23310
rect 9947 -23360 10007 -23100
rect 9937 -23370 10007 -23360
rect 9607 -23380 9687 -23370
rect 9607 -23440 9617 -23380
rect 9677 -23390 9687 -23380
rect 9927 -23380 10007 -23370
rect 9927 -23390 9937 -23380
rect 9677 -23440 9937 -23390
rect 9997 -23440 10007 -23380
rect 9607 -23450 10007 -23440
rect 10063 -23030 10463 -23020
rect 10063 -23090 10073 -23030
rect 10133 -23080 10393 -23030
rect 10133 -23090 10143 -23080
rect 10063 -23100 10143 -23090
rect 10383 -23090 10393 -23080
rect 10453 -23090 10463 -23030
rect 10383 -23100 10463 -23090
rect 10063 -23370 10123 -23100
rect 10203 -23160 10233 -23140
rect 10183 -23200 10233 -23160
rect 10293 -23160 10323 -23140
rect 10293 -23200 10343 -23160
rect 10183 -23270 10343 -23200
rect 10183 -23310 10233 -23270
rect 10203 -23330 10233 -23310
rect 10293 -23310 10343 -23270
rect 10293 -23330 10323 -23310
rect 10403 -23360 10463 -23100
rect 10393 -23370 10463 -23360
rect 10063 -23380 10143 -23370
rect 10063 -23440 10073 -23380
rect 10133 -23390 10143 -23380
rect 10383 -23380 10463 -23370
rect 10383 -23390 10393 -23380
rect 10133 -23440 10393 -23390
rect 10453 -23440 10463 -23380
rect 10063 -23450 10463 -23440
rect 10521 -23030 10921 -23020
rect 10521 -23090 10531 -23030
rect 10591 -23080 10851 -23030
rect 10591 -23090 10601 -23080
rect 10521 -23100 10601 -23090
rect 10841 -23090 10851 -23080
rect 10911 -23090 10921 -23030
rect 10841 -23100 10921 -23090
rect 10521 -23370 10581 -23100
rect 10661 -23160 10691 -23140
rect 10641 -23200 10691 -23160
rect 10751 -23160 10781 -23140
rect 10751 -23200 10801 -23160
rect 10641 -23270 10801 -23200
rect 10641 -23310 10691 -23270
rect 10661 -23330 10691 -23310
rect 10751 -23310 10801 -23270
rect 10751 -23330 10781 -23310
rect 10861 -23360 10921 -23100
rect 10851 -23370 10921 -23360
rect 10521 -23380 10601 -23370
rect 10521 -23440 10531 -23380
rect 10591 -23390 10601 -23380
rect 10841 -23380 10921 -23370
rect 10841 -23390 10851 -23380
rect 10591 -23440 10851 -23390
rect 10911 -23440 10921 -23380
rect 10521 -23450 10921 -23440
rect 10977 -23030 11377 -23020
rect 10977 -23090 10987 -23030
rect 11047 -23080 11307 -23030
rect 11047 -23090 11057 -23080
rect 10977 -23100 11057 -23090
rect 11297 -23090 11307 -23080
rect 11367 -23090 11377 -23030
rect 11297 -23100 11377 -23090
rect 10977 -23370 11037 -23100
rect 11117 -23160 11147 -23140
rect 11097 -23200 11147 -23160
rect 11207 -23160 11237 -23140
rect 11207 -23200 11257 -23160
rect 11097 -23270 11257 -23200
rect 11097 -23310 11147 -23270
rect 11117 -23330 11147 -23310
rect 11207 -23310 11257 -23270
rect 11207 -23330 11237 -23310
rect 11317 -23360 11377 -23100
rect 11307 -23370 11377 -23360
rect 10977 -23380 11057 -23370
rect 10977 -23440 10987 -23380
rect 11047 -23390 11057 -23380
rect 11297 -23380 11377 -23370
rect 11297 -23390 11307 -23380
rect 11047 -23440 11307 -23390
rect 11367 -23440 11377 -23380
rect 10977 -23450 11377 -23440
rect 11433 -23030 11833 -23020
rect 11433 -23090 11443 -23030
rect 11503 -23080 11763 -23030
rect 11503 -23090 11513 -23080
rect 11433 -23100 11513 -23090
rect 11753 -23090 11763 -23080
rect 11823 -23090 11833 -23030
rect 11753 -23100 11833 -23090
rect 11433 -23370 11493 -23100
rect 11573 -23160 11603 -23140
rect 11553 -23200 11603 -23160
rect 11663 -23160 11693 -23140
rect 11663 -23200 11713 -23160
rect 11553 -23270 11713 -23200
rect 11553 -23310 11603 -23270
rect 11573 -23330 11603 -23310
rect 11663 -23310 11713 -23270
rect 11663 -23330 11693 -23310
rect 11773 -23360 11833 -23100
rect 11763 -23370 11833 -23360
rect 11433 -23380 11513 -23370
rect 11433 -23440 11443 -23380
rect 11503 -23390 11513 -23380
rect 11753 -23380 11833 -23370
rect 11753 -23390 11763 -23380
rect 11503 -23440 11763 -23390
rect 11823 -23440 11833 -23380
rect 11433 -23450 11833 -23440
rect 11891 -23030 12291 -23020
rect 11891 -23090 11901 -23030
rect 11961 -23080 12221 -23030
rect 11961 -23090 11971 -23080
rect 11891 -23100 11971 -23090
rect 12211 -23090 12221 -23080
rect 12281 -23090 12291 -23030
rect 12211 -23100 12291 -23090
rect 11891 -23370 11951 -23100
rect 12031 -23160 12061 -23140
rect 12011 -23200 12061 -23160
rect 12121 -23160 12151 -23140
rect 12121 -23200 12171 -23160
rect 12011 -23270 12171 -23200
rect 12011 -23310 12061 -23270
rect 12031 -23330 12061 -23310
rect 12121 -23310 12171 -23270
rect 12121 -23330 12151 -23310
rect 12231 -23360 12291 -23100
rect 12221 -23370 12291 -23360
rect 11891 -23380 11971 -23370
rect 11891 -23440 11901 -23380
rect 11961 -23390 11971 -23380
rect 12211 -23380 12291 -23370
rect 12211 -23390 12221 -23380
rect 11961 -23440 12221 -23390
rect 12281 -23440 12291 -23380
rect 11891 -23450 12291 -23440
rect 12347 -23030 12747 -23020
rect 12347 -23090 12357 -23030
rect 12417 -23080 12677 -23030
rect 12417 -23090 12427 -23080
rect 12347 -23100 12427 -23090
rect 12667 -23090 12677 -23080
rect 12737 -23090 12747 -23030
rect 12667 -23100 12747 -23090
rect 12347 -23370 12407 -23100
rect 12487 -23160 12517 -23140
rect 12467 -23200 12517 -23160
rect 12577 -23160 12607 -23140
rect 12577 -23200 12627 -23160
rect 12467 -23270 12627 -23200
rect 12467 -23310 12517 -23270
rect 12487 -23330 12517 -23310
rect 12577 -23310 12627 -23270
rect 12577 -23330 12607 -23310
rect 12687 -23360 12747 -23100
rect 12677 -23370 12747 -23360
rect 12347 -23380 12427 -23370
rect 12347 -23440 12357 -23380
rect 12417 -23390 12427 -23380
rect 12667 -23380 12747 -23370
rect 12667 -23390 12677 -23380
rect 12417 -23440 12677 -23390
rect 12737 -23440 12747 -23380
rect 12347 -23450 12747 -23440
rect 12803 -23030 13203 -23020
rect 12803 -23090 12813 -23030
rect 12873 -23080 13133 -23030
rect 12873 -23090 12883 -23080
rect 12803 -23100 12883 -23090
rect 13123 -23090 13133 -23080
rect 13193 -23090 13203 -23030
rect 13123 -23100 13203 -23090
rect 12803 -23370 12863 -23100
rect 12943 -23160 12973 -23140
rect 12923 -23200 12973 -23160
rect 13033 -23160 13063 -23140
rect 13033 -23200 13083 -23160
rect 12923 -23270 13083 -23200
rect 12923 -23310 12973 -23270
rect 12943 -23330 12973 -23310
rect 13033 -23310 13083 -23270
rect 13033 -23330 13063 -23310
rect 13143 -23360 13203 -23100
rect 13133 -23370 13203 -23360
rect 12803 -23380 12883 -23370
rect 12803 -23440 12813 -23380
rect 12873 -23390 12883 -23380
rect 13123 -23380 13203 -23370
rect 13123 -23390 13133 -23380
rect 12873 -23440 13133 -23390
rect 13193 -23440 13203 -23380
rect 12803 -23450 13203 -23440
rect 13261 -23030 13661 -23020
rect 13261 -23090 13271 -23030
rect 13331 -23080 13591 -23030
rect 13331 -23090 13341 -23080
rect 13261 -23100 13341 -23090
rect 13581 -23090 13591 -23080
rect 13651 -23090 13661 -23030
rect 13581 -23100 13661 -23090
rect 13261 -23370 13321 -23100
rect 13401 -23160 13431 -23140
rect 13381 -23200 13431 -23160
rect 13491 -23160 13521 -23140
rect 13491 -23200 13541 -23160
rect 13381 -23270 13541 -23200
rect 13381 -23310 13431 -23270
rect 13401 -23330 13431 -23310
rect 13491 -23310 13541 -23270
rect 13491 -23330 13521 -23310
rect 13601 -23360 13661 -23100
rect 13591 -23370 13661 -23360
rect 13261 -23380 13341 -23370
rect 13261 -23440 13271 -23380
rect 13331 -23390 13341 -23380
rect 13581 -23380 13661 -23370
rect 13581 -23390 13591 -23380
rect 13331 -23440 13591 -23390
rect 13651 -23440 13661 -23380
rect 13261 -23450 13661 -23440
rect 13717 -23030 14117 -23020
rect 13717 -23090 13727 -23030
rect 13787 -23080 14047 -23030
rect 13787 -23090 13797 -23080
rect 13717 -23100 13797 -23090
rect 14037 -23090 14047 -23080
rect 14107 -23090 14117 -23030
rect 14037 -23100 14117 -23090
rect 13717 -23370 13777 -23100
rect 13857 -23160 13887 -23140
rect 13837 -23200 13887 -23160
rect 13947 -23160 13977 -23140
rect 13947 -23200 13997 -23160
rect 13837 -23270 13997 -23200
rect 13837 -23310 13887 -23270
rect 13857 -23330 13887 -23310
rect 13947 -23310 13997 -23270
rect 13947 -23330 13977 -23310
rect 14057 -23360 14117 -23100
rect 14047 -23370 14117 -23360
rect 13717 -23380 13797 -23370
rect 13717 -23440 13727 -23380
rect 13787 -23390 13797 -23380
rect 14037 -23380 14117 -23370
rect 14037 -23390 14047 -23380
rect 13787 -23440 14047 -23390
rect 14107 -23440 14117 -23380
rect 13717 -23450 14117 -23440
rect 14173 -23030 14573 -23020
rect 14173 -23090 14183 -23030
rect 14243 -23080 14503 -23030
rect 14243 -23090 14253 -23080
rect 14173 -23100 14253 -23090
rect 14493 -23090 14503 -23080
rect 14563 -23090 14573 -23030
rect 14493 -23100 14573 -23090
rect 14173 -23370 14233 -23100
rect 14313 -23160 14343 -23140
rect 14293 -23200 14343 -23160
rect 14403 -23160 14433 -23140
rect 14403 -23200 14453 -23160
rect 14293 -23270 14453 -23200
rect 14293 -23310 14343 -23270
rect 14313 -23330 14343 -23310
rect 14403 -23310 14453 -23270
rect 14403 -23330 14433 -23310
rect 14513 -23360 14573 -23100
rect 14503 -23370 14573 -23360
rect 14173 -23380 14253 -23370
rect 14173 -23440 14183 -23380
rect 14243 -23390 14253 -23380
rect 14493 -23380 14573 -23370
rect 14493 -23390 14503 -23380
rect 14243 -23440 14503 -23390
rect 14563 -23440 14573 -23380
rect 14173 -23450 14573 -23440
rect 14631 -23030 15031 -23020
rect 14631 -23090 14641 -23030
rect 14701 -23080 14961 -23030
rect 14701 -23090 14711 -23080
rect 14631 -23100 14711 -23090
rect 14951 -23090 14961 -23080
rect 15021 -23090 15031 -23030
rect 14951 -23100 15031 -23090
rect 14631 -23370 14691 -23100
rect 14771 -23160 14801 -23140
rect 14751 -23200 14801 -23160
rect 14861 -23160 14891 -23140
rect 14861 -23200 14911 -23160
rect 14751 -23270 14911 -23200
rect 14751 -23310 14801 -23270
rect 14771 -23330 14801 -23310
rect 14861 -23310 14911 -23270
rect 14861 -23330 14891 -23310
rect 14971 -23360 15031 -23100
rect 14961 -23370 15031 -23360
rect 14631 -23380 14711 -23370
rect 14631 -23440 14641 -23380
rect 14701 -23390 14711 -23380
rect 14951 -23380 15031 -23370
rect 14951 -23390 14961 -23380
rect 14701 -23440 14961 -23390
rect 15021 -23440 15031 -23380
rect 14631 -23450 15031 -23440
rect 15087 -23030 15487 -23020
rect 15087 -23090 15097 -23030
rect 15157 -23080 15417 -23030
rect 15157 -23090 15167 -23080
rect 15087 -23100 15167 -23090
rect 15407 -23090 15417 -23080
rect 15477 -23090 15487 -23030
rect 15407 -23100 15487 -23090
rect 15087 -23370 15147 -23100
rect 15227 -23160 15257 -23140
rect 15207 -23200 15257 -23160
rect 15317 -23160 15347 -23140
rect 15317 -23200 15367 -23160
rect 15207 -23270 15367 -23200
rect 15207 -23310 15257 -23270
rect 15227 -23330 15257 -23310
rect 15317 -23310 15367 -23270
rect 15317 -23330 15347 -23310
rect 15427 -23360 15487 -23100
rect 15417 -23370 15487 -23360
rect 15087 -23380 15167 -23370
rect 15087 -23440 15097 -23380
rect 15157 -23390 15167 -23380
rect 15407 -23380 15487 -23370
rect 15407 -23390 15417 -23380
rect 15157 -23440 15417 -23390
rect 15477 -23440 15487 -23380
rect 15087 -23450 15487 -23440
rect 1 -23524 401 -23514
rect 1 -23584 11 -23524
rect 71 -23574 331 -23524
rect 71 -23584 81 -23574
rect 1 -23594 81 -23584
rect 321 -23584 331 -23574
rect 391 -23584 401 -23524
rect 321 -23594 401 -23584
rect 1 -23864 61 -23594
rect 141 -23654 171 -23634
rect 121 -23694 171 -23654
rect 231 -23654 261 -23634
rect 231 -23694 281 -23654
rect 121 -23764 281 -23694
rect 121 -23804 171 -23764
rect 141 -23824 171 -23804
rect 231 -23804 281 -23764
rect 231 -23824 261 -23804
rect 341 -23854 401 -23594
rect 331 -23864 401 -23854
rect 1 -23874 81 -23864
rect 1 -23934 11 -23874
rect 71 -23884 81 -23874
rect 321 -23874 401 -23864
rect 321 -23884 331 -23874
rect 71 -23934 331 -23884
rect 391 -23934 401 -23874
rect 1 -23944 401 -23934
rect 457 -23524 857 -23514
rect 457 -23584 467 -23524
rect 527 -23574 787 -23524
rect 527 -23584 537 -23574
rect 457 -23594 537 -23584
rect 777 -23584 787 -23574
rect 847 -23584 857 -23524
rect 777 -23594 857 -23584
rect 457 -23864 517 -23594
rect 597 -23654 627 -23634
rect 577 -23694 627 -23654
rect 687 -23654 717 -23634
rect 687 -23694 737 -23654
rect 577 -23764 737 -23694
rect 577 -23804 627 -23764
rect 597 -23824 627 -23804
rect 687 -23804 737 -23764
rect 687 -23824 717 -23804
rect 797 -23854 857 -23594
rect 787 -23864 857 -23854
rect 457 -23874 537 -23864
rect 457 -23934 467 -23874
rect 527 -23884 537 -23874
rect 777 -23874 857 -23864
rect 777 -23884 787 -23874
rect 527 -23934 787 -23884
rect 847 -23934 857 -23874
rect 457 -23944 857 -23934
rect 913 -23524 1313 -23514
rect 913 -23584 923 -23524
rect 983 -23574 1243 -23524
rect 983 -23584 993 -23574
rect 913 -23594 993 -23584
rect 1233 -23584 1243 -23574
rect 1303 -23584 1313 -23524
rect 1233 -23594 1313 -23584
rect 913 -23864 973 -23594
rect 1053 -23654 1083 -23634
rect 1033 -23694 1083 -23654
rect 1143 -23654 1173 -23634
rect 1143 -23694 1193 -23654
rect 1033 -23764 1193 -23694
rect 1033 -23804 1083 -23764
rect 1053 -23824 1083 -23804
rect 1143 -23804 1193 -23764
rect 1143 -23824 1173 -23804
rect 1253 -23854 1313 -23594
rect 1243 -23864 1313 -23854
rect 913 -23874 993 -23864
rect 913 -23934 923 -23874
rect 983 -23884 993 -23874
rect 1233 -23874 1313 -23864
rect 1233 -23884 1243 -23874
rect 983 -23934 1243 -23884
rect 1303 -23934 1313 -23874
rect 913 -23944 1313 -23934
rect 1371 -23524 1771 -23514
rect 1371 -23584 1381 -23524
rect 1441 -23574 1701 -23524
rect 1441 -23584 1451 -23574
rect 1371 -23594 1451 -23584
rect 1691 -23584 1701 -23574
rect 1761 -23584 1771 -23524
rect 1691 -23594 1771 -23584
rect 1371 -23864 1431 -23594
rect 1511 -23654 1541 -23634
rect 1491 -23694 1541 -23654
rect 1601 -23654 1631 -23634
rect 1601 -23694 1651 -23654
rect 1491 -23764 1651 -23694
rect 1491 -23804 1541 -23764
rect 1511 -23824 1541 -23804
rect 1601 -23804 1651 -23764
rect 1601 -23824 1631 -23804
rect 1711 -23854 1771 -23594
rect 1701 -23864 1771 -23854
rect 1371 -23874 1451 -23864
rect 1371 -23934 1381 -23874
rect 1441 -23884 1451 -23874
rect 1691 -23874 1771 -23864
rect 1691 -23884 1701 -23874
rect 1441 -23934 1701 -23884
rect 1761 -23934 1771 -23874
rect 1371 -23944 1771 -23934
rect 1827 -23524 2227 -23514
rect 1827 -23584 1837 -23524
rect 1897 -23574 2157 -23524
rect 1897 -23584 1907 -23574
rect 1827 -23594 1907 -23584
rect 2147 -23584 2157 -23574
rect 2217 -23584 2227 -23524
rect 2147 -23594 2227 -23584
rect 1827 -23864 1887 -23594
rect 1967 -23654 1997 -23634
rect 1947 -23694 1997 -23654
rect 2057 -23654 2087 -23634
rect 2057 -23694 2107 -23654
rect 1947 -23764 2107 -23694
rect 1947 -23804 1997 -23764
rect 1967 -23824 1997 -23804
rect 2057 -23804 2107 -23764
rect 2057 -23824 2087 -23804
rect 2167 -23854 2227 -23594
rect 2157 -23864 2227 -23854
rect 1827 -23874 1907 -23864
rect 1827 -23934 1837 -23874
rect 1897 -23884 1907 -23874
rect 2147 -23874 2227 -23864
rect 2147 -23884 2157 -23874
rect 1897 -23934 2157 -23884
rect 2217 -23934 2227 -23874
rect 1827 -23944 2227 -23934
rect 2283 -23524 2683 -23514
rect 2283 -23584 2293 -23524
rect 2353 -23574 2613 -23524
rect 2353 -23584 2363 -23574
rect 2283 -23594 2363 -23584
rect 2603 -23584 2613 -23574
rect 2673 -23584 2683 -23524
rect 2603 -23594 2683 -23584
rect 2283 -23864 2343 -23594
rect 2423 -23654 2453 -23634
rect 2403 -23694 2453 -23654
rect 2513 -23654 2543 -23634
rect 2513 -23694 2563 -23654
rect 2403 -23764 2563 -23694
rect 2403 -23804 2453 -23764
rect 2423 -23824 2453 -23804
rect 2513 -23804 2563 -23764
rect 2513 -23824 2543 -23804
rect 2623 -23854 2683 -23594
rect 2613 -23864 2683 -23854
rect 2283 -23874 2363 -23864
rect 2283 -23934 2293 -23874
rect 2353 -23884 2363 -23874
rect 2603 -23874 2683 -23864
rect 2603 -23884 2613 -23874
rect 2353 -23934 2613 -23884
rect 2673 -23934 2683 -23874
rect 2283 -23944 2683 -23934
rect 2741 -23524 3141 -23514
rect 2741 -23584 2751 -23524
rect 2811 -23574 3071 -23524
rect 2811 -23584 2821 -23574
rect 2741 -23594 2821 -23584
rect 3061 -23584 3071 -23574
rect 3131 -23584 3141 -23524
rect 3061 -23594 3141 -23584
rect 2741 -23864 2801 -23594
rect 2881 -23654 2911 -23634
rect 2861 -23694 2911 -23654
rect 2971 -23654 3001 -23634
rect 2971 -23694 3021 -23654
rect 2861 -23764 3021 -23694
rect 2861 -23804 2911 -23764
rect 2881 -23824 2911 -23804
rect 2971 -23804 3021 -23764
rect 2971 -23824 3001 -23804
rect 3081 -23854 3141 -23594
rect 3071 -23864 3141 -23854
rect 2741 -23874 2821 -23864
rect 2741 -23934 2751 -23874
rect 2811 -23884 2821 -23874
rect 3061 -23874 3141 -23864
rect 3061 -23884 3071 -23874
rect 2811 -23934 3071 -23884
rect 3131 -23934 3141 -23874
rect 2741 -23944 3141 -23934
rect 3197 -23524 3597 -23514
rect 3197 -23584 3207 -23524
rect 3267 -23574 3527 -23524
rect 3267 -23584 3277 -23574
rect 3197 -23594 3277 -23584
rect 3517 -23584 3527 -23574
rect 3587 -23584 3597 -23524
rect 3517 -23594 3597 -23584
rect 3197 -23864 3257 -23594
rect 3337 -23654 3367 -23634
rect 3317 -23694 3367 -23654
rect 3427 -23654 3457 -23634
rect 3427 -23694 3477 -23654
rect 3317 -23764 3477 -23694
rect 3317 -23804 3367 -23764
rect 3337 -23824 3367 -23804
rect 3427 -23804 3477 -23764
rect 3427 -23824 3457 -23804
rect 3537 -23854 3597 -23594
rect 3527 -23864 3597 -23854
rect 3197 -23874 3277 -23864
rect 3197 -23934 3207 -23874
rect 3267 -23884 3277 -23874
rect 3517 -23874 3597 -23864
rect 3517 -23884 3527 -23874
rect 3267 -23934 3527 -23884
rect 3587 -23934 3597 -23874
rect 3197 -23944 3597 -23934
rect 3653 -23524 4053 -23514
rect 3653 -23584 3663 -23524
rect 3723 -23574 3983 -23524
rect 3723 -23584 3733 -23574
rect 3653 -23594 3733 -23584
rect 3973 -23584 3983 -23574
rect 4043 -23584 4053 -23524
rect 3973 -23594 4053 -23584
rect 3653 -23864 3713 -23594
rect 3793 -23654 3823 -23634
rect 3773 -23694 3823 -23654
rect 3883 -23654 3913 -23634
rect 3883 -23694 3933 -23654
rect 3773 -23764 3933 -23694
rect 3773 -23804 3823 -23764
rect 3793 -23824 3823 -23804
rect 3883 -23804 3933 -23764
rect 3883 -23824 3913 -23804
rect 3993 -23854 4053 -23594
rect 3983 -23864 4053 -23854
rect 3653 -23874 3733 -23864
rect 3653 -23934 3663 -23874
rect 3723 -23884 3733 -23874
rect 3973 -23874 4053 -23864
rect 3973 -23884 3983 -23874
rect 3723 -23934 3983 -23884
rect 4043 -23934 4053 -23874
rect 3653 -23944 4053 -23934
rect 4111 -23524 4511 -23514
rect 4111 -23584 4121 -23524
rect 4181 -23574 4441 -23524
rect 4181 -23584 4191 -23574
rect 4111 -23594 4191 -23584
rect 4431 -23584 4441 -23574
rect 4501 -23584 4511 -23524
rect 4431 -23594 4511 -23584
rect 4111 -23864 4171 -23594
rect 4251 -23654 4281 -23634
rect 4231 -23694 4281 -23654
rect 4341 -23654 4371 -23634
rect 4341 -23694 4391 -23654
rect 4231 -23764 4391 -23694
rect 4231 -23804 4281 -23764
rect 4251 -23824 4281 -23804
rect 4341 -23804 4391 -23764
rect 4341 -23824 4371 -23804
rect 4451 -23854 4511 -23594
rect 4441 -23864 4511 -23854
rect 4111 -23874 4191 -23864
rect 4111 -23934 4121 -23874
rect 4181 -23884 4191 -23874
rect 4431 -23874 4511 -23864
rect 4431 -23884 4441 -23874
rect 4181 -23934 4441 -23884
rect 4501 -23934 4511 -23874
rect 4111 -23944 4511 -23934
rect 4567 -23524 4967 -23514
rect 4567 -23584 4577 -23524
rect 4637 -23574 4897 -23524
rect 4637 -23584 4647 -23574
rect 4567 -23594 4647 -23584
rect 4887 -23584 4897 -23574
rect 4957 -23584 4967 -23524
rect 4887 -23594 4967 -23584
rect 4567 -23864 4627 -23594
rect 4707 -23654 4737 -23634
rect 4687 -23694 4737 -23654
rect 4797 -23654 4827 -23634
rect 4797 -23694 4847 -23654
rect 4687 -23764 4847 -23694
rect 4687 -23804 4737 -23764
rect 4707 -23824 4737 -23804
rect 4797 -23804 4847 -23764
rect 4797 -23824 4827 -23804
rect 4907 -23854 4967 -23594
rect 4897 -23864 4967 -23854
rect 4567 -23874 4647 -23864
rect 4567 -23934 4577 -23874
rect 4637 -23884 4647 -23874
rect 4887 -23874 4967 -23864
rect 4887 -23884 4897 -23874
rect 4637 -23934 4897 -23884
rect 4957 -23934 4967 -23874
rect 4567 -23944 4967 -23934
rect 5023 -23524 5423 -23514
rect 5023 -23584 5033 -23524
rect 5093 -23574 5353 -23524
rect 5093 -23584 5103 -23574
rect 5023 -23594 5103 -23584
rect 5343 -23584 5353 -23574
rect 5413 -23584 5423 -23524
rect 5343 -23594 5423 -23584
rect 5023 -23864 5083 -23594
rect 5163 -23654 5193 -23634
rect 5143 -23694 5193 -23654
rect 5253 -23654 5283 -23634
rect 5253 -23694 5303 -23654
rect 5143 -23764 5303 -23694
rect 5143 -23804 5193 -23764
rect 5163 -23824 5193 -23804
rect 5253 -23804 5303 -23764
rect 5253 -23824 5283 -23804
rect 5363 -23854 5423 -23594
rect 5353 -23864 5423 -23854
rect 5023 -23874 5103 -23864
rect 5023 -23934 5033 -23874
rect 5093 -23884 5103 -23874
rect 5343 -23874 5423 -23864
rect 5343 -23884 5353 -23874
rect 5093 -23934 5353 -23884
rect 5413 -23934 5423 -23874
rect 5023 -23944 5423 -23934
rect 5481 -23524 5881 -23514
rect 5481 -23584 5491 -23524
rect 5551 -23574 5811 -23524
rect 5551 -23584 5561 -23574
rect 5481 -23594 5561 -23584
rect 5801 -23584 5811 -23574
rect 5871 -23584 5881 -23524
rect 5801 -23594 5881 -23584
rect 5481 -23864 5541 -23594
rect 5621 -23654 5651 -23634
rect 5601 -23694 5651 -23654
rect 5711 -23654 5741 -23634
rect 5711 -23694 5761 -23654
rect 5601 -23764 5761 -23694
rect 5601 -23804 5651 -23764
rect 5621 -23824 5651 -23804
rect 5711 -23804 5761 -23764
rect 5711 -23824 5741 -23804
rect 5821 -23854 5881 -23594
rect 5811 -23864 5881 -23854
rect 5481 -23874 5561 -23864
rect 5481 -23934 5491 -23874
rect 5551 -23884 5561 -23874
rect 5801 -23874 5881 -23864
rect 5801 -23884 5811 -23874
rect 5551 -23934 5811 -23884
rect 5871 -23934 5881 -23874
rect 5481 -23944 5881 -23934
rect 5937 -23524 6337 -23514
rect 5937 -23584 5947 -23524
rect 6007 -23574 6267 -23524
rect 6007 -23584 6017 -23574
rect 5937 -23594 6017 -23584
rect 6257 -23584 6267 -23574
rect 6327 -23584 6337 -23524
rect 6257 -23594 6337 -23584
rect 5937 -23864 5997 -23594
rect 6077 -23654 6107 -23634
rect 6057 -23694 6107 -23654
rect 6167 -23654 6197 -23634
rect 6167 -23694 6217 -23654
rect 6057 -23764 6217 -23694
rect 6057 -23804 6107 -23764
rect 6077 -23824 6107 -23804
rect 6167 -23804 6217 -23764
rect 6167 -23824 6197 -23804
rect 6277 -23854 6337 -23594
rect 6267 -23864 6337 -23854
rect 5937 -23874 6017 -23864
rect 5937 -23934 5947 -23874
rect 6007 -23884 6017 -23874
rect 6257 -23874 6337 -23864
rect 6257 -23884 6267 -23874
rect 6007 -23934 6267 -23884
rect 6327 -23934 6337 -23874
rect 5937 -23944 6337 -23934
rect 6393 -23524 6793 -23514
rect 6393 -23584 6403 -23524
rect 6463 -23574 6723 -23524
rect 6463 -23584 6473 -23574
rect 6393 -23594 6473 -23584
rect 6713 -23584 6723 -23574
rect 6783 -23584 6793 -23524
rect 6713 -23594 6793 -23584
rect 6393 -23864 6453 -23594
rect 6533 -23654 6563 -23634
rect 6513 -23694 6563 -23654
rect 6623 -23654 6653 -23634
rect 6623 -23694 6673 -23654
rect 6513 -23764 6673 -23694
rect 6513 -23804 6563 -23764
rect 6533 -23824 6563 -23804
rect 6623 -23804 6673 -23764
rect 6623 -23824 6653 -23804
rect 6733 -23854 6793 -23594
rect 6723 -23864 6793 -23854
rect 6393 -23874 6473 -23864
rect 6393 -23934 6403 -23874
rect 6463 -23884 6473 -23874
rect 6713 -23874 6793 -23864
rect 6713 -23884 6723 -23874
rect 6463 -23934 6723 -23884
rect 6783 -23934 6793 -23874
rect 6393 -23944 6793 -23934
rect 6851 -23524 7251 -23514
rect 6851 -23584 6861 -23524
rect 6921 -23574 7181 -23524
rect 6921 -23584 6931 -23574
rect 6851 -23594 6931 -23584
rect 7171 -23584 7181 -23574
rect 7241 -23584 7251 -23524
rect 7171 -23594 7251 -23584
rect 6851 -23864 6911 -23594
rect 6991 -23654 7021 -23634
rect 6971 -23694 7021 -23654
rect 7081 -23654 7111 -23634
rect 7081 -23694 7131 -23654
rect 6971 -23764 7131 -23694
rect 6971 -23804 7021 -23764
rect 6991 -23824 7021 -23804
rect 7081 -23804 7131 -23764
rect 7081 -23824 7111 -23804
rect 7191 -23854 7251 -23594
rect 7181 -23864 7251 -23854
rect 6851 -23874 6931 -23864
rect 6851 -23934 6861 -23874
rect 6921 -23884 6931 -23874
rect 7171 -23874 7251 -23864
rect 7171 -23884 7181 -23874
rect 6921 -23934 7181 -23884
rect 7241 -23934 7251 -23874
rect 6851 -23944 7251 -23934
rect 7307 -23524 7707 -23514
rect 7307 -23584 7317 -23524
rect 7377 -23574 7637 -23524
rect 7377 -23584 7387 -23574
rect 7307 -23594 7387 -23584
rect 7627 -23584 7637 -23574
rect 7697 -23584 7707 -23524
rect 7627 -23594 7707 -23584
rect 7307 -23864 7367 -23594
rect 7447 -23654 7477 -23634
rect 7427 -23694 7477 -23654
rect 7537 -23654 7567 -23634
rect 7537 -23694 7587 -23654
rect 7427 -23764 7587 -23694
rect 7427 -23804 7477 -23764
rect 7447 -23824 7477 -23804
rect 7537 -23804 7587 -23764
rect 7537 -23824 7567 -23804
rect 7647 -23854 7707 -23594
rect 7637 -23864 7707 -23854
rect 7307 -23874 7387 -23864
rect 7307 -23934 7317 -23874
rect 7377 -23884 7387 -23874
rect 7627 -23874 7707 -23864
rect 7627 -23884 7637 -23874
rect 7377 -23934 7637 -23884
rect 7697 -23934 7707 -23874
rect 7307 -23944 7707 -23934
rect 7763 -23524 8163 -23514
rect 7763 -23584 7773 -23524
rect 7833 -23574 8093 -23524
rect 7833 -23584 7843 -23574
rect 7763 -23594 7843 -23584
rect 8083 -23584 8093 -23574
rect 8153 -23584 8163 -23524
rect 8083 -23594 8163 -23584
rect 7763 -23864 7823 -23594
rect 7903 -23654 7933 -23634
rect 7883 -23694 7933 -23654
rect 7993 -23654 8023 -23634
rect 7993 -23694 8043 -23654
rect 7883 -23764 8043 -23694
rect 7883 -23804 7933 -23764
rect 7903 -23824 7933 -23804
rect 7993 -23804 8043 -23764
rect 7993 -23824 8023 -23804
rect 8103 -23854 8163 -23594
rect 8093 -23864 8163 -23854
rect 7763 -23874 7843 -23864
rect 7763 -23934 7773 -23874
rect 7833 -23884 7843 -23874
rect 8083 -23874 8163 -23864
rect 8083 -23884 8093 -23874
rect 7833 -23934 8093 -23884
rect 8153 -23934 8163 -23874
rect 7763 -23944 8163 -23934
rect 8237 -23524 8637 -23514
rect 8237 -23584 8247 -23524
rect 8307 -23574 8567 -23524
rect 8307 -23584 8317 -23574
rect 8237 -23594 8317 -23584
rect 8557 -23584 8567 -23574
rect 8627 -23584 8637 -23524
rect 8557 -23594 8637 -23584
rect 8237 -23864 8297 -23594
rect 8377 -23654 8407 -23634
rect 8357 -23694 8407 -23654
rect 8467 -23654 8497 -23634
rect 8467 -23694 8517 -23654
rect 8357 -23764 8517 -23694
rect 8357 -23804 8407 -23764
rect 8377 -23824 8407 -23804
rect 8467 -23804 8517 -23764
rect 8467 -23824 8497 -23804
rect 8577 -23854 8637 -23594
rect 8567 -23864 8637 -23854
rect 8237 -23874 8317 -23864
rect 8237 -23934 8247 -23874
rect 8307 -23884 8317 -23874
rect 8557 -23874 8637 -23864
rect 8557 -23884 8567 -23874
rect 8307 -23934 8567 -23884
rect 8627 -23934 8637 -23874
rect 8237 -23944 8637 -23934
rect 8693 -23524 9093 -23514
rect 8693 -23584 8703 -23524
rect 8763 -23574 9023 -23524
rect 8763 -23584 8773 -23574
rect 8693 -23594 8773 -23584
rect 9013 -23584 9023 -23574
rect 9083 -23584 9093 -23524
rect 9013 -23594 9093 -23584
rect 8693 -23864 8753 -23594
rect 8833 -23654 8863 -23634
rect 8813 -23694 8863 -23654
rect 8923 -23654 8953 -23634
rect 8923 -23694 8973 -23654
rect 8813 -23764 8973 -23694
rect 8813 -23804 8863 -23764
rect 8833 -23824 8863 -23804
rect 8923 -23804 8973 -23764
rect 8923 -23824 8953 -23804
rect 9033 -23854 9093 -23594
rect 9023 -23864 9093 -23854
rect 8693 -23874 8773 -23864
rect 8693 -23934 8703 -23874
rect 8763 -23884 8773 -23874
rect 9013 -23874 9093 -23864
rect 9013 -23884 9023 -23874
rect 8763 -23934 9023 -23884
rect 9083 -23934 9093 -23874
rect 8693 -23944 9093 -23934
rect 9151 -23524 9551 -23514
rect 9151 -23584 9161 -23524
rect 9221 -23574 9481 -23524
rect 9221 -23584 9231 -23574
rect 9151 -23594 9231 -23584
rect 9471 -23584 9481 -23574
rect 9541 -23584 9551 -23524
rect 9471 -23594 9551 -23584
rect 9151 -23864 9211 -23594
rect 9291 -23654 9321 -23634
rect 9271 -23694 9321 -23654
rect 9381 -23654 9411 -23634
rect 9381 -23694 9431 -23654
rect 9271 -23764 9431 -23694
rect 9271 -23804 9321 -23764
rect 9291 -23824 9321 -23804
rect 9381 -23804 9431 -23764
rect 9381 -23824 9411 -23804
rect 9491 -23854 9551 -23594
rect 9481 -23864 9551 -23854
rect 9151 -23874 9231 -23864
rect 9151 -23934 9161 -23874
rect 9221 -23884 9231 -23874
rect 9471 -23874 9551 -23864
rect 9471 -23884 9481 -23874
rect 9221 -23934 9481 -23884
rect 9541 -23934 9551 -23874
rect 9151 -23944 9551 -23934
rect 9607 -23524 10007 -23514
rect 9607 -23584 9617 -23524
rect 9677 -23574 9937 -23524
rect 9677 -23584 9687 -23574
rect 9607 -23594 9687 -23584
rect 9927 -23584 9937 -23574
rect 9997 -23584 10007 -23524
rect 9927 -23594 10007 -23584
rect 9607 -23864 9667 -23594
rect 9747 -23654 9777 -23634
rect 9727 -23694 9777 -23654
rect 9837 -23654 9867 -23634
rect 9837 -23694 9887 -23654
rect 9727 -23764 9887 -23694
rect 9727 -23804 9777 -23764
rect 9747 -23824 9777 -23804
rect 9837 -23804 9887 -23764
rect 9837 -23824 9867 -23804
rect 9947 -23854 10007 -23594
rect 9937 -23864 10007 -23854
rect 9607 -23874 9687 -23864
rect 9607 -23934 9617 -23874
rect 9677 -23884 9687 -23874
rect 9927 -23874 10007 -23864
rect 9927 -23884 9937 -23874
rect 9677 -23934 9937 -23884
rect 9997 -23934 10007 -23874
rect 9607 -23944 10007 -23934
rect 10063 -23524 10463 -23514
rect 10063 -23584 10073 -23524
rect 10133 -23574 10393 -23524
rect 10133 -23584 10143 -23574
rect 10063 -23594 10143 -23584
rect 10383 -23584 10393 -23574
rect 10453 -23584 10463 -23524
rect 10383 -23594 10463 -23584
rect 10063 -23864 10123 -23594
rect 10203 -23654 10233 -23634
rect 10183 -23694 10233 -23654
rect 10293 -23654 10323 -23634
rect 10293 -23694 10343 -23654
rect 10183 -23764 10343 -23694
rect 10183 -23804 10233 -23764
rect 10203 -23824 10233 -23804
rect 10293 -23804 10343 -23764
rect 10293 -23824 10323 -23804
rect 10403 -23854 10463 -23594
rect 10393 -23864 10463 -23854
rect 10063 -23874 10143 -23864
rect 10063 -23934 10073 -23874
rect 10133 -23884 10143 -23874
rect 10383 -23874 10463 -23864
rect 10383 -23884 10393 -23874
rect 10133 -23934 10393 -23884
rect 10453 -23934 10463 -23874
rect 10063 -23944 10463 -23934
rect 10521 -23524 10921 -23514
rect 10521 -23584 10531 -23524
rect 10591 -23574 10851 -23524
rect 10591 -23584 10601 -23574
rect 10521 -23594 10601 -23584
rect 10841 -23584 10851 -23574
rect 10911 -23584 10921 -23524
rect 10841 -23594 10921 -23584
rect 10521 -23864 10581 -23594
rect 10661 -23654 10691 -23634
rect 10641 -23694 10691 -23654
rect 10751 -23654 10781 -23634
rect 10751 -23694 10801 -23654
rect 10641 -23764 10801 -23694
rect 10641 -23804 10691 -23764
rect 10661 -23824 10691 -23804
rect 10751 -23804 10801 -23764
rect 10751 -23824 10781 -23804
rect 10861 -23854 10921 -23594
rect 10851 -23864 10921 -23854
rect 10521 -23874 10601 -23864
rect 10521 -23934 10531 -23874
rect 10591 -23884 10601 -23874
rect 10841 -23874 10921 -23864
rect 10841 -23884 10851 -23874
rect 10591 -23934 10851 -23884
rect 10911 -23934 10921 -23874
rect 10521 -23944 10921 -23934
rect 10977 -23524 11377 -23514
rect 10977 -23584 10987 -23524
rect 11047 -23574 11307 -23524
rect 11047 -23584 11057 -23574
rect 10977 -23594 11057 -23584
rect 11297 -23584 11307 -23574
rect 11367 -23584 11377 -23524
rect 11297 -23594 11377 -23584
rect 10977 -23864 11037 -23594
rect 11117 -23654 11147 -23634
rect 11097 -23694 11147 -23654
rect 11207 -23654 11237 -23634
rect 11207 -23694 11257 -23654
rect 11097 -23764 11257 -23694
rect 11097 -23804 11147 -23764
rect 11117 -23824 11147 -23804
rect 11207 -23804 11257 -23764
rect 11207 -23824 11237 -23804
rect 11317 -23854 11377 -23594
rect 11307 -23864 11377 -23854
rect 10977 -23874 11057 -23864
rect 10977 -23934 10987 -23874
rect 11047 -23884 11057 -23874
rect 11297 -23874 11377 -23864
rect 11297 -23884 11307 -23874
rect 11047 -23934 11307 -23884
rect 11367 -23934 11377 -23874
rect 10977 -23944 11377 -23934
rect 11433 -23524 11833 -23514
rect 11433 -23584 11443 -23524
rect 11503 -23574 11763 -23524
rect 11503 -23584 11513 -23574
rect 11433 -23594 11513 -23584
rect 11753 -23584 11763 -23574
rect 11823 -23584 11833 -23524
rect 11753 -23594 11833 -23584
rect 11433 -23864 11493 -23594
rect 11573 -23654 11603 -23634
rect 11553 -23694 11603 -23654
rect 11663 -23654 11693 -23634
rect 11663 -23694 11713 -23654
rect 11553 -23764 11713 -23694
rect 11553 -23804 11603 -23764
rect 11573 -23824 11603 -23804
rect 11663 -23804 11713 -23764
rect 11663 -23824 11693 -23804
rect 11773 -23854 11833 -23594
rect 11763 -23864 11833 -23854
rect 11433 -23874 11513 -23864
rect 11433 -23934 11443 -23874
rect 11503 -23884 11513 -23874
rect 11753 -23874 11833 -23864
rect 11753 -23884 11763 -23874
rect 11503 -23934 11763 -23884
rect 11823 -23934 11833 -23874
rect 11433 -23944 11833 -23934
rect 11891 -23524 12291 -23514
rect 11891 -23584 11901 -23524
rect 11961 -23574 12221 -23524
rect 11961 -23584 11971 -23574
rect 11891 -23594 11971 -23584
rect 12211 -23584 12221 -23574
rect 12281 -23584 12291 -23524
rect 12211 -23594 12291 -23584
rect 11891 -23864 11951 -23594
rect 12031 -23654 12061 -23634
rect 12011 -23694 12061 -23654
rect 12121 -23654 12151 -23634
rect 12121 -23694 12171 -23654
rect 12011 -23764 12171 -23694
rect 12011 -23804 12061 -23764
rect 12031 -23824 12061 -23804
rect 12121 -23804 12171 -23764
rect 12121 -23824 12151 -23804
rect 12231 -23854 12291 -23594
rect 12221 -23864 12291 -23854
rect 11891 -23874 11971 -23864
rect 11891 -23934 11901 -23874
rect 11961 -23884 11971 -23874
rect 12211 -23874 12291 -23864
rect 12211 -23884 12221 -23874
rect 11961 -23934 12221 -23884
rect 12281 -23934 12291 -23874
rect 11891 -23944 12291 -23934
rect 12347 -23524 12747 -23514
rect 12347 -23584 12357 -23524
rect 12417 -23574 12677 -23524
rect 12417 -23584 12427 -23574
rect 12347 -23594 12427 -23584
rect 12667 -23584 12677 -23574
rect 12737 -23584 12747 -23524
rect 12667 -23594 12747 -23584
rect 12347 -23864 12407 -23594
rect 12487 -23654 12517 -23634
rect 12467 -23694 12517 -23654
rect 12577 -23654 12607 -23634
rect 12577 -23694 12627 -23654
rect 12467 -23764 12627 -23694
rect 12467 -23804 12517 -23764
rect 12487 -23824 12517 -23804
rect 12577 -23804 12627 -23764
rect 12577 -23824 12607 -23804
rect 12687 -23854 12747 -23594
rect 12677 -23864 12747 -23854
rect 12347 -23874 12427 -23864
rect 12347 -23934 12357 -23874
rect 12417 -23884 12427 -23874
rect 12667 -23874 12747 -23864
rect 12667 -23884 12677 -23874
rect 12417 -23934 12677 -23884
rect 12737 -23934 12747 -23874
rect 12347 -23944 12747 -23934
rect 12803 -23524 13203 -23514
rect 12803 -23584 12813 -23524
rect 12873 -23574 13133 -23524
rect 12873 -23584 12883 -23574
rect 12803 -23594 12883 -23584
rect 13123 -23584 13133 -23574
rect 13193 -23584 13203 -23524
rect 13123 -23594 13203 -23584
rect 12803 -23864 12863 -23594
rect 12943 -23654 12973 -23634
rect 12923 -23694 12973 -23654
rect 13033 -23654 13063 -23634
rect 13033 -23694 13083 -23654
rect 12923 -23764 13083 -23694
rect 12923 -23804 12973 -23764
rect 12943 -23824 12973 -23804
rect 13033 -23804 13083 -23764
rect 13033 -23824 13063 -23804
rect 13143 -23854 13203 -23594
rect 13133 -23864 13203 -23854
rect 12803 -23874 12883 -23864
rect 12803 -23934 12813 -23874
rect 12873 -23884 12883 -23874
rect 13123 -23874 13203 -23864
rect 13123 -23884 13133 -23874
rect 12873 -23934 13133 -23884
rect 13193 -23934 13203 -23874
rect 12803 -23944 13203 -23934
rect 13261 -23524 13661 -23514
rect 13261 -23584 13271 -23524
rect 13331 -23574 13591 -23524
rect 13331 -23584 13341 -23574
rect 13261 -23594 13341 -23584
rect 13581 -23584 13591 -23574
rect 13651 -23584 13661 -23524
rect 13581 -23594 13661 -23584
rect 13261 -23864 13321 -23594
rect 13401 -23654 13431 -23634
rect 13381 -23694 13431 -23654
rect 13491 -23654 13521 -23634
rect 13491 -23694 13541 -23654
rect 13381 -23764 13541 -23694
rect 13381 -23804 13431 -23764
rect 13401 -23824 13431 -23804
rect 13491 -23804 13541 -23764
rect 13491 -23824 13521 -23804
rect 13601 -23854 13661 -23594
rect 13591 -23864 13661 -23854
rect 13261 -23874 13341 -23864
rect 13261 -23934 13271 -23874
rect 13331 -23884 13341 -23874
rect 13581 -23874 13661 -23864
rect 13581 -23884 13591 -23874
rect 13331 -23934 13591 -23884
rect 13651 -23934 13661 -23874
rect 13261 -23944 13661 -23934
rect 13717 -23524 14117 -23514
rect 13717 -23584 13727 -23524
rect 13787 -23574 14047 -23524
rect 13787 -23584 13797 -23574
rect 13717 -23594 13797 -23584
rect 14037 -23584 14047 -23574
rect 14107 -23584 14117 -23524
rect 14037 -23594 14117 -23584
rect 13717 -23864 13777 -23594
rect 13857 -23654 13887 -23634
rect 13837 -23694 13887 -23654
rect 13947 -23654 13977 -23634
rect 13947 -23694 13997 -23654
rect 13837 -23764 13997 -23694
rect 13837 -23804 13887 -23764
rect 13857 -23824 13887 -23804
rect 13947 -23804 13997 -23764
rect 13947 -23824 13977 -23804
rect 14057 -23854 14117 -23594
rect 14047 -23864 14117 -23854
rect 13717 -23874 13797 -23864
rect 13717 -23934 13727 -23874
rect 13787 -23884 13797 -23874
rect 14037 -23874 14117 -23864
rect 14037 -23884 14047 -23874
rect 13787 -23934 14047 -23884
rect 14107 -23934 14117 -23874
rect 13717 -23944 14117 -23934
rect 14173 -23524 14573 -23514
rect 14173 -23584 14183 -23524
rect 14243 -23574 14503 -23524
rect 14243 -23584 14253 -23574
rect 14173 -23594 14253 -23584
rect 14493 -23584 14503 -23574
rect 14563 -23584 14573 -23524
rect 14493 -23594 14573 -23584
rect 14173 -23864 14233 -23594
rect 14313 -23654 14343 -23634
rect 14293 -23694 14343 -23654
rect 14403 -23654 14433 -23634
rect 14403 -23694 14453 -23654
rect 14293 -23764 14453 -23694
rect 14293 -23804 14343 -23764
rect 14313 -23824 14343 -23804
rect 14403 -23804 14453 -23764
rect 14403 -23824 14433 -23804
rect 14513 -23854 14573 -23594
rect 14503 -23864 14573 -23854
rect 14173 -23874 14253 -23864
rect 14173 -23934 14183 -23874
rect 14243 -23884 14253 -23874
rect 14493 -23874 14573 -23864
rect 14493 -23884 14503 -23874
rect 14243 -23934 14503 -23884
rect 14563 -23934 14573 -23874
rect 14173 -23944 14573 -23934
rect 14631 -23524 15031 -23514
rect 14631 -23584 14641 -23524
rect 14701 -23574 14961 -23524
rect 14701 -23584 14711 -23574
rect 14631 -23594 14711 -23584
rect 14951 -23584 14961 -23574
rect 15021 -23584 15031 -23524
rect 14951 -23594 15031 -23584
rect 14631 -23864 14691 -23594
rect 14771 -23654 14801 -23634
rect 14751 -23694 14801 -23654
rect 14861 -23654 14891 -23634
rect 14861 -23694 14911 -23654
rect 14751 -23764 14911 -23694
rect 14751 -23804 14801 -23764
rect 14771 -23824 14801 -23804
rect 14861 -23804 14911 -23764
rect 14861 -23824 14891 -23804
rect 14971 -23854 15031 -23594
rect 14961 -23864 15031 -23854
rect 14631 -23874 14711 -23864
rect 14631 -23934 14641 -23874
rect 14701 -23884 14711 -23874
rect 14951 -23874 15031 -23864
rect 14951 -23884 14961 -23874
rect 14701 -23934 14961 -23884
rect 15021 -23934 15031 -23874
rect 14631 -23944 15031 -23934
rect 15087 -23524 15487 -23514
rect 15087 -23584 15097 -23524
rect 15157 -23574 15417 -23524
rect 15157 -23584 15167 -23574
rect 15087 -23594 15167 -23584
rect 15407 -23584 15417 -23574
rect 15477 -23584 15487 -23524
rect 15407 -23594 15487 -23584
rect 15087 -23864 15147 -23594
rect 15227 -23654 15257 -23634
rect 15207 -23694 15257 -23654
rect 15317 -23654 15347 -23634
rect 15317 -23694 15367 -23654
rect 15207 -23764 15367 -23694
rect 15207 -23804 15257 -23764
rect 15227 -23824 15257 -23804
rect 15317 -23804 15367 -23764
rect 15317 -23824 15347 -23804
rect 15427 -23854 15487 -23594
rect 15417 -23864 15487 -23854
rect 15087 -23874 15167 -23864
rect 15087 -23934 15097 -23874
rect 15157 -23884 15167 -23874
rect 15407 -23874 15487 -23864
rect 15407 -23884 15417 -23874
rect 15157 -23934 15417 -23884
rect 15477 -23934 15487 -23874
rect 15087 -23944 15487 -23934
rect 1 -24016 401 -24006
rect 1 -24076 11 -24016
rect 71 -24066 331 -24016
rect 71 -24076 81 -24066
rect 1 -24086 81 -24076
rect 321 -24076 331 -24066
rect 391 -24076 401 -24016
rect 321 -24086 401 -24076
rect 1 -24356 61 -24086
rect 141 -24146 171 -24126
rect 121 -24186 171 -24146
rect 231 -24146 261 -24126
rect 231 -24186 281 -24146
rect 121 -24256 281 -24186
rect 121 -24296 171 -24256
rect 141 -24316 171 -24296
rect 231 -24296 281 -24256
rect 231 -24316 261 -24296
rect 341 -24346 401 -24086
rect 331 -24356 401 -24346
rect 1 -24366 81 -24356
rect 1 -24426 11 -24366
rect 71 -24376 81 -24366
rect 321 -24366 401 -24356
rect 321 -24376 331 -24366
rect 71 -24426 331 -24376
rect 391 -24426 401 -24366
rect 1 -24436 401 -24426
rect 457 -24016 857 -24006
rect 457 -24076 467 -24016
rect 527 -24066 787 -24016
rect 527 -24076 537 -24066
rect 457 -24086 537 -24076
rect 777 -24076 787 -24066
rect 847 -24076 857 -24016
rect 777 -24086 857 -24076
rect 457 -24356 517 -24086
rect 597 -24146 627 -24126
rect 577 -24186 627 -24146
rect 687 -24146 717 -24126
rect 687 -24186 737 -24146
rect 577 -24256 737 -24186
rect 577 -24296 627 -24256
rect 597 -24316 627 -24296
rect 687 -24296 737 -24256
rect 687 -24316 717 -24296
rect 797 -24346 857 -24086
rect 787 -24356 857 -24346
rect 457 -24366 537 -24356
rect 457 -24426 467 -24366
rect 527 -24376 537 -24366
rect 777 -24366 857 -24356
rect 777 -24376 787 -24366
rect 527 -24426 787 -24376
rect 847 -24426 857 -24366
rect 457 -24436 857 -24426
rect 913 -24016 1313 -24006
rect 913 -24076 923 -24016
rect 983 -24066 1243 -24016
rect 983 -24076 993 -24066
rect 913 -24086 993 -24076
rect 1233 -24076 1243 -24066
rect 1303 -24076 1313 -24016
rect 1233 -24086 1313 -24076
rect 913 -24356 973 -24086
rect 1053 -24146 1083 -24126
rect 1033 -24186 1083 -24146
rect 1143 -24146 1173 -24126
rect 1143 -24186 1193 -24146
rect 1033 -24256 1193 -24186
rect 1033 -24296 1083 -24256
rect 1053 -24316 1083 -24296
rect 1143 -24296 1193 -24256
rect 1143 -24316 1173 -24296
rect 1253 -24346 1313 -24086
rect 1243 -24356 1313 -24346
rect 913 -24366 993 -24356
rect 913 -24426 923 -24366
rect 983 -24376 993 -24366
rect 1233 -24366 1313 -24356
rect 1233 -24376 1243 -24366
rect 983 -24426 1243 -24376
rect 1303 -24426 1313 -24366
rect 913 -24436 1313 -24426
rect 1371 -24016 1771 -24006
rect 1371 -24076 1381 -24016
rect 1441 -24066 1701 -24016
rect 1441 -24076 1451 -24066
rect 1371 -24086 1451 -24076
rect 1691 -24076 1701 -24066
rect 1761 -24076 1771 -24016
rect 1691 -24086 1771 -24076
rect 1371 -24356 1431 -24086
rect 1511 -24146 1541 -24126
rect 1491 -24186 1541 -24146
rect 1601 -24146 1631 -24126
rect 1601 -24186 1651 -24146
rect 1491 -24256 1651 -24186
rect 1491 -24296 1541 -24256
rect 1511 -24316 1541 -24296
rect 1601 -24296 1651 -24256
rect 1601 -24316 1631 -24296
rect 1711 -24346 1771 -24086
rect 1701 -24356 1771 -24346
rect 1371 -24366 1451 -24356
rect 1371 -24426 1381 -24366
rect 1441 -24376 1451 -24366
rect 1691 -24366 1771 -24356
rect 1691 -24376 1701 -24366
rect 1441 -24426 1701 -24376
rect 1761 -24426 1771 -24366
rect 1371 -24436 1771 -24426
rect 1827 -24016 2227 -24006
rect 1827 -24076 1837 -24016
rect 1897 -24066 2157 -24016
rect 1897 -24076 1907 -24066
rect 1827 -24086 1907 -24076
rect 2147 -24076 2157 -24066
rect 2217 -24076 2227 -24016
rect 2147 -24086 2227 -24076
rect 1827 -24356 1887 -24086
rect 1967 -24146 1997 -24126
rect 1947 -24186 1997 -24146
rect 2057 -24146 2087 -24126
rect 2057 -24186 2107 -24146
rect 1947 -24256 2107 -24186
rect 1947 -24296 1997 -24256
rect 1967 -24316 1997 -24296
rect 2057 -24296 2107 -24256
rect 2057 -24316 2087 -24296
rect 2167 -24346 2227 -24086
rect 2157 -24356 2227 -24346
rect 1827 -24366 1907 -24356
rect 1827 -24426 1837 -24366
rect 1897 -24376 1907 -24366
rect 2147 -24366 2227 -24356
rect 2147 -24376 2157 -24366
rect 1897 -24426 2157 -24376
rect 2217 -24426 2227 -24366
rect 1827 -24436 2227 -24426
rect 2283 -24016 2683 -24006
rect 2283 -24076 2293 -24016
rect 2353 -24066 2613 -24016
rect 2353 -24076 2363 -24066
rect 2283 -24086 2363 -24076
rect 2603 -24076 2613 -24066
rect 2673 -24076 2683 -24016
rect 2603 -24086 2683 -24076
rect 2283 -24356 2343 -24086
rect 2423 -24146 2453 -24126
rect 2403 -24186 2453 -24146
rect 2513 -24146 2543 -24126
rect 2513 -24186 2563 -24146
rect 2403 -24256 2563 -24186
rect 2403 -24296 2453 -24256
rect 2423 -24316 2453 -24296
rect 2513 -24296 2563 -24256
rect 2513 -24316 2543 -24296
rect 2623 -24346 2683 -24086
rect 2613 -24356 2683 -24346
rect 2283 -24366 2363 -24356
rect 2283 -24426 2293 -24366
rect 2353 -24376 2363 -24366
rect 2603 -24366 2683 -24356
rect 2603 -24376 2613 -24366
rect 2353 -24426 2613 -24376
rect 2673 -24426 2683 -24366
rect 2283 -24436 2683 -24426
rect 2741 -24016 3141 -24006
rect 2741 -24076 2751 -24016
rect 2811 -24066 3071 -24016
rect 2811 -24076 2821 -24066
rect 2741 -24086 2821 -24076
rect 3061 -24076 3071 -24066
rect 3131 -24076 3141 -24016
rect 3061 -24086 3141 -24076
rect 2741 -24356 2801 -24086
rect 2881 -24146 2911 -24126
rect 2861 -24186 2911 -24146
rect 2971 -24146 3001 -24126
rect 2971 -24186 3021 -24146
rect 2861 -24256 3021 -24186
rect 2861 -24296 2911 -24256
rect 2881 -24316 2911 -24296
rect 2971 -24296 3021 -24256
rect 2971 -24316 3001 -24296
rect 3081 -24346 3141 -24086
rect 3071 -24356 3141 -24346
rect 2741 -24366 2821 -24356
rect 2741 -24426 2751 -24366
rect 2811 -24376 2821 -24366
rect 3061 -24366 3141 -24356
rect 3061 -24376 3071 -24366
rect 2811 -24426 3071 -24376
rect 3131 -24426 3141 -24366
rect 2741 -24436 3141 -24426
rect 3197 -24016 3597 -24006
rect 3197 -24076 3207 -24016
rect 3267 -24066 3527 -24016
rect 3267 -24076 3277 -24066
rect 3197 -24086 3277 -24076
rect 3517 -24076 3527 -24066
rect 3587 -24076 3597 -24016
rect 3517 -24086 3597 -24076
rect 3197 -24356 3257 -24086
rect 3337 -24146 3367 -24126
rect 3317 -24186 3367 -24146
rect 3427 -24146 3457 -24126
rect 3427 -24186 3477 -24146
rect 3317 -24256 3477 -24186
rect 3317 -24296 3367 -24256
rect 3337 -24316 3367 -24296
rect 3427 -24296 3477 -24256
rect 3427 -24316 3457 -24296
rect 3537 -24346 3597 -24086
rect 3527 -24356 3597 -24346
rect 3197 -24366 3277 -24356
rect 3197 -24426 3207 -24366
rect 3267 -24376 3277 -24366
rect 3517 -24366 3597 -24356
rect 3517 -24376 3527 -24366
rect 3267 -24426 3527 -24376
rect 3587 -24426 3597 -24366
rect 3197 -24436 3597 -24426
rect 3653 -24016 4053 -24006
rect 3653 -24076 3663 -24016
rect 3723 -24066 3983 -24016
rect 3723 -24076 3733 -24066
rect 3653 -24086 3733 -24076
rect 3973 -24076 3983 -24066
rect 4043 -24076 4053 -24016
rect 3973 -24086 4053 -24076
rect 3653 -24356 3713 -24086
rect 3793 -24146 3823 -24126
rect 3773 -24186 3823 -24146
rect 3883 -24146 3913 -24126
rect 3883 -24186 3933 -24146
rect 3773 -24256 3933 -24186
rect 3773 -24296 3823 -24256
rect 3793 -24316 3823 -24296
rect 3883 -24296 3933 -24256
rect 3883 -24316 3913 -24296
rect 3993 -24346 4053 -24086
rect 3983 -24356 4053 -24346
rect 3653 -24366 3733 -24356
rect 3653 -24426 3663 -24366
rect 3723 -24376 3733 -24366
rect 3973 -24366 4053 -24356
rect 3973 -24376 3983 -24366
rect 3723 -24426 3983 -24376
rect 4043 -24426 4053 -24366
rect 3653 -24436 4053 -24426
rect 4111 -24016 4511 -24006
rect 4111 -24076 4121 -24016
rect 4181 -24066 4441 -24016
rect 4181 -24076 4191 -24066
rect 4111 -24086 4191 -24076
rect 4431 -24076 4441 -24066
rect 4501 -24076 4511 -24016
rect 4431 -24086 4511 -24076
rect 4111 -24356 4171 -24086
rect 4251 -24146 4281 -24126
rect 4231 -24186 4281 -24146
rect 4341 -24146 4371 -24126
rect 4341 -24186 4391 -24146
rect 4231 -24256 4391 -24186
rect 4231 -24296 4281 -24256
rect 4251 -24316 4281 -24296
rect 4341 -24296 4391 -24256
rect 4341 -24316 4371 -24296
rect 4451 -24346 4511 -24086
rect 4441 -24356 4511 -24346
rect 4111 -24366 4191 -24356
rect 4111 -24426 4121 -24366
rect 4181 -24376 4191 -24366
rect 4431 -24366 4511 -24356
rect 4431 -24376 4441 -24366
rect 4181 -24426 4441 -24376
rect 4501 -24426 4511 -24366
rect 4111 -24436 4511 -24426
rect 4567 -24016 4967 -24006
rect 4567 -24076 4577 -24016
rect 4637 -24066 4897 -24016
rect 4637 -24076 4647 -24066
rect 4567 -24086 4647 -24076
rect 4887 -24076 4897 -24066
rect 4957 -24076 4967 -24016
rect 4887 -24086 4967 -24076
rect 4567 -24356 4627 -24086
rect 4707 -24146 4737 -24126
rect 4687 -24186 4737 -24146
rect 4797 -24146 4827 -24126
rect 4797 -24186 4847 -24146
rect 4687 -24256 4847 -24186
rect 4687 -24296 4737 -24256
rect 4707 -24316 4737 -24296
rect 4797 -24296 4847 -24256
rect 4797 -24316 4827 -24296
rect 4907 -24346 4967 -24086
rect 4897 -24356 4967 -24346
rect 4567 -24366 4647 -24356
rect 4567 -24426 4577 -24366
rect 4637 -24376 4647 -24366
rect 4887 -24366 4967 -24356
rect 4887 -24376 4897 -24366
rect 4637 -24426 4897 -24376
rect 4957 -24426 4967 -24366
rect 4567 -24436 4967 -24426
rect 5023 -24016 5423 -24006
rect 5023 -24076 5033 -24016
rect 5093 -24066 5353 -24016
rect 5093 -24076 5103 -24066
rect 5023 -24086 5103 -24076
rect 5343 -24076 5353 -24066
rect 5413 -24076 5423 -24016
rect 5343 -24086 5423 -24076
rect 5023 -24356 5083 -24086
rect 5163 -24146 5193 -24126
rect 5143 -24186 5193 -24146
rect 5253 -24146 5283 -24126
rect 5253 -24186 5303 -24146
rect 5143 -24256 5303 -24186
rect 5143 -24296 5193 -24256
rect 5163 -24316 5193 -24296
rect 5253 -24296 5303 -24256
rect 5253 -24316 5283 -24296
rect 5363 -24346 5423 -24086
rect 5353 -24356 5423 -24346
rect 5023 -24366 5103 -24356
rect 5023 -24426 5033 -24366
rect 5093 -24376 5103 -24366
rect 5343 -24366 5423 -24356
rect 5343 -24376 5353 -24366
rect 5093 -24426 5353 -24376
rect 5413 -24426 5423 -24366
rect 5023 -24436 5423 -24426
rect 5481 -24016 5881 -24006
rect 5481 -24076 5491 -24016
rect 5551 -24066 5811 -24016
rect 5551 -24076 5561 -24066
rect 5481 -24086 5561 -24076
rect 5801 -24076 5811 -24066
rect 5871 -24076 5881 -24016
rect 5801 -24086 5881 -24076
rect 5481 -24356 5541 -24086
rect 5621 -24146 5651 -24126
rect 5601 -24186 5651 -24146
rect 5711 -24146 5741 -24126
rect 5711 -24186 5761 -24146
rect 5601 -24256 5761 -24186
rect 5601 -24296 5651 -24256
rect 5621 -24316 5651 -24296
rect 5711 -24296 5761 -24256
rect 5711 -24316 5741 -24296
rect 5821 -24346 5881 -24086
rect 5811 -24356 5881 -24346
rect 5481 -24366 5561 -24356
rect 5481 -24426 5491 -24366
rect 5551 -24376 5561 -24366
rect 5801 -24366 5881 -24356
rect 5801 -24376 5811 -24366
rect 5551 -24426 5811 -24376
rect 5871 -24426 5881 -24366
rect 5481 -24436 5881 -24426
rect 5937 -24016 6337 -24006
rect 5937 -24076 5947 -24016
rect 6007 -24066 6267 -24016
rect 6007 -24076 6017 -24066
rect 5937 -24086 6017 -24076
rect 6257 -24076 6267 -24066
rect 6327 -24076 6337 -24016
rect 6257 -24086 6337 -24076
rect 5937 -24356 5997 -24086
rect 6077 -24146 6107 -24126
rect 6057 -24186 6107 -24146
rect 6167 -24146 6197 -24126
rect 6167 -24186 6217 -24146
rect 6057 -24256 6217 -24186
rect 6057 -24296 6107 -24256
rect 6077 -24316 6107 -24296
rect 6167 -24296 6217 -24256
rect 6167 -24316 6197 -24296
rect 6277 -24346 6337 -24086
rect 6267 -24356 6337 -24346
rect 5937 -24366 6017 -24356
rect 5937 -24426 5947 -24366
rect 6007 -24376 6017 -24366
rect 6257 -24366 6337 -24356
rect 6257 -24376 6267 -24366
rect 6007 -24426 6267 -24376
rect 6327 -24426 6337 -24366
rect 5937 -24436 6337 -24426
rect 6393 -24016 6793 -24006
rect 6393 -24076 6403 -24016
rect 6463 -24066 6723 -24016
rect 6463 -24076 6473 -24066
rect 6393 -24086 6473 -24076
rect 6713 -24076 6723 -24066
rect 6783 -24076 6793 -24016
rect 6713 -24086 6793 -24076
rect 6393 -24356 6453 -24086
rect 6533 -24146 6563 -24126
rect 6513 -24186 6563 -24146
rect 6623 -24146 6653 -24126
rect 6623 -24186 6673 -24146
rect 6513 -24256 6673 -24186
rect 6513 -24296 6563 -24256
rect 6533 -24316 6563 -24296
rect 6623 -24296 6673 -24256
rect 6623 -24316 6653 -24296
rect 6733 -24346 6793 -24086
rect 6723 -24356 6793 -24346
rect 6393 -24366 6473 -24356
rect 6393 -24426 6403 -24366
rect 6463 -24376 6473 -24366
rect 6713 -24366 6793 -24356
rect 6713 -24376 6723 -24366
rect 6463 -24426 6723 -24376
rect 6783 -24426 6793 -24366
rect 6393 -24436 6793 -24426
rect 6851 -24016 7251 -24006
rect 6851 -24076 6861 -24016
rect 6921 -24066 7181 -24016
rect 6921 -24076 6931 -24066
rect 6851 -24086 6931 -24076
rect 7171 -24076 7181 -24066
rect 7241 -24076 7251 -24016
rect 7171 -24086 7251 -24076
rect 6851 -24356 6911 -24086
rect 6991 -24146 7021 -24126
rect 6971 -24186 7021 -24146
rect 7081 -24146 7111 -24126
rect 7081 -24186 7131 -24146
rect 6971 -24256 7131 -24186
rect 6971 -24296 7021 -24256
rect 6991 -24316 7021 -24296
rect 7081 -24296 7131 -24256
rect 7081 -24316 7111 -24296
rect 7191 -24346 7251 -24086
rect 7181 -24356 7251 -24346
rect 6851 -24366 6931 -24356
rect 6851 -24426 6861 -24366
rect 6921 -24376 6931 -24366
rect 7171 -24366 7251 -24356
rect 7171 -24376 7181 -24366
rect 6921 -24426 7181 -24376
rect 7241 -24426 7251 -24366
rect 6851 -24436 7251 -24426
rect 7307 -24016 7707 -24006
rect 7307 -24076 7317 -24016
rect 7377 -24066 7637 -24016
rect 7377 -24076 7387 -24066
rect 7307 -24086 7387 -24076
rect 7627 -24076 7637 -24066
rect 7697 -24076 7707 -24016
rect 7627 -24086 7707 -24076
rect 7307 -24356 7367 -24086
rect 7447 -24146 7477 -24126
rect 7427 -24186 7477 -24146
rect 7537 -24146 7567 -24126
rect 7537 -24186 7587 -24146
rect 7427 -24256 7587 -24186
rect 7427 -24296 7477 -24256
rect 7447 -24316 7477 -24296
rect 7537 -24296 7587 -24256
rect 7537 -24316 7567 -24296
rect 7647 -24346 7707 -24086
rect 7637 -24356 7707 -24346
rect 7307 -24366 7387 -24356
rect 7307 -24426 7317 -24366
rect 7377 -24376 7387 -24366
rect 7627 -24366 7707 -24356
rect 7627 -24376 7637 -24366
rect 7377 -24426 7637 -24376
rect 7697 -24426 7707 -24366
rect 7307 -24436 7707 -24426
rect 7763 -24016 8163 -24006
rect 7763 -24076 7773 -24016
rect 7833 -24066 8093 -24016
rect 7833 -24076 7843 -24066
rect 7763 -24086 7843 -24076
rect 8083 -24076 8093 -24066
rect 8153 -24076 8163 -24016
rect 8083 -24086 8163 -24076
rect 7763 -24356 7823 -24086
rect 7903 -24146 7933 -24126
rect 7883 -24186 7933 -24146
rect 7993 -24146 8023 -24126
rect 7993 -24186 8043 -24146
rect 7883 -24256 8043 -24186
rect 7883 -24296 7933 -24256
rect 7903 -24316 7933 -24296
rect 7993 -24296 8043 -24256
rect 7993 -24316 8023 -24296
rect 8103 -24346 8163 -24086
rect 8093 -24356 8163 -24346
rect 7763 -24366 7843 -24356
rect 7763 -24426 7773 -24366
rect 7833 -24376 7843 -24366
rect 8083 -24366 8163 -24356
rect 8083 -24376 8093 -24366
rect 7833 -24426 8093 -24376
rect 8153 -24426 8163 -24366
rect 7763 -24436 8163 -24426
rect 8237 -24016 8637 -24006
rect 8237 -24076 8247 -24016
rect 8307 -24066 8567 -24016
rect 8307 -24076 8317 -24066
rect 8237 -24086 8317 -24076
rect 8557 -24076 8567 -24066
rect 8627 -24076 8637 -24016
rect 8557 -24086 8637 -24076
rect 8237 -24356 8297 -24086
rect 8377 -24146 8407 -24126
rect 8357 -24186 8407 -24146
rect 8467 -24146 8497 -24126
rect 8467 -24186 8517 -24146
rect 8357 -24256 8517 -24186
rect 8357 -24296 8407 -24256
rect 8377 -24316 8407 -24296
rect 8467 -24296 8517 -24256
rect 8467 -24316 8497 -24296
rect 8577 -24346 8637 -24086
rect 8567 -24356 8637 -24346
rect 8237 -24366 8317 -24356
rect 8237 -24426 8247 -24366
rect 8307 -24376 8317 -24366
rect 8557 -24366 8637 -24356
rect 8557 -24376 8567 -24366
rect 8307 -24426 8567 -24376
rect 8627 -24426 8637 -24366
rect 8237 -24436 8637 -24426
rect 8693 -24016 9093 -24006
rect 8693 -24076 8703 -24016
rect 8763 -24066 9023 -24016
rect 8763 -24076 8773 -24066
rect 8693 -24086 8773 -24076
rect 9013 -24076 9023 -24066
rect 9083 -24076 9093 -24016
rect 9013 -24086 9093 -24076
rect 8693 -24356 8753 -24086
rect 8833 -24146 8863 -24126
rect 8813 -24186 8863 -24146
rect 8923 -24146 8953 -24126
rect 8923 -24186 8973 -24146
rect 8813 -24256 8973 -24186
rect 8813 -24296 8863 -24256
rect 8833 -24316 8863 -24296
rect 8923 -24296 8973 -24256
rect 8923 -24316 8953 -24296
rect 9033 -24346 9093 -24086
rect 9023 -24356 9093 -24346
rect 8693 -24366 8773 -24356
rect 8693 -24426 8703 -24366
rect 8763 -24376 8773 -24366
rect 9013 -24366 9093 -24356
rect 9013 -24376 9023 -24366
rect 8763 -24426 9023 -24376
rect 9083 -24426 9093 -24366
rect 8693 -24436 9093 -24426
rect 9151 -24016 9551 -24006
rect 9151 -24076 9161 -24016
rect 9221 -24066 9481 -24016
rect 9221 -24076 9231 -24066
rect 9151 -24086 9231 -24076
rect 9471 -24076 9481 -24066
rect 9541 -24076 9551 -24016
rect 9471 -24086 9551 -24076
rect 9151 -24356 9211 -24086
rect 9291 -24146 9321 -24126
rect 9271 -24186 9321 -24146
rect 9381 -24146 9411 -24126
rect 9381 -24186 9431 -24146
rect 9271 -24256 9431 -24186
rect 9271 -24296 9321 -24256
rect 9291 -24316 9321 -24296
rect 9381 -24296 9431 -24256
rect 9381 -24316 9411 -24296
rect 9491 -24346 9551 -24086
rect 9481 -24356 9551 -24346
rect 9151 -24366 9231 -24356
rect 9151 -24426 9161 -24366
rect 9221 -24376 9231 -24366
rect 9471 -24366 9551 -24356
rect 9471 -24376 9481 -24366
rect 9221 -24426 9481 -24376
rect 9541 -24426 9551 -24366
rect 9151 -24436 9551 -24426
rect 9607 -24016 10007 -24006
rect 9607 -24076 9617 -24016
rect 9677 -24066 9937 -24016
rect 9677 -24076 9687 -24066
rect 9607 -24086 9687 -24076
rect 9927 -24076 9937 -24066
rect 9997 -24076 10007 -24016
rect 9927 -24086 10007 -24076
rect 9607 -24356 9667 -24086
rect 9747 -24146 9777 -24126
rect 9727 -24186 9777 -24146
rect 9837 -24146 9867 -24126
rect 9837 -24186 9887 -24146
rect 9727 -24256 9887 -24186
rect 9727 -24296 9777 -24256
rect 9747 -24316 9777 -24296
rect 9837 -24296 9887 -24256
rect 9837 -24316 9867 -24296
rect 9947 -24346 10007 -24086
rect 9937 -24356 10007 -24346
rect 9607 -24366 9687 -24356
rect 9607 -24426 9617 -24366
rect 9677 -24376 9687 -24366
rect 9927 -24366 10007 -24356
rect 9927 -24376 9937 -24366
rect 9677 -24426 9937 -24376
rect 9997 -24426 10007 -24366
rect 9607 -24436 10007 -24426
rect 10063 -24016 10463 -24006
rect 10063 -24076 10073 -24016
rect 10133 -24066 10393 -24016
rect 10133 -24076 10143 -24066
rect 10063 -24086 10143 -24076
rect 10383 -24076 10393 -24066
rect 10453 -24076 10463 -24016
rect 10383 -24086 10463 -24076
rect 10063 -24356 10123 -24086
rect 10203 -24146 10233 -24126
rect 10183 -24186 10233 -24146
rect 10293 -24146 10323 -24126
rect 10293 -24186 10343 -24146
rect 10183 -24256 10343 -24186
rect 10183 -24296 10233 -24256
rect 10203 -24316 10233 -24296
rect 10293 -24296 10343 -24256
rect 10293 -24316 10323 -24296
rect 10403 -24346 10463 -24086
rect 10393 -24356 10463 -24346
rect 10063 -24366 10143 -24356
rect 10063 -24426 10073 -24366
rect 10133 -24376 10143 -24366
rect 10383 -24366 10463 -24356
rect 10383 -24376 10393 -24366
rect 10133 -24426 10393 -24376
rect 10453 -24426 10463 -24366
rect 10063 -24436 10463 -24426
rect 10521 -24016 10921 -24006
rect 10521 -24076 10531 -24016
rect 10591 -24066 10851 -24016
rect 10591 -24076 10601 -24066
rect 10521 -24086 10601 -24076
rect 10841 -24076 10851 -24066
rect 10911 -24076 10921 -24016
rect 10841 -24086 10921 -24076
rect 10521 -24356 10581 -24086
rect 10661 -24146 10691 -24126
rect 10641 -24186 10691 -24146
rect 10751 -24146 10781 -24126
rect 10751 -24186 10801 -24146
rect 10641 -24256 10801 -24186
rect 10641 -24296 10691 -24256
rect 10661 -24316 10691 -24296
rect 10751 -24296 10801 -24256
rect 10751 -24316 10781 -24296
rect 10861 -24346 10921 -24086
rect 10851 -24356 10921 -24346
rect 10521 -24366 10601 -24356
rect 10521 -24426 10531 -24366
rect 10591 -24376 10601 -24366
rect 10841 -24366 10921 -24356
rect 10841 -24376 10851 -24366
rect 10591 -24426 10851 -24376
rect 10911 -24426 10921 -24366
rect 10521 -24436 10921 -24426
rect 10977 -24016 11377 -24006
rect 10977 -24076 10987 -24016
rect 11047 -24066 11307 -24016
rect 11047 -24076 11057 -24066
rect 10977 -24086 11057 -24076
rect 11297 -24076 11307 -24066
rect 11367 -24076 11377 -24016
rect 11297 -24086 11377 -24076
rect 10977 -24356 11037 -24086
rect 11117 -24146 11147 -24126
rect 11097 -24186 11147 -24146
rect 11207 -24146 11237 -24126
rect 11207 -24186 11257 -24146
rect 11097 -24256 11257 -24186
rect 11097 -24296 11147 -24256
rect 11117 -24316 11147 -24296
rect 11207 -24296 11257 -24256
rect 11207 -24316 11237 -24296
rect 11317 -24346 11377 -24086
rect 11307 -24356 11377 -24346
rect 10977 -24366 11057 -24356
rect 10977 -24426 10987 -24366
rect 11047 -24376 11057 -24366
rect 11297 -24366 11377 -24356
rect 11297 -24376 11307 -24366
rect 11047 -24426 11307 -24376
rect 11367 -24426 11377 -24366
rect 10977 -24436 11377 -24426
rect 11433 -24016 11833 -24006
rect 11433 -24076 11443 -24016
rect 11503 -24066 11763 -24016
rect 11503 -24076 11513 -24066
rect 11433 -24086 11513 -24076
rect 11753 -24076 11763 -24066
rect 11823 -24076 11833 -24016
rect 11753 -24086 11833 -24076
rect 11433 -24356 11493 -24086
rect 11573 -24146 11603 -24126
rect 11553 -24186 11603 -24146
rect 11663 -24146 11693 -24126
rect 11663 -24186 11713 -24146
rect 11553 -24256 11713 -24186
rect 11553 -24296 11603 -24256
rect 11573 -24316 11603 -24296
rect 11663 -24296 11713 -24256
rect 11663 -24316 11693 -24296
rect 11773 -24346 11833 -24086
rect 11763 -24356 11833 -24346
rect 11433 -24366 11513 -24356
rect 11433 -24426 11443 -24366
rect 11503 -24376 11513 -24366
rect 11753 -24366 11833 -24356
rect 11753 -24376 11763 -24366
rect 11503 -24426 11763 -24376
rect 11823 -24426 11833 -24366
rect 11433 -24436 11833 -24426
rect 11891 -24016 12291 -24006
rect 11891 -24076 11901 -24016
rect 11961 -24066 12221 -24016
rect 11961 -24076 11971 -24066
rect 11891 -24086 11971 -24076
rect 12211 -24076 12221 -24066
rect 12281 -24076 12291 -24016
rect 12211 -24086 12291 -24076
rect 11891 -24356 11951 -24086
rect 12031 -24146 12061 -24126
rect 12011 -24186 12061 -24146
rect 12121 -24146 12151 -24126
rect 12121 -24186 12171 -24146
rect 12011 -24256 12171 -24186
rect 12011 -24296 12061 -24256
rect 12031 -24316 12061 -24296
rect 12121 -24296 12171 -24256
rect 12121 -24316 12151 -24296
rect 12231 -24346 12291 -24086
rect 12221 -24356 12291 -24346
rect 11891 -24366 11971 -24356
rect 11891 -24426 11901 -24366
rect 11961 -24376 11971 -24366
rect 12211 -24366 12291 -24356
rect 12211 -24376 12221 -24366
rect 11961 -24426 12221 -24376
rect 12281 -24426 12291 -24366
rect 11891 -24436 12291 -24426
rect 12347 -24016 12747 -24006
rect 12347 -24076 12357 -24016
rect 12417 -24066 12677 -24016
rect 12417 -24076 12427 -24066
rect 12347 -24086 12427 -24076
rect 12667 -24076 12677 -24066
rect 12737 -24076 12747 -24016
rect 12667 -24086 12747 -24076
rect 12347 -24356 12407 -24086
rect 12487 -24146 12517 -24126
rect 12467 -24186 12517 -24146
rect 12577 -24146 12607 -24126
rect 12577 -24186 12627 -24146
rect 12467 -24256 12627 -24186
rect 12467 -24296 12517 -24256
rect 12487 -24316 12517 -24296
rect 12577 -24296 12627 -24256
rect 12577 -24316 12607 -24296
rect 12687 -24346 12747 -24086
rect 12677 -24356 12747 -24346
rect 12347 -24366 12427 -24356
rect 12347 -24426 12357 -24366
rect 12417 -24376 12427 -24366
rect 12667 -24366 12747 -24356
rect 12667 -24376 12677 -24366
rect 12417 -24426 12677 -24376
rect 12737 -24426 12747 -24366
rect 12347 -24436 12747 -24426
rect 12803 -24016 13203 -24006
rect 12803 -24076 12813 -24016
rect 12873 -24066 13133 -24016
rect 12873 -24076 12883 -24066
rect 12803 -24086 12883 -24076
rect 13123 -24076 13133 -24066
rect 13193 -24076 13203 -24016
rect 13123 -24086 13203 -24076
rect 12803 -24356 12863 -24086
rect 12943 -24146 12973 -24126
rect 12923 -24186 12973 -24146
rect 13033 -24146 13063 -24126
rect 13033 -24186 13083 -24146
rect 12923 -24256 13083 -24186
rect 12923 -24296 12973 -24256
rect 12943 -24316 12973 -24296
rect 13033 -24296 13083 -24256
rect 13033 -24316 13063 -24296
rect 13143 -24346 13203 -24086
rect 13133 -24356 13203 -24346
rect 12803 -24366 12883 -24356
rect 12803 -24426 12813 -24366
rect 12873 -24376 12883 -24366
rect 13123 -24366 13203 -24356
rect 13123 -24376 13133 -24366
rect 12873 -24426 13133 -24376
rect 13193 -24426 13203 -24366
rect 12803 -24436 13203 -24426
rect 13261 -24016 13661 -24006
rect 13261 -24076 13271 -24016
rect 13331 -24066 13591 -24016
rect 13331 -24076 13341 -24066
rect 13261 -24086 13341 -24076
rect 13581 -24076 13591 -24066
rect 13651 -24076 13661 -24016
rect 13581 -24086 13661 -24076
rect 13261 -24356 13321 -24086
rect 13401 -24146 13431 -24126
rect 13381 -24186 13431 -24146
rect 13491 -24146 13521 -24126
rect 13491 -24186 13541 -24146
rect 13381 -24256 13541 -24186
rect 13381 -24296 13431 -24256
rect 13401 -24316 13431 -24296
rect 13491 -24296 13541 -24256
rect 13491 -24316 13521 -24296
rect 13601 -24346 13661 -24086
rect 13591 -24356 13661 -24346
rect 13261 -24366 13341 -24356
rect 13261 -24426 13271 -24366
rect 13331 -24376 13341 -24366
rect 13581 -24366 13661 -24356
rect 13581 -24376 13591 -24366
rect 13331 -24426 13591 -24376
rect 13651 -24426 13661 -24366
rect 13261 -24436 13661 -24426
rect 13717 -24016 14117 -24006
rect 13717 -24076 13727 -24016
rect 13787 -24066 14047 -24016
rect 13787 -24076 13797 -24066
rect 13717 -24086 13797 -24076
rect 14037 -24076 14047 -24066
rect 14107 -24076 14117 -24016
rect 14037 -24086 14117 -24076
rect 13717 -24356 13777 -24086
rect 13857 -24146 13887 -24126
rect 13837 -24186 13887 -24146
rect 13947 -24146 13977 -24126
rect 13947 -24186 13997 -24146
rect 13837 -24256 13997 -24186
rect 13837 -24296 13887 -24256
rect 13857 -24316 13887 -24296
rect 13947 -24296 13997 -24256
rect 13947 -24316 13977 -24296
rect 14057 -24346 14117 -24086
rect 14047 -24356 14117 -24346
rect 13717 -24366 13797 -24356
rect 13717 -24426 13727 -24366
rect 13787 -24376 13797 -24366
rect 14037 -24366 14117 -24356
rect 14037 -24376 14047 -24366
rect 13787 -24426 14047 -24376
rect 14107 -24426 14117 -24366
rect 13717 -24436 14117 -24426
rect 14173 -24016 14573 -24006
rect 14173 -24076 14183 -24016
rect 14243 -24066 14503 -24016
rect 14243 -24076 14253 -24066
rect 14173 -24086 14253 -24076
rect 14493 -24076 14503 -24066
rect 14563 -24076 14573 -24016
rect 14493 -24086 14573 -24076
rect 14173 -24356 14233 -24086
rect 14313 -24146 14343 -24126
rect 14293 -24186 14343 -24146
rect 14403 -24146 14433 -24126
rect 14403 -24186 14453 -24146
rect 14293 -24256 14453 -24186
rect 14293 -24296 14343 -24256
rect 14313 -24316 14343 -24296
rect 14403 -24296 14453 -24256
rect 14403 -24316 14433 -24296
rect 14513 -24346 14573 -24086
rect 14503 -24356 14573 -24346
rect 14173 -24366 14253 -24356
rect 14173 -24426 14183 -24366
rect 14243 -24376 14253 -24366
rect 14493 -24366 14573 -24356
rect 14493 -24376 14503 -24366
rect 14243 -24426 14503 -24376
rect 14563 -24426 14573 -24366
rect 14173 -24436 14573 -24426
rect 14631 -24016 15031 -24006
rect 14631 -24076 14641 -24016
rect 14701 -24066 14961 -24016
rect 14701 -24076 14711 -24066
rect 14631 -24086 14711 -24076
rect 14951 -24076 14961 -24066
rect 15021 -24076 15031 -24016
rect 14951 -24086 15031 -24076
rect 14631 -24356 14691 -24086
rect 14771 -24146 14801 -24126
rect 14751 -24186 14801 -24146
rect 14861 -24146 14891 -24126
rect 14861 -24186 14911 -24146
rect 14751 -24256 14911 -24186
rect 14751 -24296 14801 -24256
rect 14771 -24316 14801 -24296
rect 14861 -24296 14911 -24256
rect 14861 -24316 14891 -24296
rect 14971 -24346 15031 -24086
rect 14961 -24356 15031 -24346
rect 14631 -24366 14711 -24356
rect 14631 -24426 14641 -24366
rect 14701 -24376 14711 -24366
rect 14951 -24366 15031 -24356
rect 14951 -24376 14961 -24366
rect 14701 -24426 14961 -24376
rect 15021 -24426 15031 -24366
rect 14631 -24436 15031 -24426
rect 15087 -24016 15487 -24006
rect 15087 -24076 15097 -24016
rect 15157 -24066 15417 -24016
rect 15157 -24076 15167 -24066
rect 15087 -24086 15167 -24076
rect 15407 -24076 15417 -24066
rect 15477 -24076 15487 -24016
rect 15407 -24086 15487 -24076
rect 15087 -24356 15147 -24086
rect 15227 -24146 15257 -24126
rect 15207 -24186 15257 -24146
rect 15317 -24146 15347 -24126
rect 15317 -24186 15367 -24146
rect 15207 -24256 15367 -24186
rect 15207 -24296 15257 -24256
rect 15227 -24316 15257 -24296
rect 15317 -24296 15367 -24256
rect 15317 -24316 15347 -24296
rect 15427 -24346 15487 -24086
rect 15417 -24356 15487 -24346
rect 15087 -24366 15167 -24356
rect 15087 -24426 15097 -24366
rect 15157 -24376 15167 -24366
rect 15407 -24366 15487 -24356
rect 15407 -24376 15417 -24366
rect 15157 -24426 15417 -24376
rect 15477 -24426 15487 -24366
rect 15087 -24436 15487 -24426
rect 1 -24518 401 -24508
rect 1 -24578 11 -24518
rect 71 -24568 331 -24518
rect 71 -24578 81 -24568
rect 1 -24588 81 -24578
rect 321 -24578 331 -24568
rect 391 -24578 401 -24518
rect 321 -24588 401 -24578
rect 1 -24858 61 -24588
rect 141 -24648 171 -24628
rect 121 -24688 171 -24648
rect 231 -24648 261 -24628
rect 231 -24688 281 -24648
rect 121 -24758 281 -24688
rect 121 -24798 171 -24758
rect 141 -24818 171 -24798
rect 231 -24798 281 -24758
rect 231 -24818 261 -24798
rect 341 -24848 401 -24588
rect 331 -24858 401 -24848
rect 1 -24868 81 -24858
rect 1 -24928 11 -24868
rect 71 -24878 81 -24868
rect 321 -24868 401 -24858
rect 321 -24878 331 -24868
rect 71 -24928 331 -24878
rect 391 -24928 401 -24868
rect 1 -24938 401 -24928
rect 457 -24518 857 -24508
rect 457 -24578 467 -24518
rect 527 -24568 787 -24518
rect 527 -24578 537 -24568
rect 457 -24588 537 -24578
rect 777 -24578 787 -24568
rect 847 -24578 857 -24518
rect 777 -24588 857 -24578
rect 457 -24858 517 -24588
rect 597 -24648 627 -24628
rect 577 -24688 627 -24648
rect 687 -24648 717 -24628
rect 687 -24688 737 -24648
rect 577 -24758 737 -24688
rect 577 -24798 627 -24758
rect 597 -24818 627 -24798
rect 687 -24798 737 -24758
rect 687 -24818 717 -24798
rect 797 -24848 857 -24588
rect 787 -24858 857 -24848
rect 457 -24868 537 -24858
rect 457 -24928 467 -24868
rect 527 -24878 537 -24868
rect 777 -24868 857 -24858
rect 777 -24878 787 -24868
rect 527 -24928 787 -24878
rect 847 -24928 857 -24868
rect 457 -24938 857 -24928
rect 913 -24518 1313 -24508
rect 913 -24578 923 -24518
rect 983 -24568 1243 -24518
rect 983 -24578 993 -24568
rect 913 -24588 993 -24578
rect 1233 -24578 1243 -24568
rect 1303 -24578 1313 -24518
rect 1233 -24588 1313 -24578
rect 913 -24858 973 -24588
rect 1053 -24648 1083 -24628
rect 1033 -24688 1083 -24648
rect 1143 -24648 1173 -24628
rect 1143 -24688 1193 -24648
rect 1033 -24758 1193 -24688
rect 1033 -24798 1083 -24758
rect 1053 -24818 1083 -24798
rect 1143 -24798 1193 -24758
rect 1143 -24818 1173 -24798
rect 1253 -24848 1313 -24588
rect 1243 -24858 1313 -24848
rect 913 -24868 993 -24858
rect 913 -24928 923 -24868
rect 983 -24878 993 -24868
rect 1233 -24868 1313 -24858
rect 1233 -24878 1243 -24868
rect 983 -24928 1243 -24878
rect 1303 -24928 1313 -24868
rect 913 -24938 1313 -24928
rect 1371 -24518 1771 -24508
rect 1371 -24578 1381 -24518
rect 1441 -24568 1701 -24518
rect 1441 -24578 1451 -24568
rect 1371 -24588 1451 -24578
rect 1691 -24578 1701 -24568
rect 1761 -24578 1771 -24518
rect 1691 -24588 1771 -24578
rect 1371 -24858 1431 -24588
rect 1511 -24648 1541 -24628
rect 1491 -24688 1541 -24648
rect 1601 -24648 1631 -24628
rect 1601 -24688 1651 -24648
rect 1491 -24758 1651 -24688
rect 1491 -24798 1541 -24758
rect 1511 -24818 1541 -24798
rect 1601 -24798 1651 -24758
rect 1601 -24818 1631 -24798
rect 1711 -24848 1771 -24588
rect 1701 -24858 1771 -24848
rect 1371 -24868 1451 -24858
rect 1371 -24928 1381 -24868
rect 1441 -24878 1451 -24868
rect 1691 -24868 1771 -24858
rect 1691 -24878 1701 -24868
rect 1441 -24928 1701 -24878
rect 1761 -24928 1771 -24868
rect 1371 -24938 1771 -24928
rect 1827 -24518 2227 -24508
rect 1827 -24578 1837 -24518
rect 1897 -24568 2157 -24518
rect 1897 -24578 1907 -24568
rect 1827 -24588 1907 -24578
rect 2147 -24578 2157 -24568
rect 2217 -24578 2227 -24518
rect 2147 -24588 2227 -24578
rect 1827 -24858 1887 -24588
rect 1967 -24648 1997 -24628
rect 1947 -24688 1997 -24648
rect 2057 -24648 2087 -24628
rect 2057 -24688 2107 -24648
rect 1947 -24758 2107 -24688
rect 1947 -24798 1997 -24758
rect 1967 -24818 1997 -24798
rect 2057 -24798 2107 -24758
rect 2057 -24818 2087 -24798
rect 2167 -24848 2227 -24588
rect 2157 -24858 2227 -24848
rect 1827 -24868 1907 -24858
rect 1827 -24928 1837 -24868
rect 1897 -24878 1907 -24868
rect 2147 -24868 2227 -24858
rect 2147 -24878 2157 -24868
rect 1897 -24928 2157 -24878
rect 2217 -24928 2227 -24868
rect 1827 -24938 2227 -24928
rect 2283 -24518 2683 -24508
rect 2283 -24578 2293 -24518
rect 2353 -24568 2613 -24518
rect 2353 -24578 2363 -24568
rect 2283 -24588 2363 -24578
rect 2603 -24578 2613 -24568
rect 2673 -24578 2683 -24518
rect 2603 -24588 2683 -24578
rect 2283 -24858 2343 -24588
rect 2423 -24648 2453 -24628
rect 2403 -24688 2453 -24648
rect 2513 -24648 2543 -24628
rect 2513 -24688 2563 -24648
rect 2403 -24758 2563 -24688
rect 2403 -24798 2453 -24758
rect 2423 -24818 2453 -24798
rect 2513 -24798 2563 -24758
rect 2513 -24818 2543 -24798
rect 2623 -24848 2683 -24588
rect 2613 -24858 2683 -24848
rect 2283 -24868 2363 -24858
rect 2283 -24928 2293 -24868
rect 2353 -24878 2363 -24868
rect 2603 -24868 2683 -24858
rect 2603 -24878 2613 -24868
rect 2353 -24928 2613 -24878
rect 2673 -24928 2683 -24868
rect 2283 -24938 2683 -24928
rect 2741 -24518 3141 -24508
rect 2741 -24578 2751 -24518
rect 2811 -24568 3071 -24518
rect 2811 -24578 2821 -24568
rect 2741 -24588 2821 -24578
rect 3061 -24578 3071 -24568
rect 3131 -24578 3141 -24518
rect 3061 -24588 3141 -24578
rect 2741 -24858 2801 -24588
rect 2881 -24648 2911 -24628
rect 2861 -24688 2911 -24648
rect 2971 -24648 3001 -24628
rect 2971 -24688 3021 -24648
rect 2861 -24758 3021 -24688
rect 2861 -24798 2911 -24758
rect 2881 -24818 2911 -24798
rect 2971 -24798 3021 -24758
rect 2971 -24818 3001 -24798
rect 3081 -24848 3141 -24588
rect 3071 -24858 3141 -24848
rect 2741 -24868 2821 -24858
rect 2741 -24928 2751 -24868
rect 2811 -24878 2821 -24868
rect 3061 -24868 3141 -24858
rect 3061 -24878 3071 -24868
rect 2811 -24928 3071 -24878
rect 3131 -24928 3141 -24868
rect 2741 -24938 3141 -24928
rect 3197 -24518 3597 -24508
rect 3197 -24578 3207 -24518
rect 3267 -24568 3527 -24518
rect 3267 -24578 3277 -24568
rect 3197 -24588 3277 -24578
rect 3517 -24578 3527 -24568
rect 3587 -24578 3597 -24518
rect 3517 -24588 3597 -24578
rect 3197 -24858 3257 -24588
rect 3337 -24648 3367 -24628
rect 3317 -24688 3367 -24648
rect 3427 -24648 3457 -24628
rect 3427 -24688 3477 -24648
rect 3317 -24758 3477 -24688
rect 3317 -24798 3367 -24758
rect 3337 -24818 3367 -24798
rect 3427 -24798 3477 -24758
rect 3427 -24818 3457 -24798
rect 3537 -24848 3597 -24588
rect 3527 -24858 3597 -24848
rect 3197 -24868 3277 -24858
rect 3197 -24928 3207 -24868
rect 3267 -24878 3277 -24868
rect 3517 -24868 3597 -24858
rect 3517 -24878 3527 -24868
rect 3267 -24928 3527 -24878
rect 3587 -24928 3597 -24868
rect 3197 -24938 3597 -24928
rect 3653 -24518 4053 -24508
rect 3653 -24578 3663 -24518
rect 3723 -24568 3983 -24518
rect 3723 -24578 3733 -24568
rect 3653 -24588 3733 -24578
rect 3973 -24578 3983 -24568
rect 4043 -24578 4053 -24518
rect 3973 -24588 4053 -24578
rect 3653 -24858 3713 -24588
rect 3793 -24648 3823 -24628
rect 3773 -24688 3823 -24648
rect 3883 -24648 3913 -24628
rect 3883 -24688 3933 -24648
rect 3773 -24758 3933 -24688
rect 3773 -24798 3823 -24758
rect 3793 -24818 3823 -24798
rect 3883 -24798 3933 -24758
rect 3883 -24818 3913 -24798
rect 3993 -24848 4053 -24588
rect 3983 -24858 4053 -24848
rect 3653 -24868 3733 -24858
rect 3653 -24928 3663 -24868
rect 3723 -24878 3733 -24868
rect 3973 -24868 4053 -24858
rect 3973 -24878 3983 -24868
rect 3723 -24928 3983 -24878
rect 4043 -24928 4053 -24868
rect 3653 -24938 4053 -24928
rect 4111 -24518 4511 -24508
rect 4111 -24578 4121 -24518
rect 4181 -24568 4441 -24518
rect 4181 -24578 4191 -24568
rect 4111 -24588 4191 -24578
rect 4431 -24578 4441 -24568
rect 4501 -24578 4511 -24518
rect 4431 -24588 4511 -24578
rect 4111 -24858 4171 -24588
rect 4251 -24648 4281 -24628
rect 4231 -24688 4281 -24648
rect 4341 -24648 4371 -24628
rect 4341 -24688 4391 -24648
rect 4231 -24758 4391 -24688
rect 4231 -24798 4281 -24758
rect 4251 -24818 4281 -24798
rect 4341 -24798 4391 -24758
rect 4341 -24818 4371 -24798
rect 4451 -24848 4511 -24588
rect 4441 -24858 4511 -24848
rect 4111 -24868 4191 -24858
rect 4111 -24928 4121 -24868
rect 4181 -24878 4191 -24868
rect 4431 -24868 4511 -24858
rect 4431 -24878 4441 -24868
rect 4181 -24928 4441 -24878
rect 4501 -24928 4511 -24868
rect 4111 -24938 4511 -24928
rect 4567 -24518 4967 -24508
rect 4567 -24578 4577 -24518
rect 4637 -24568 4897 -24518
rect 4637 -24578 4647 -24568
rect 4567 -24588 4647 -24578
rect 4887 -24578 4897 -24568
rect 4957 -24578 4967 -24518
rect 4887 -24588 4967 -24578
rect 4567 -24858 4627 -24588
rect 4707 -24648 4737 -24628
rect 4687 -24688 4737 -24648
rect 4797 -24648 4827 -24628
rect 4797 -24688 4847 -24648
rect 4687 -24758 4847 -24688
rect 4687 -24798 4737 -24758
rect 4707 -24818 4737 -24798
rect 4797 -24798 4847 -24758
rect 4797 -24818 4827 -24798
rect 4907 -24848 4967 -24588
rect 4897 -24858 4967 -24848
rect 4567 -24868 4647 -24858
rect 4567 -24928 4577 -24868
rect 4637 -24878 4647 -24868
rect 4887 -24868 4967 -24858
rect 4887 -24878 4897 -24868
rect 4637 -24928 4897 -24878
rect 4957 -24928 4967 -24868
rect 4567 -24938 4967 -24928
rect 5023 -24518 5423 -24508
rect 5023 -24578 5033 -24518
rect 5093 -24568 5353 -24518
rect 5093 -24578 5103 -24568
rect 5023 -24588 5103 -24578
rect 5343 -24578 5353 -24568
rect 5413 -24578 5423 -24518
rect 5343 -24588 5423 -24578
rect 5023 -24858 5083 -24588
rect 5163 -24648 5193 -24628
rect 5143 -24688 5193 -24648
rect 5253 -24648 5283 -24628
rect 5253 -24688 5303 -24648
rect 5143 -24758 5303 -24688
rect 5143 -24798 5193 -24758
rect 5163 -24818 5193 -24798
rect 5253 -24798 5303 -24758
rect 5253 -24818 5283 -24798
rect 5363 -24848 5423 -24588
rect 5353 -24858 5423 -24848
rect 5023 -24868 5103 -24858
rect 5023 -24928 5033 -24868
rect 5093 -24878 5103 -24868
rect 5343 -24868 5423 -24858
rect 5343 -24878 5353 -24868
rect 5093 -24928 5353 -24878
rect 5413 -24928 5423 -24868
rect 5023 -24938 5423 -24928
rect 5481 -24518 5881 -24508
rect 5481 -24578 5491 -24518
rect 5551 -24568 5811 -24518
rect 5551 -24578 5561 -24568
rect 5481 -24588 5561 -24578
rect 5801 -24578 5811 -24568
rect 5871 -24578 5881 -24518
rect 5801 -24588 5881 -24578
rect 5481 -24858 5541 -24588
rect 5621 -24648 5651 -24628
rect 5601 -24688 5651 -24648
rect 5711 -24648 5741 -24628
rect 5711 -24688 5761 -24648
rect 5601 -24758 5761 -24688
rect 5601 -24798 5651 -24758
rect 5621 -24818 5651 -24798
rect 5711 -24798 5761 -24758
rect 5711 -24818 5741 -24798
rect 5821 -24848 5881 -24588
rect 5811 -24858 5881 -24848
rect 5481 -24868 5561 -24858
rect 5481 -24928 5491 -24868
rect 5551 -24878 5561 -24868
rect 5801 -24868 5881 -24858
rect 5801 -24878 5811 -24868
rect 5551 -24928 5811 -24878
rect 5871 -24928 5881 -24868
rect 5481 -24938 5881 -24928
rect 5937 -24518 6337 -24508
rect 5937 -24578 5947 -24518
rect 6007 -24568 6267 -24518
rect 6007 -24578 6017 -24568
rect 5937 -24588 6017 -24578
rect 6257 -24578 6267 -24568
rect 6327 -24578 6337 -24518
rect 6257 -24588 6337 -24578
rect 5937 -24858 5997 -24588
rect 6077 -24648 6107 -24628
rect 6057 -24688 6107 -24648
rect 6167 -24648 6197 -24628
rect 6167 -24688 6217 -24648
rect 6057 -24758 6217 -24688
rect 6057 -24798 6107 -24758
rect 6077 -24818 6107 -24798
rect 6167 -24798 6217 -24758
rect 6167 -24818 6197 -24798
rect 6277 -24848 6337 -24588
rect 6267 -24858 6337 -24848
rect 5937 -24868 6017 -24858
rect 5937 -24928 5947 -24868
rect 6007 -24878 6017 -24868
rect 6257 -24868 6337 -24858
rect 6257 -24878 6267 -24868
rect 6007 -24928 6267 -24878
rect 6327 -24928 6337 -24868
rect 5937 -24938 6337 -24928
rect 6393 -24518 6793 -24508
rect 6393 -24578 6403 -24518
rect 6463 -24568 6723 -24518
rect 6463 -24578 6473 -24568
rect 6393 -24588 6473 -24578
rect 6713 -24578 6723 -24568
rect 6783 -24578 6793 -24518
rect 6713 -24588 6793 -24578
rect 6393 -24858 6453 -24588
rect 6533 -24648 6563 -24628
rect 6513 -24688 6563 -24648
rect 6623 -24648 6653 -24628
rect 6623 -24688 6673 -24648
rect 6513 -24758 6673 -24688
rect 6513 -24798 6563 -24758
rect 6533 -24818 6563 -24798
rect 6623 -24798 6673 -24758
rect 6623 -24818 6653 -24798
rect 6733 -24848 6793 -24588
rect 6723 -24858 6793 -24848
rect 6393 -24868 6473 -24858
rect 6393 -24928 6403 -24868
rect 6463 -24878 6473 -24868
rect 6713 -24868 6793 -24858
rect 6713 -24878 6723 -24868
rect 6463 -24928 6723 -24878
rect 6783 -24928 6793 -24868
rect 6393 -24938 6793 -24928
rect 6851 -24518 7251 -24508
rect 6851 -24578 6861 -24518
rect 6921 -24568 7181 -24518
rect 6921 -24578 6931 -24568
rect 6851 -24588 6931 -24578
rect 7171 -24578 7181 -24568
rect 7241 -24578 7251 -24518
rect 7171 -24588 7251 -24578
rect 6851 -24858 6911 -24588
rect 6991 -24648 7021 -24628
rect 6971 -24688 7021 -24648
rect 7081 -24648 7111 -24628
rect 7081 -24688 7131 -24648
rect 6971 -24758 7131 -24688
rect 6971 -24798 7021 -24758
rect 6991 -24818 7021 -24798
rect 7081 -24798 7131 -24758
rect 7081 -24818 7111 -24798
rect 7191 -24848 7251 -24588
rect 7181 -24858 7251 -24848
rect 6851 -24868 6931 -24858
rect 6851 -24928 6861 -24868
rect 6921 -24878 6931 -24868
rect 7171 -24868 7251 -24858
rect 7171 -24878 7181 -24868
rect 6921 -24928 7181 -24878
rect 7241 -24928 7251 -24868
rect 6851 -24938 7251 -24928
rect 7307 -24518 7707 -24508
rect 7307 -24578 7317 -24518
rect 7377 -24568 7637 -24518
rect 7377 -24578 7387 -24568
rect 7307 -24588 7387 -24578
rect 7627 -24578 7637 -24568
rect 7697 -24578 7707 -24518
rect 7627 -24588 7707 -24578
rect 7307 -24858 7367 -24588
rect 7447 -24648 7477 -24628
rect 7427 -24688 7477 -24648
rect 7537 -24648 7567 -24628
rect 7537 -24688 7587 -24648
rect 7427 -24758 7587 -24688
rect 7427 -24798 7477 -24758
rect 7447 -24818 7477 -24798
rect 7537 -24798 7587 -24758
rect 7537 -24818 7567 -24798
rect 7647 -24848 7707 -24588
rect 7637 -24858 7707 -24848
rect 7307 -24868 7387 -24858
rect 7307 -24928 7317 -24868
rect 7377 -24878 7387 -24868
rect 7627 -24868 7707 -24858
rect 7627 -24878 7637 -24868
rect 7377 -24928 7637 -24878
rect 7697 -24928 7707 -24868
rect 7307 -24938 7707 -24928
rect 7763 -24518 8163 -24508
rect 7763 -24578 7773 -24518
rect 7833 -24568 8093 -24518
rect 7833 -24578 7843 -24568
rect 7763 -24588 7843 -24578
rect 8083 -24578 8093 -24568
rect 8153 -24578 8163 -24518
rect 8083 -24588 8163 -24578
rect 7763 -24858 7823 -24588
rect 7903 -24648 7933 -24628
rect 7883 -24688 7933 -24648
rect 7993 -24648 8023 -24628
rect 7993 -24688 8043 -24648
rect 7883 -24758 8043 -24688
rect 7883 -24798 7933 -24758
rect 7903 -24818 7933 -24798
rect 7993 -24798 8043 -24758
rect 7993 -24818 8023 -24798
rect 8103 -24848 8163 -24588
rect 8093 -24858 8163 -24848
rect 7763 -24868 7843 -24858
rect 7763 -24928 7773 -24868
rect 7833 -24878 7843 -24868
rect 8083 -24868 8163 -24858
rect 8083 -24878 8093 -24868
rect 7833 -24928 8093 -24878
rect 8153 -24928 8163 -24868
rect 7763 -24938 8163 -24928
rect 8237 -24518 8637 -24508
rect 8237 -24578 8247 -24518
rect 8307 -24568 8567 -24518
rect 8307 -24578 8317 -24568
rect 8237 -24588 8317 -24578
rect 8557 -24578 8567 -24568
rect 8627 -24578 8637 -24518
rect 8557 -24588 8637 -24578
rect 8237 -24858 8297 -24588
rect 8377 -24648 8407 -24628
rect 8357 -24688 8407 -24648
rect 8467 -24648 8497 -24628
rect 8467 -24688 8517 -24648
rect 8357 -24758 8517 -24688
rect 8357 -24798 8407 -24758
rect 8377 -24818 8407 -24798
rect 8467 -24798 8517 -24758
rect 8467 -24818 8497 -24798
rect 8577 -24848 8637 -24588
rect 8567 -24858 8637 -24848
rect 8237 -24868 8317 -24858
rect 8237 -24928 8247 -24868
rect 8307 -24878 8317 -24868
rect 8557 -24868 8637 -24858
rect 8557 -24878 8567 -24868
rect 8307 -24928 8567 -24878
rect 8627 -24928 8637 -24868
rect 8237 -24938 8637 -24928
rect 8693 -24518 9093 -24508
rect 8693 -24578 8703 -24518
rect 8763 -24568 9023 -24518
rect 8763 -24578 8773 -24568
rect 8693 -24588 8773 -24578
rect 9013 -24578 9023 -24568
rect 9083 -24578 9093 -24518
rect 9013 -24588 9093 -24578
rect 8693 -24858 8753 -24588
rect 8833 -24648 8863 -24628
rect 8813 -24688 8863 -24648
rect 8923 -24648 8953 -24628
rect 8923 -24688 8973 -24648
rect 8813 -24758 8973 -24688
rect 8813 -24798 8863 -24758
rect 8833 -24818 8863 -24798
rect 8923 -24798 8973 -24758
rect 8923 -24818 8953 -24798
rect 9033 -24848 9093 -24588
rect 9023 -24858 9093 -24848
rect 8693 -24868 8773 -24858
rect 8693 -24928 8703 -24868
rect 8763 -24878 8773 -24868
rect 9013 -24868 9093 -24858
rect 9013 -24878 9023 -24868
rect 8763 -24928 9023 -24878
rect 9083 -24928 9093 -24868
rect 8693 -24938 9093 -24928
rect 9151 -24518 9551 -24508
rect 9151 -24578 9161 -24518
rect 9221 -24568 9481 -24518
rect 9221 -24578 9231 -24568
rect 9151 -24588 9231 -24578
rect 9471 -24578 9481 -24568
rect 9541 -24578 9551 -24518
rect 9471 -24588 9551 -24578
rect 9151 -24858 9211 -24588
rect 9291 -24648 9321 -24628
rect 9271 -24688 9321 -24648
rect 9381 -24648 9411 -24628
rect 9381 -24688 9431 -24648
rect 9271 -24758 9431 -24688
rect 9271 -24798 9321 -24758
rect 9291 -24818 9321 -24798
rect 9381 -24798 9431 -24758
rect 9381 -24818 9411 -24798
rect 9491 -24848 9551 -24588
rect 9481 -24858 9551 -24848
rect 9151 -24868 9231 -24858
rect 9151 -24928 9161 -24868
rect 9221 -24878 9231 -24868
rect 9471 -24868 9551 -24858
rect 9471 -24878 9481 -24868
rect 9221 -24928 9481 -24878
rect 9541 -24928 9551 -24868
rect 9151 -24938 9551 -24928
rect 9607 -24518 10007 -24508
rect 9607 -24578 9617 -24518
rect 9677 -24568 9937 -24518
rect 9677 -24578 9687 -24568
rect 9607 -24588 9687 -24578
rect 9927 -24578 9937 -24568
rect 9997 -24578 10007 -24518
rect 9927 -24588 10007 -24578
rect 9607 -24858 9667 -24588
rect 9747 -24648 9777 -24628
rect 9727 -24688 9777 -24648
rect 9837 -24648 9867 -24628
rect 9837 -24688 9887 -24648
rect 9727 -24758 9887 -24688
rect 9727 -24798 9777 -24758
rect 9747 -24818 9777 -24798
rect 9837 -24798 9887 -24758
rect 9837 -24818 9867 -24798
rect 9947 -24848 10007 -24588
rect 9937 -24858 10007 -24848
rect 9607 -24868 9687 -24858
rect 9607 -24928 9617 -24868
rect 9677 -24878 9687 -24868
rect 9927 -24868 10007 -24858
rect 9927 -24878 9937 -24868
rect 9677 -24928 9937 -24878
rect 9997 -24928 10007 -24868
rect 9607 -24938 10007 -24928
rect 10063 -24518 10463 -24508
rect 10063 -24578 10073 -24518
rect 10133 -24568 10393 -24518
rect 10133 -24578 10143 -24568
rect 10063 -24588 10143 -24578
rect 10383 -24578 10393 -24568
rect 10453 -24578 10463 -24518
rect 10383 -24588 10463 -24578
rect 10063 -24858 10123 -24588
rect 10203 -24648 10233 -24628
rect 10183 -24688 10233 -24648
rect 10293 -24648 10323 -24628
rect 10293 -24688 10343 -24648
rect 10183 -24758 10343 -24688
rect 10183 -24798 10233 -24758
rect 10203 -24818 10233 -24798
rect 10293 -24798 10343 -24758
rect 10293 -24818 10323 -24798
rect 10403 -24848 10463 -24588
rect 10393 -24858 10463 -24848
rect 10063 -24868 10143 -24858
rect 10063 -24928 10073 -24868
rect 10133 -24878 10143 -24868
rect 10383 -24868 10463 -24858
rect 10383 -24878 10393 -24868
rect 10133 -24928 10393 -24878
rect 10453 -24928 10463 -24868
rect 10063 -24938 10463 -24928
rect 10521 -24518 10921 -24508
rect 10521 -24578 10531 -24518
rect 10591 -24568 10851 -24518
rect 10591 -24578 10601 -24568
rect 10521 -24588 10601 -24578
rect 10841 -24578 10851 -24568
rect 10911 -24578 10921 -24518
rect 10841 -24588 10921 -24578
rect 10521 -24858 10581 -24588
rect 10661 -24648 10691 -24628
rect 10641 -24688 10691 -24648
rect 10751 -24648 10781 -24628
rect 10751 -24688 10801 -24648
rect 10641 -24758 10801 -24688
rect 10641 -24798 10691 -24758
rect 10661 -24818 10691 -24798
rect 10751 -24798 10801 -24758
rect 10751 -24818 10781 -24798
rect 10861 -24848 10921 -24588
rect 10851 -24858 10921 -24848
rect 10521 -24868 10601 -24858
rect 10521 -24928 10531 -24868
rect 10591 -24878 10601 -24868
rect 10841 -24868 10921 -24858
rect 10841 -24878 10851 -24868
rect 10591 -24928 10851 -24878
rect 10911 -24928 10921 -24868
rect 10521 -24938 10921 -24928
rect 10977 -24518 11377 -24508
rect 10977 -24578 10987 -24518
rect 11047 -24568 11307 -24518
rect 11047 -24578 11057 -24568
rect 10977 -24588 11057 -24578
rect 11297 -24578 11307 -24568
rect 11367 -24578 11377 -24518
rect 11297 -24588 11377 -24578
rect 10977 -24858 11037 -24588
rect 11117 -24648 11147 -24628
rect 11097 -24688 11147 -24648
rect 11207 -24648 11237 -24628
rect 11207 -24688 11257 -24648
rect 11097 -24758 11257 -24688
rect 11097 -24798 11147 -24758
rect 11117 -24818 11147 -24798
rect 11207 -24798 11257 -24758
rect 11207 -24818 11237 -24798
rect 11317 -24848 11377 -24588
rect 11307 -24858 11377 -24848
rect 10977 -24868 11057 -24858
rect 10977 -24928 10987 -24868
rect 11047 -24878 11057 -24868
rect 11297 -24868 11377 -24858
rect 11297 -24878 11307 -24868
rect 11047 -24928 11307 -24878
rect 11367 -24928 11377 -24868
rect 10977 -24938 11377 -24928
rect 11433 -24518 11833 -24508
rect 11433 -24578 11443 -24518
rect 11503 -24568 11763 -24518
rect 11503 -24578 11513 -24568
rect 11433 -24588 11513 -24578
rect 11753 -24578 11763 -24568
rect 11823 -24578 11833 -24518
rect 11753 -24588 11833 -24578
rect 11433 -24858 11493 -24588
rect 11573 -24648 11603 -24628
rect 11553 -24688 11603 -24648
rect 11663 -24648 11693 -24628
rect 11663 -24688 11713 -24648
rect 11553 -24758 11713 -24688
rect 11553 -24798 11603 -24758
rect 11573 -24818 11603 -24798
rect 11663 -24798 11713 -24758
rect 11663 -24818 11693 -24798
rect 11773 -24848 11833 -24588
rect 11763 -24858 11833 -24848
rect 11433 -24868 11513 -24858
rect 11433 -24928 11443 -24868
rect 11503 -24878 11513 -24868
rect 11753 -24868 11833 -24858
rect 11753 -24878 11763 -24868
rect 11503 -24928 11763 -24878
rect 11823 -24928 11833 -24868
rect 11433 -24938 11833 -24928
rect 11891 -24518 12291 -24508
rect 11891 -24578 11901 -24518
rect 11961 -24568 12221 -24518
rect 11961 -24578 11971 -24568
rect 11891 -24588 11971 -24578
rect 12211 -24578 12221 -24568
rect 12281 -24578 12291 -24518
rect 12211 -24588 12291 -24578
rect 11891 -24858 11951 -24588
rect 12031 -24648 12061 -24628
rect 12011 -24688 12061 -24648
rect 12121 -24648 12151 -24628
rect 12121 -24688 12171 -24648
rect 12011 -24758 12171 -24688
rect 12011 -24798 12061 -24758
rect 12031 -24818 12061 -24798
rect 12121 -24798 12171 -24758
rect 12121 -24818 12151 -24798
rect 12231 -24848 12291 -24588
rect 12221 -24858 12291 -24848
rect 11891 -24868 11971 -24858
rect 11891 -24928 11901 -24868
rect 11961 -24878 11971 -24868
rect 12211 -24868 12291 -24858
rect 12211 -24878 12221 -24868
rect 11961 -24928 12221 -24878
rect 12281 -24928 12291 -24868
rect 11891 -24938 12291 -24928
rect 12347 -24518 12747 -24508
rect 12347 -24578 12357 -24518
rect 12417 -24568 12677 -24518
rect 12417 -24578 12427 -24568
rect 12347 -24588 12427 -24578
rect 12667 -24578 12677 -24568
rect 12737 -24578 12747 -24518
rect 12667 -24588 12747 -24578
rect 12347 -24858 12407 -24588
rect 12487 -24648 12517 -24628
rect 12467 -24688 12517 -24648
rect 12577 -24648 12607 -24628
rect 12577 -24688 12627 -24648
rect 12467 -24758 12627 -24688
rect 12467 -24798 12517 -24758
rect 12487 -24818 12517 -24798
rect 12577 -24798 12627 -24758
rect 12577 -24818 12607 -24798
rect 12687 -24848 12747 -24588
rect 12677 -24858 12747 -24848
rect 12347 -24868 12427 -24858
rect 12347 -24928 12357 -24868
rect 12417 -24878 12427 -24868
rect 12667 -24868 12747 -24858
rect 12667 -24878 12677 -24868
rect 12417 -24928 12677 -24878
rect 12737 -24928 12747 -24868
rect 12347 -24938 12747 -24928
rect 12803 -24518 13203 -24508
rect 12803 -24578 12813 -24518
rect 12873 -24568 13133 -24518
rect 12873 -24578 12883 -24568
rect 12803 -24588 12883 -24578
rect 13123 -24578 13133 -24568
rect 13193 -24578 13203 -24518
rect 13123 -24588 13203 -24578
rect 12803 -24858 12863 -24588
rect 12943 -24648 12973 -24628
rect 12923 -24688 12973 -24648
rect 13033 -24648 13063 -24628
rect 13033 -24688 13083 -24648
rect 12923 -24758 13083 -24688
rect 12923 -24798 12973 -24758
rect 12943 -24818 12973 -24798
rect 13033 -24798 13083 -24758
rect 13033 -24818 13063 -24798
rect 13143 -24848 13203 -24588
rect 13133 -24858 13203 -24848
rect 12803 -24868 12883 -24858
rect 12803 -24928 12813 -24868
rect 12873 -24878 12883 -24868
rect 13123 -24868 13203 -24858
rect 13123 -24878 13133 -24868
rect 12873 -24928 13133 -24878
rect 13193 -24928 13203 -24868
rect 12803 -24938 13203 -24928
rect 13261 -24518 13661 -24508
rect 13261 -24578 13271 -24518
rect 13331 -24568 13591 -24518
rect 13331 -24578 13341 -24568
rect 13261 -24588 13341 -24578
rect 13581 -24578 13591 -24568
rect 13651 -24578 13661 -24518
rect 13581 -24588 13661 -24578
rect 13261 -24858 13321 -24588
rect 13401 -24648 13431 -24628
rect 13381 -24688 13431 -24648
rect 13491 -24648 13521 -24628
rect 13491 -24688 13541 -24648
rect 13381 -24758 13541 -24688
rect 13381 -24798 13431 -24758
rect 13401 -24818 13431 -24798
rect 13491 -24798 13541 -24758
rect 13491 -24818 13521 -24798
rect 13601 -24848 13661 -24588
rect 13591 -24858 13661 -24848
rect 13261 -24868 13341 -24858
rect 13261 -24928 13271 -24868
rect 13331 -24878 13341 -24868
rect 13581 -24868 13661 -24858
rect 13581 -24878 13591 -24868
rect 13331 -24928 13591 -24878
rect 13651 -24928 13661 -24868
rect 13261 -24938 13661 -24928
rect 13717 -24518 14117 -24508
rect 13717 -24578 13727 -24518
rect 13787 -24568 14047 -24518
rect 13787 -24578 13797 -24568
rect 13717 -24588 13797 -24578
rect 14037 -24578 14047 -24568
rect 14107 -24578 14117 -24518
rect 14037 -24588 14117 -24578
rect 13717 -24858 13777 -24588
rect 13857 -24648 13887 -24628
rect 13837 -24688 13887 -24648
rect 13947 -24648 13977 -24628
rect 13947 -24688 13997 -24648
rect 13837 -24758 13997 -24688
rect 13837 -24798 13887 -24758
rect 13857 -24818 13887 -24798
rect 13947 -24798 13997 -24758
rect 13947 -24818 13977 -24798
rect 14057 -24848 14117 -24588
rect 14047 -24858 14117 -24848
rect 13717 -24868 13797 -24858
rect 13717 -24928 13727 -24868
rect 13787 -24878 13797 -24868
rect 14037 -24868 14117 -24858
rect 14037 -24878 14047 -24868
rect 13787 -24928 14047 -24878
rect 14107 -24928 14117 -24868
rect 13717 -24938 14117 -24928
rect 14173 -24518 14573 -24508
rect 14173 -24578 14183 -24518
rect 14243 -24568 14503 -24518
rect 14243 -24578 14253 -24568
rect 14173 -24588 14253 -24578
rect 14493 -24578 14503 -24568
rect 14563 -24578 14573 -24518
rect 14493 -24588 14573 -24578
rect 14173 -24858 14233 -24588
rect 14313 -24648 14343 -24628
rect 14293 -24688 14343 -24648
rect 14403 -24648 14433 -24628
rect 14403 -24688 14453 -24648
rect 14293 -24758 14453 -24688
rect 14293 -24798 14343 -24758
rect 14313 -24818 14343 -24798
rect 14403 -24798 14453 -24758
rect 14403 -24818 14433 -24798
rect 14513 -24848 14573 -24588
rect 14503 -24858 14573 -24848
rect 14173 -24868 14253 -24858
rect 14173 -24928 14183 -24868
rect 14243 -24878 14253 -24868
rect 14493 -24868 14573 -24858
rect 14493 -24878 14503 -24868
rect 14243 -24928 14503 -24878
rect 14563 -24928 14573 -24868
rect 14173 -24938 14573 -24928
rect 14631 -24518 15031 -24508
rect 14631 -24578 14641 -24518
rect 14701 -24568 14961 -24518
rect 14701 -24578 14711 -24568
rect 14631 -24588 14711 -24578
rect 14951 -24578 14961 -24568
rect 15021 -24578 15031 -24518
rect 14951 -24588 15031 -24578
rect 14631 -24858 14691 -24588
rect 14771 -24648 14801 -24628
rect 14751 -24688 14801 -24648
rect 14861 -24648 14891 -24628
rect 14861 -24688 14911 -24648
rect 14751 -24758 14911 -24688
rect 14751 -24798 14801 -24758
rect 14771 -24818 14801 -24798
rect 14861 -24798 14911 -24758
rect 14861 -24818 14891 -24798
rect 14971 -24848 15031 -24588
rect 14961 -24858 15031 -24848
rect 14631 -24868 14711 -24858
rect 14631 -24928 14641 -24868
rect 14701 -24878 14711 -24868
rect 14951 -24868 15031 -24858
rect 14951 -24878 14961 -24868
rect 14701 -24928 14961 -24878
rect 15021 -24928 15031 -24868
rect 14631 -24938 15031 -24928
rect 15087 -24518 15487 -24508
rect 15087 -24578 15097 -24518
rect 15157 -24568 15417 -24518
rect 15157 -24578 15167 -24568
rect 15087 -24588 15167 -24578
rect 15407 -24578 15417 -24568
rect 15477 -24578 15487 -24518
rect 15407 -24588 15487 -24578
rect 15087 -24858 15147 -24588
rect 15227 -24648 15257 -24628
rect 15207 -24688 15257 -24648
rect 15317 -24648 15347 -24628
rect 15317 -24688 15367 -24648
rect 15207 -24758 15367 -24688
rect 15207 -24798 15257 -24758
rect 15227 -24818 15257 -24798
rect 15317 -24798 15367 -24758
rect 15317 -24818 15347 -24798
rect 15427 -24848 15487 -24588
rect 15417 -24858 15487 -24848
rect 15087 -24868 15167 -24858
rect 15087 -24928 15097 -24868
rect 15157 -24878 15167 -24868
rect 15407 -24868 15487 -24858
rect 15407 -24878 15417 -24868
rect 15157 -24928 15417 -24878
rect 15477 -24928 15487 -24868
rect 15087 -24938 15487 -24928
rect 1 -25034 401 -25024
rect 1 -25094 11 -25034
rect 71 -25084 331 -25034
rect 71 -25094 81 -25084
rect 1 -25104 81 -25094
rect 321 -25094 331 -25084
rect 391 -25094 401 -25034
rect 321 -25104 401 -25094
rect 1 -25374 61 -25104
rect 141 -25164 171 -25144
rect 121 -25204 171 -25164
rect 231 -25164 261 -25144
rect 231 -25204 281 -25164
rect 121 -25274 281 -25204
rect 121 -25314 171 -25274
rect 141 -25334 171 -25314
rect 231 -25314 281 -25274
rect 231 -25334 261 -25314
rect 341 -25364 401 -25104
rect 331 -25374 401 -25364
rect 1 -25384 81 -25374
rect 1 -25444 11 -25384
rect 71 -25394 81 -25384
rect 321 -25384 401 -25374
rect 321 -25394 331 -25384
rect 71 -25444 331 -25394
rect 391 -25444 401 -25384
rect 1 -25454 401 -25444
rect 457 -25034 857 -25024
rect 457 -25094 467 -25034
rect 527 -25084 787 -25034
rect 527 -25094 537 -25084
rect 457 -25104 537 -25094
rect 777 -25094 787 -25084
rect 847 -25094 857 -25034
rect 777 -25104 857 -25094
rect 457 -25374 517 -25104
rect 597 -25164 627 -25144
rect 577 -25204 627 -25164
rect 687 -25164 717 -25144
rect 687 -25204 737 -25164
rect 577 -25274 737 -25204
rect 577 -25314 627 -25274
rect 597 -25334 627 -25314
rect 687 -25314 737 -25274
rect 687 -25334 717 -25314
rect 797 -25364 857 -25104
rect 787 -25374 857 -25364
rect 457 -25384 537 -25374
rect 457 -25444 467 -25384
rect 527 -25394 537 -25384
rect 777 -25384 857 -25374
rect 777 -25394 787 -25384
rect 527 -25444 787 -25394
rect 847 -25444 857 -25384
rect 457 -25454 857 -25444
rect 913 -25034 1313 -25024
rect 913 -25094 923 -25034
rect 983 -25084 1243 -25034
rect 983 -25094 993 -25084
rect 913 -25104 993 -25094
rect 1233 -25094 1243 -25084
rect 1303 -25094 1313 -25034
rect 1233 -25104 1313 -25094
rect 913 -25374 973 -25104
rect 1053 -25164 1083 -25144
rect 1033 -25204 1083 -25164
rect 1143 -25164 1173 -25144
rect 1143 -25204 1193 -25164
rect 1033 -25274 1193 -25204
rect 1033 -25314 1083 -25274
rect 1053 -25334 1083 -25314
rect 1143 -25314 1193 -25274
rect 1143 -25334 1173 -25314
rect 1253 -25364 1313 -25104
rect 1243 -25374 1313 -25364
rect 913 -25384 993 -25374
rect 913 -25444 923 -25384
rect 983 -25394 993 -25384
rect 1233 -25384 1313 -25374
rect 1233 -25394 1243 -25384
rect 983 -25444 1243 -25394
rect 1303 -25444 1313 -25384
rect 913 -25454 1313 -25444
rect 1371 -25034 1771 -25024
rect 1371 -25094 1381 -25034
rect 1441 -25084 1701 -25034
rect 1441 -25094 1451 -25084
rect 1371 -25104 1451 -25094
rect 1691 -25094 1701 -25084
rect 1761 -25094 1771 -25034
rect 1691 -25104 1771 -25094
rect 1371 -25374 1431 -25104
rect 1511 -25164 1541 -25144
rect 1491 -25204 1541 -25164
rect 1601 -25164 1631 -25144
rect 1601 -25204 1651 -25164
rect 1491 -25274 1651 -25204
rect 1491 -25314 1541 -25274
rect 1511 -25334 1541 -25314
rect 1601 -25314 1651 -25274
rect 1601 -25334 1631 -25314
rect 1711 -25364 1771 -25104
rect 1701 -25374 1771 -25364
rect 1371 -25384 1451 -25374
rect 1371 -25444 1381 -25384
rect 1441 -25394 1451 -25384
rect 1691 -25384 1771 -25374
rect 1691 -25394 1701 -25384
rect 1441 -25444 1701 -25394
rect 1761 -25444 1771 -25384
rect 1371 -25454 1771 -25444
rect 1827 -25034 2227 -25024
rect 1827 -25094 1837 -25034
rect 1897 -25084 2157 -25034
rect 1897 -25094 1907 -25084
rect 1827 -25104 1907 -25094
rect 2147 -25094 2157 -25084
rect 2217 -25094 2227 -25034
rect 2147 -25104 2227 -25094
rect 1827 -25374 1887 -25104
rect 1967 -25164 1997 -25144
rect 1947 -25204 1997 -25164
rect 2057 -25164 2087 -25144
rect 2057 -25204 2107 -25164
rect 1947 -25274 2107 -25204
rect 1947 -25314 1997 -25274
rect 1967 -25334 1997 -25314
rect 2057 -25314 2107 -25274
rect 2057 -25334 2087 -25314
rect 2167 -25364 2227 -25104
rect 2157 -25374 2227 -25364
rect 1827 -25384 1907 -25374
rect 1827 -25444 1837 -25384
rect 1897 -25394 1907 -25384
rect 2147 -25384 2227 -25374
rect 2147 -25394 2157 -25384
rect 1897 -25444 2157 -25394
rect 2217 -25444 2227 -25384
rect 1827 -25454 2227 -25444
rect 2283 -25034 2683 -25024
rect 2283 -25094 2293 -25034
rect 2353 -25084 2613 -25034
rect 2353 -25094 2363 -25084
rect 2283 -25104 2363 -25094
rect 2603 -25094 2613 -25084
rect 2673 -25094 2683 -25034
rect 2603 -25104 2683 -25094
rect 2283 -25374 2343 -25104
rect 2423 -25164 2453 -25144
rect 2403 -25204 2453 -25164
rect 2513 -25164 2543 -25144
rect 2513 -25204 2563 -25164
rect 2403 -25274 2563 -25204
rect 2403 -25314 2453 -25274
rect 2423 -25334 2453 -25314
rect 2513 -25314 2563 -25274
rect 2513 -25334 2543 -25314
rect 2623 -25364 2683 -25104
rect 2613 -25374 2683 -25364
rect 2283 -25384 2363 -25374
rect 2283 -25444 2293 -25384
rect 2353 -25394 2363 -25384
rect 2603 -25384 2683 -25374
rect 2603 -25394 2613 -25384
rect 2353 -25444 2613 -25394
rect 2673 -25444 2683 -25384
rect 2283 -25454 2683 -25444
rect 2741 -25034 3141 -25024
rect 2741 -25094 2751 -25034
rect 2811 -25084 3071 -25034
rect 2811 -25094 2821 -25084
rect 2741 -25104 2821 -25094
rect 3061 -25094 3071 -25084
rect 3131 -25094 3141 -25034
rect 3061 -25104 3141 -25094
rect 2741 -25374 2801 -25104
rect 2881 -25164 2911 -25144
rect 2861 -25204 2911 -25164
rect 2971 -25164 3001 -25144
rect 2971 -25204 3021 -25164
rect 2861 -25274 3021 -25204
rect 2861 -25314 2911 -25274
rect 2881 -25334 2911 -25314
rect 2971 -25314 3021 -25274
rect 2971 -25334 3001 -25314
rect 3081 -25364 3141 -25104
rect 3071 -25374 3141 -25364
rect 2741 -25384 2821 -25374
rect 2741 -25444 2751 -25384
rect 2811 -25394 2821 -25384
rect 3061 -25384 3141 -25374
rect 3061 -25394 3071 -25384
rect 2811 -25444 3071 -25394
rect 3131 -25444 3141 -25384
rect 2741 -25454 3141 -25444
rect 3197 -25034 3597 -25024
rect 3197 -25094 3207 -25034
rect 3267 -25084 3527 -25034
rect 3267 -25094 3277 -25084
rect 3197 -25104 3277 -25094
rect 3517 -25094 3527 -25084
rect 3587 -25094 3597 -25034
rect 3517 -25104 3597 -25094
rect 3197 -25374 3257 -25104
rect 3337 -25164 3367 -25144
rect 3317 -25204 3367 -25164
rect 3427 -25164 3457 -25144
rect 3427 -25204 3477 -25164
rect 3317 -25274 3477 -25204
rect 3317 -25314 3367 -25274
rect 3337 -25334 3367 -25314
rect 3427 -25314 3477 -25274
rect 3427 -25334 3457 -25314
rect 3537 -25364 3597 -25104
rect 3527 -25374 3597 -25364
rect 3197 -25384 3277 -25374
rect 3197 -25444 3207 -25384
rect 3267 -25394 3277 -25384
rect 3517 -25384 3597 -25374
rect 3517 -25394 3527 -25384
rect 3267 -25444 3527 -25394
rect 3587 -25444 3597 -25384
rect 3197 -25454 3597 -25444
rect 3653 -25034 4053 -25024
rect 3653 -25094 3663 -25034
rect 3723 -25084 3983 -25034
rect 3723 -25094 3733 -25084
rect 3653 -25104 3733 -25094
rect 3973 -25094 3983 -25084
rect 4043 -25094 4053 -25034
rect 3973 -25104 4053 -25094
rect 3653 -25374 3713 -25104
rect 3793 -25164 3823 -25144
rect 3773 -25204 3823 -25164
rect 3883 -25164 3913 -25144
rect 3883 -25204 3933 -25164
rect 3773 -25274 3933 -25204
rect 3773 -25314 3823 -25274
rect 3793 -25334 3823 -25314
rect 3883 -25314 3933 -25274
rect 3883 -25334 3913 -25314
rect 3993 -25364 4053 -25104
rect 3983 -25374 4053 -25364
rect 3653 -25384 3733 -25374
rect 3653 -25444 3663 -25384
rect 3723 -25394 3733 -25384
rect 3973 -25384 4053 -25374
rect 3973 -25394 3983 -25384
rect 3723 -25444 3983 -25394
rect 4043 -25444 4053 -25384
rect 3653 -25454 4053 -25444
rect 4111 -25034 4511 -25024
rect 4111 -25094 4121 -25034
rect 4181 -25084 4441 -25034
rect 4181 -25094 4191 -25084
rect 4111 -25104 4191 -25094
rect 4431 -25094 4441 -25084
rect 4501 -25094 4511 -25034
rect 4431 -25104 4511 -25094
rect 4111 -25374 4171 -25104
rect 4251 -25164 4281 -25144
rect 4231 -25204 4281 -25164
rect 4341 -25164 4371 -25144
rect 4341 -25204 4391 -25164
rect 4231 -25274 4391 -25204
rect 4231 -25314 4281 -25274
rect 4251 -25334 4281 -25314
rect 4341 -25314 4391 -25274
rect 4341 -25334 4371 -25314
rect 4451 -25364 4511 -25104
rect 4441 -25374 4511 -25364
rect 4111 -25384 4191 -25374
rect 4111 -25444 4121 -25384
rect 4181 -25394 4191 -25384
rect 4431 -25384 4511 -25374
rect 4431 -25394 4441 -25384
rect 4181 -25444 4441 -25394
rect 4501 -25444 4511 -25384
rect 4111 -25454 4511 -25444
rect 4567 -25034 4967 -25024
rect 4567 -25094 4577 -25034
rect 4637 -25084 4897 -25034
rect 4637 -25094 4647 -25084
rect 4567 -25104 4647 -25094
rect 4887 -25094 4897 -25084
rect 4957 -25094 4967 -25034
rect 4887 -25104 4967 -25094
rect 4567 -25374 4627 -25104
rect 4707 -25164 4737 -25144
rect 4687 -25204 4737 -25164
rect 4797 -25164 4827 -25144
rect 4797 -25204 4847 -25164
rect 4687 -25274 4847 -25204
rect 4687 -25314 4737 -25274
rect 4707 -25334 4737 -25314
rect 4797 -25314 4847 -25274
rect 4797 -25334 4827 -25314
rect 4907 -25364 4967 -25104
rect 4897 -25374 4967 -25364
rect 4567 -25384 4647 -25374
rect 4567 -25444 4577 -25384
rect 4637 -25394 4647 -25384
rect 4887 -25384 4967 -25374
rect 4887 -25394 4897 -25384
rect 4637 -25444 4897 -25394
rect 4957 -25444 4967 -25384
rect 4567 -25454 4967 -25444
rect 5023 -25034 5423 -25024
rect 5023 -25094 5033 -25034
rect 5093 -25084 5353 -25034
rect 5093 -25094 5103 -25084
rect 5023 -25104 5103 -25094
rect 5343 -25094 5353 -25084
rect 5413 -25094 5423 -25034
rect 5343 -25104 5423 -25094
rect 5023 -25374 5083 -25104
rect 5163 -25164 5193 -25144
rect 5143 -25204 5193 -25164
rect 5253 -25164 5283 -25144
rect 5253 -25204 5303 -25164
rect 5143 -25274 5303 -25204
rect 5143 -25314 5193 -25274
rect 5163 -25334 5193 -25314
rect 5253 -25314 5303 -25274
rect 5253 -25334 5283 -25314
rect 5363 -25364 5423 -25104
rect 5353 -25374 5423 -25364
rect 5023 -25384 5103 -25374
rect 5023 -25444 5033 -25384
rect 5093 -25394 5103 -25384
rect 5343 -25384 5423 -25374
rect 5343 -25394 5353 -25384
rect 5093 -25444 5353 -25394
rect 5413 -25444 5423 -25384
rect 5023 -25454 5423 -25444
rect 5481 -25034 5881 -25024
rect 5481 -25094 5491 -25034
rect 5551 -25084 5811 -25034
rect 5551 -25094 5561 -25084
rect 5481 -25104 5561 -25094
rect 5801 -25094 5811 -25084
rect 5871 -25094 5881 -25034
rect 5801 -25104 5881 -25094
rect 5481 -25374 5541 -25104
rect 5621 -25164 5651 -25144
rect 5601 -25204 5651 -25164
rect 5711 -25164 5741 -25144
rect 5711 -25204 5761 -25164
rect 5601 -25274 5761 -25204
rect 5601 -25314 5651 -25274
rect 5621 -25334 5651 -25314
rect 5711 -25314 5761 -25274
rect 5711 -25334 5741 -25314
rect 5821 -25364 5881 -25104
rect 5811 -25374 5881 -25364
rect 5481 -25384 5561 -25374
rect 5481 -25444 5491 -25384
rect 5551 -25394 5561 -25384
rect 5801 -25384 5881 -25374
rect 5801 -25394 5811 -25384
rect 5551 -25444 5811 -25394
rect 5871 -25444 5881 -25384
rect 5481 -25454 5881 -25444
rect 5937 -25034 6337 -25024
rect 5937 -25094 5947 -25034
rect 6007 -25084 6267 -25034
rect 6007 -25094 6017 -25084
rect 5937 -25104 6017 -25094
rect 6257 -25094 6267 -25084
rect 6327 -25094 6337 -25034
rect 6257 -25104 6337 -25094
rect 5937 -25374 5997 -25104
rect 6077 -25164 6107 -25144
rect 6057 -25204 6107 -25164
rect 6167 -25164 6197 -25144
rect 6167 -25204 6217 -25164
rect 6057 -25274 6217 -25204
rect 6057 -25314 6107 -25274
rect 6077 -25334 6107 -25314
rect 6167 -25314 6217 -25274
rect 6167 -25334 6197 -25314
rect 6277 -25364 6337 -25104
rect 6267 -25374 6337 -25364
rect 5937 -25384 6017 -25374
rect 5937 -25444 5947 -25384
rect 6007 -25394 6017 -25384
rect 6257 -25384 6337 -25374
rect 6257 -25394 6267 -25384
rect 6007 -25444 6267 -25394
rect 6327 -25444 6337 -25384
rect 5937 -25454 6337 -25444
rect 6393 -25034 6793 -25024
rect 6393 -25094 6403 -25034
rect 6463 -25084 6723 -25034
rect 6463 -25094 6473 -25084
rect 6393 -25104 6473 -25094
rect 6713 -25094 6723 -25084
rect 6783 -25094 6793 -25034
rect 6713 -25104 6793 -25094
rect 6393 -25374 6453 -25104
rect 6533 -25164 6563 -25144
rect 6513 -25204 6563 -25164
rect 6623 -25164 6653 -25144
rect 6623 -25204 6673 -25164
rect 6513 -25274 6673 -25204
rect 6513 -25314 6563 -25274
rect 6533 -25334 6563 -25314
rect 6623 -25314 6673 -25274
rect 6623 -25334 6653 -25314
rect 6733 -25364 6793 -25104
rect 6723 -25374 6793 -25364
rect 6393 -25384 6473 -25374
rect 6393 -25444 6403 -25384
rect 6463 -25394 6473 -25384
rect 6713 -25384 6793 -25374
rect 6713 -25394 6723 -25384
rect 6463 -25444 6723 -25394
rect 6783 -25444 6793 -25384
rect 6393 -25454 6793 -25444
rect 6851 -25034 7251 -25024
rect 6851 -25094 6861 -25034
rect 6921 -25084 7181 -25034
rect 6921 -25094 6931 -25084
rect 6851 -25104 6931 -25094
rect 7171 -25094 7181 -25084
rect 7241 -25094 7251 -25034
rect 7171 -25104 7251 -25094
rect 6851 -25374 6911 -25104
rect 6991 -25164 7021 -25144
rect 6971 -25204 7021 -25164
rect 7081 -25164 7111 -25144
rect 7081 -25204 7131 -25164
rect 6971 -25274 7131 -25204
rect 6971 -25314 7021 -25274
rect 6991 -25334 7021 -25314
rect 7081 -25314 7131 -25274
rect 7081 -25334 7111 -25314
rect 7191 -25364 7251 -25104
rect 7181 -25374 7251 -25364
rect 6851 -25384 6931 -25374
rect 6851 -25444 6861 -25384
rect 6921 -25394 6931 -25384
rect 7171 -25384 7251 -25374
rect 7171 -25394 7181 -25384
rect 6921 -25444 7181 -25394
rect 7241 -25444 7251 -25384
rect 6851 -25454 7251 -25444
rect 7307 -25034 7707 -25024
rect 7307 -25094 7317 -25034
rect 7377 -25084 7637 -25034
rect 7377 -25094 7387 -25084
rect 7307 -25104 7387 -25094
rect 7627 -25094 7637 -25084
rect 7697 -25094 7707 -25034
rect 7627 -25104 7707 -25094
rect 7307 -25374 7367 -25104
rect 7447 -25164 7477 -25144
rect 7427 -25204 7477 -25164
rect 7537 -25164 7567 -25144
rect 7537 -25204 7587 -25164
rect 7427 -25274 7587 -25204
rect 7427 -25314 7477 -25274
rect 7447 -25334 7477 -25314
rect 7537 -25314 7587 -25274
rect 7537 -25334 7567 -25314
rect 7647 -25364 7707 -25104
rect 7637 -25374 7707 -25364
rect 7307 -25384 7387 -25374
rect 7307 -25444 7317 -25384
rect 7377 -25394 7387 -25384
rect 7627 -25384 7707 -25374
rect 7627 -25394 7637 -25384
rect 7377 -25444 7637 -25394
rect 7697 -25444 7707 -25384
rect 7307 -25454 7707 -25444
rect 7763 -25034 8163 -25024
rect 7763 -25094 7773 -25034
rect 7833 -25084 8093 -25034
rect 7833 -25094 7843 -25084
rect 7763 -25104 7843 -25094
rect 8083 -25094 8093 -25084
rect 8153 -25094 8163 -25034
rect 8083 -25104 8163 -25094
rect 7763 -25374 7823 -25104
rect 7903 -25164 7933 -25144
rect 7883 -25204 7933 -25164
rect 7993 -25164 8023 -25144
rect 7993 -25204 8043 -25164
rect 7883 -25274 8043 -25204
rect 7883 -25314 7933 -25274
rect 7903 -25334 7933 -25314
rect 7993 -25314 8043 -25274
rect 7993 -25334 8023 -25314
rect 8103 -25364 8163 -25104
rect 8093 -25374 8163 -25364
rect 7763 -25384 7843 -25374
rect 7763 -25444 7773 -25384
rect 7833 -25394 7843 -25384
rect 8083 -25384 8163 -25374
rect 8083 -25394 8093 -25384
rect 7833 -25444 8093 -25394
rect 8153 -25444 8163 -25384
rect 7763 -25454 8163 -25444
rect 8237 -25034 8637 -25024
rect 8237 -25094 8247 -25034
rect 8307 -25084 8567 -25034
rect 8307 -25094 8317 -25084
rect 8237 -25104 8317 -25094
rect 8557 -25094 8567 -25084
rect 8627 -25094 8637 -25034
rect 8557 -25104 8637 -25094
rect 8237 -25374 8297 -25104
rect 8377 -25164 8407 -25144
rect 8357 -25204 8407 -25164
rect 8467 -25164 8497 -25144
rect 8467 -25204 8517 -25164
rect 8357 -25274 8517 -25204
rect 8357 -25314 8407 -25274
rect 8377 -25334 8407 -25314
rect 8467 -25314 8517 -25274
rect 8467 -25334 8497 -25314
rect 8577 -25364 8637 -25104
rect 8567 -25374 8637 -25364
rect 8237 -25384 8317 -25374
rect 8237 -25444 8247 -25384
rect 8307 -25394 8317 -25384
rect 8557 -25384 8637 -25374
rect 8557 -25394 8567 -25384
rect 8307 -25444 8567 -25394
rect 8627 -25444 8637 -25384
rect 8237 -25454 8637 -25444
rect 8693 -25034 9093 -25024
rect 8693 -25094 8703 -25034
rect 8763 -25084 9023 -25034
rect 8763 -25094 8773 -25084
rect 8693 -25104 8773 -25094
rect 9013 -25094 9023 -25084
rect 9083 -25094 9093 -25034
rect 9013 -25104 9093 -25094
rect 8693 -25374 8753 -25104
rect 8833 -25164 8863 -25144
rect 8813 -25204 8863 -25164
rect 8923 -25164 8953 -25144
rect 8923 -25204 8973 -25164
rect 8813 -25274 8973 -25204
rect 8813 -25314 8863 -25274
rect 8833 -25334 8863 -25314
rect 8923 -25314 8973 -25274
rect 8923 -25334 8953 -25314
rect 9033 -25364 9093 -25104
rect 9023 -25374 9093 -25364
rect 8693 -25384 8773 -25374
rect 8693 -25444 8703 -25384
rect 8763 -25394 8773 -25384
rect 9013 -25384 9093 -25374
rect 9013 -25394 9023 -25384
rect 8763 -25444 9023 -25394
rect 9083 -25444 9093 -25384
rect 8693 -25454 9093 -25444
rect 9151 -25034 9551 -25024
rect 9151 -25094 9161 -25034
rect 9221 -25084 9481 -25034
rect 9221 -25094 9231 -25084
rect 9151 -25104 9231 -25094
rect 9471 -25094 9481 -25084
rect 9541 -25094 9551 -25034
rect 9471 -25104 9551 -25094
rect 9151 -25374 9211 -25104
rect 9291 -25164 9321 -25144
rect 9271 -25204 9321 -25164
rect 9381 -25164 9411 -25144
rect 9381 -25204 9431 -25164
rect 9271 -25274 9431 -25204
rect 9271 -25314 9321 -25274
rect 9291 -25334 9321 -25314
rect 9381 -25314 9431 -25274
rect 9381 -25334 9411 -25314
rect 9491 -25364 9551 -25104
rect 9481 -25374 9551 -25364
rect 9151 -25384 9231 -25374
rect 9151 -25444 9161 -25384
rect 9221 -25394 9231 -25384
rect 9471 -25384 9551 -25374
rect 9471 -25394 9481 -25384
rect 9221 -25444 9481 -25394
rect 9541 -25444 9551 -25384
rect 9151 -25454 9551 -25444
rect 9607 -25034 10007 -25024
rect 9607 -25094 9617 -25034
rect 9677 -25084 9937 -25034
rect 9677 -25094 9687 -25084
rect 9607 -25104 9687 -25094
rect 9927 -25094 9937 -25084
rect 9997 -25094 10007 -25034
rect 9927 -25104 10007 -25094
rect 9607 -25374 9667 -25104
rect 9747 -25164 9777 -25144
rect 9727 -25204 9777 -25164
rect 9837 -25164 9867 -25144
rect 9837 -25204 9887 -25164
rect 9727 -25274 9887 -25204
rect 9727 -25314 9777 -25274
rect 9747 -25334 9777 -25314
rect 9837 -25314 9887 -25274
rect 9837 -25334 9867 -25314
rect 9947 -25364 10007 -25104
rect 9937 -25374 10007 -25364
rect 9607 -25384 9687 -25374
rect 9607 -25444 9617 -25384
rect 9677 -25394 9687 -25384
rect 9927 -25384 10007 -25374
rect 9927 -25394 9937 -25384
rect 9677 -25444 9937 -25394
rect 9997 -25444 10007 -25384
rect 9607 -25454 10007 -25444
rect 10063 -25034 10463 -25024
rect 10063 -25094 10073 -25034
rect 10133 -25084 10393 -25034
rect 10133 -25094 10143 -25084
rect 10063 -25104 10143 -25094
rect 10383 -25094 10393 -25084
rect 10453 -25094 10463 -25034
rect 10383 -25104 10463 -25094
rect 10063 -25374 10123 -25104
rect 10203 -25164 10233 -25144
rect 10183 -25204 10233 -25164
rect 10293 -25164 10323 -25144
rect 10293 -25204 10343 -25164
rect 10183 -25274 10343 -25204
rect 10183 -25314 10233 -25274
rect 10203 -25334 10233 -25314
rect 10293 -25314 10343 -25274
rect 10293 -25334 10323 -25314
rect 10403 -25364 10463 -25104
rect 10393 -25374 10463 -25364
rect 10063 -25384 10143 -25374
rect 10063 -25444 10073 -25384
rect 10133 -25394 10143 -25384
rect 10383 -25384 10463 -25374
rect 10383 -25394 10393 -25384
rect 10133 -25444 10393 -25394
rect 10453 -25444 10463 -25384
rect 10063 -25454 10463 -25444
rect 10521 -25034 10921 -25024
rect 10521 -25094 10531 -25034
rect 10591 -25084 10851 -25034
rect 10591 -25094 10601 -25084
rect 10521 -25104 10601 -25094
rect 10841 -25094 10851 -25084
rect 10911 -25094 10921 -25034
rect 10841 -25104 10921 -25094
rect 10521 -25374 10581 -25104
rect 10661 -25164 10691 -25144
rect 10641 -25204 10691 -25164
rect 10751 -25164 10781 -25144
rect 10751 -25204 10801 -25164
rect 10641 -25274 10801 -25204
rect 10641 -25314 10691 -25274
rect 10661 -25334 10691 -25314
rect 10751 -25314 10801 -25274
rect 10751 -25334 10781 -25314
rect 10861 -25364 10921 -25104
rect 10851 -25374 10921 -25364
rect 10521 -25384 10601 -25374
rect 10521 -25444 10531 -25384
rect 10591 -25394 10601 -25384
rect 10841 -25384 10921 -25374
rect 10841 -25394 10851 -25384
rect 10591 -25444 10851 -25394
rect 10911 -25444 10921 -25384
rect 10521 -25454 10921 -25444
rect 10977 -25034 11377 -25024
rect 10977 -25094 10987 -25034
rect 11047 -25084 11307 -25034
rect 11047 -25094 11057 -25084
rect 10977 -25104 11057 -25094
rect 11297 -25094 11307 -25084
rect 11367 -25094 11377 -25034
rect 11297 -25104 11377 -25094
rect 10977 -25374 11037 -25104
rect 11117 -25164 11147 -25144
rect 11097 -25204 11147 -25164
rect 11207 -25164 11237 -25144
rect 11207 -25204 11257 -25164
rect 11097 -25274 11257 -25204
rect 11097 -25314 11147 -25274
rect 11117 -25334 11147 -25314
rect 11207 -25314 11257 -25274
rect 11207 -25334 11237 -25314
rect 11317 -25364 11377 -25104
rect 11307 -25374 11377 -25364
rect 10977 -25384 11057 -25374
rect 10977 -25444 10987 -25384
rect 11047 -25394 11057 -25384
rect 11297 -25384 11377 -25374
rect 11297 -25394 11307 -25384
rect 11047 -25444 11307 -25394
rect 11367 -25444 11377 -25384
rect 10977 -25454 11377 -25444
rect 11433 -25034 11833 -25024
rect 11433 -25094 11443 -25034
rect 11503 -25084 11763 -25034
rect 11503 -25094 11513 -25084
rect 11433 -25104 11513 -25094
rect 11753 -25094 11763 -25084
rect 11823 -25094 11833 -25034
rect 11753 -25104 11833 -25094
rect 11433 -25374 11493 -25104
rect 11573 -25164 11603 -25144
rect 11553 -25204 11603 -25164
rect 11663 -25164 11693 -25144
rect 11663 -25204 11713 -25164
rect 11553 -25274 11713 -25204
rect 11553 -25314 11603 -25274
rect 11573 -25334 11603 -25314
rect 11663 -25314 11713 -25274
rect 11663 -25334 11693 -25314
rect 11773 -25364 11833 -25104
rect 11763 -25374 11833 -25364
rect 11433 -25384 11513 -25374
rect 11433 -25444 11443 -25384
rect 11503 -25394 11513 -25384
rect 11753 -25384 11833 -25374
rect 11753 -25394 11763 -25384
rect 11503 -25444 11763 -25394
rect 11823 -25444 11833 -25384
rect 11433 -25454 11833 -25444
rect 11891 -25034 12291 -25024
rect 11891 -25094 11901 -25034
rect 11961 -25084 12221 -25034
rect 11961 -25094 11971 -25084
rect 11891 -25104 11971 -25094
rect 12211 -25094 12221 -25084
rect 12281 -25094 12291 -25034
rect 12211 -25104 12291 -25094
rect 11891 -25374 11951 -25104
rect 12031 -25164 12061 -25144
rect 12011 -25204 12061 -25164
rect 12121 -25164 12151 -25144
rect 12121 -25204 12171 -25164
rect 12011 -25274 12171 -25204
rect 12011 -25314 12061 -25274
rect 12031 -25334 12061 -25314
rect 12121 -25314 12171 -25274
rect 12121 -25334 12151 -25314
rect 12231 -25364 12291 -25104
rect 12221 -25374 12291 -25364
rect 11891 -25384 11971 -25374
rect 11891 -25444 11901 -25384
rect 11961 -25394 11971 -25384
rect 12211 -25384 12291 -25374
rect 12211 -25394 12221 -25384
rect 11961 -25444 12221 -25394
rect 12281 -25444 12291 -25384
rect 11891 -25454 12291 -25444
rect 12347 -25034 12747 -25024
rect 12347 -25094 12357 -25034
rect 12417 -25084 12677 -25034
rect 12417 -25094 12427 -25084
rect 12347 -25104 12427 -25094
rect 12667 -25094 12677 -25084
rect 12737 -25094 12747 -25034
rect 12667 -25104 12747 -25094
rect 12347 -25374 12407 -25104
rect 12487 -25164 12517 -25144
rect 12467 -25204 12517 -25164
rect 12577 -25164 12607 -25144
rect 12577 -25204 12627 -25164
rect 12467 -25274 12627 -25204
rect 12467 -25314 12517 -25274
rect 12487 -25334 12517 -25314
rect 12577 -25314 12627 -25274
rect 12577 -25334 12607 -25314
rect 12687 -25364 12747 -25104
rect 12677 -25374 12747 -25364
rect 12347 -25384 12427 -25374
rect 12347 -25444 12357 -25384
rect 12417 -25394 12427 -25384
rect 12667 -25384 12747 -25374
rect 12667 -25394 12677 -25384
rect 12417 -25444 12677 -25394
rect 12737 -25444 12747 -25384
rect 12347 -25454 12747 -25444
rect 12803 -25034 13203 -25024
rect 12803 -25094 12813 -25034
rect 12873 -25084 13133 -25034
rect 12873 -25094 12883 -25084
rect 12803 -25104 12883 -25094
rect 13123 -25094 13133 -25084
rect 13193 -25094 13203 -25034
rect 13123 -25104 13203 -25094
rect 12803 -25374 12863 -25104
rect 12943 -25164 12973 -25144
rect 12923 -25204 12973 -25164
rect 13033 -25164 13063 -25144
rect 13033 -25204 13083 -25164
rect 12923 -25274 13083 -25204
rect 12923 -25314 12973 -25274
rect 12943 -25334 12973 -25314
rect 13033 -25314 13083 -25274
rect 13033 -25334 13063 -25314
rect 13143 -25364 13203 -25104
rect 13133 -25374 13203 -25364
rect 12803 -25384 12883 -25374
rect 12803 -25444 12813 -25384
rect 12873 -25394 12883 -25384
rect 13123 -25384 13203 -25374
rect 13123 -25394 13133 -25384
rect 12873 -25444 13133 -25394
rect 13193 -25444 13203 -25384
rect 12803 -25454 13203 -25444
rect 13261 -25034 13661 -25024
rect 13261 -25094 13271 -25034
rect 13331 -25084 13591 -25034
rect 13331 -25094 13341 -25084
rect 13261 -25104 13341 -25094
rect 13581 -25094 13591 -25084
rect 13651 -25094 13661 -25034
rect 13581 -25104 13661 -25094
rect 13261 -25374 13321 -25104
rect 13401 -25164 13431 -25144
rect 13381 -25204 13431 -25164
rect 13491 -25164 13521 -25144
rect 13491 -25204 13541 -25164
rect 13381 -25274 13541 -25204
rect 13381 -25314 13431 -25274
rect 13401 -25334 13431 -25314
rect 13491 -25314 13541 -25274
rect 13491 -25334 13521 -25314
rect 13601 -25364 13661 -25104
rect 13591 -25374 13661 -25364
rect 13261 -25384 13341 -25374
rect 13261 -25444 13271 -25384
rect 13331 -25394 13341 -25384
rect 13581 -25384 13661 -25374
rect 13581 -25394 13591 -25384
rect 13331 -25444 13591 -25394
rect 13651 -25444 13661 -25384
rect 13261 -25454 13661 -25444
rect 13717 -25034 14117 -25024
rect 13717 -25094 13727 -25034
rect 13787 -25084 14047 -25034
rect 13787 -25094 13797 -25084
rect 13717 -25104 13797 -25094
rect 14037 -25094 14047 -25084
rect 14107 -25094 14117 -25034
rect 14037 -25104 14117 -25094
rect 13717 -25374 13777 -25104
rect 13857 -25164 13887 -25144
rect 13837 -25204 13887 -25164
rect 13947 -25164 13977 -25144
rect 13947 -25204 13997 -25164
rect 13837 -25274 13997 -25204
rect 13837 -25314 13887 -25274
rect 13857 -25334 13887 -25314
rect 13947 -25314 13997 -25274
rect 13947 -25334 13977 -25314
rect 14057 -25364 14117 -25104
rect 14047 -25374 14117 -25364
rect 13717 -25384 13797 -25374
rect 13717 -25444 13727 -25384
rect 13787 -25394 13797 -25384
rect 14037 -25384 14117 -25374
rect 14037 -25394 14047 -25384
rect 13787 -25444 14047 -25394
rect 14107 -25444 14117 -25384
rect 13717 -25454 14117 -25444
rect 14173 -25034 14573 -25024
rect 14173 -25094 14183 -25034
rect 14243 -25084 14503 -25034
rect 14243 -25094 14253 -25084
rect 14173 -25104 14253 -25094
rect 14493 -25094 14503 -25084
rect 14563 -25094 14573 -25034
rect 14493 -25104 14573 -25094
rect 14173 -25374 14233 -25104
rect 14313 -25164 14343 -25144
rect 14293 -25204 14343 -25164
rect 14403 -25164 14433 -25144
rect 14403 -25204 14453 -25164
rect 14293 -25274 14453 -25204
rect 14293 -25314 14343 -25274
rect 14313 -25334 14343 -25314
rect 14403 -25314 14453 -25274
rect 14403 -25334 14433 -25314
rect 14513 -25364 14573 -25104
rect 14503 -25374 14573 -25364
rect 14173 -25384 14253 -25374
rect 14173 -25444 14183 -25384
rect 14243 -25394 14253 -25384
rect 14493 -25384 14573 -25374
rect 14493 -25394 14503 -25384
rect 14243 -25444 14503 -25394
rect 14563 -25444 14573 -25384
rect 14173 -25454 14573 -25444
rect 14631 -25034 15031 -25024
rect 14631 -25094 14641 -25034
rect 14701 -25084 14961 -25034
rect 14701 -25094 14711 -25084
rect 14631 -25104 14711 -25094
rect 14951 -25094 14961 -25084
rect 15021 -25094 15031 -25034
rect 14951 -25104 15031 -25094
rect 14631 -25374 14691 -25104
rect 14771 -25164 14801 -25144
rect 14751 -25204 14801 -25164
rect 14861 -25164 14891 -25144
rect 14861 -25204 14911 -25164
rect 14751 -25274 14911 -25204
rect 14751 -25314 14801 -25274
rect 14771 -25334 14801 -25314
rect 14861 -25314 14911 -25274
rect 14861 -25334 14891 -25314
rect 14971 -25364 15031 -25104
rect 14961 -25374 15031 -25364
rect 14631 -25384 14711 -25374
rect 14631 -25444 14641 -25384
rect 14701 -25394 14711 -25384
rect 14951 -25384 15031 -25374
rect 14951 -25394 14961 -25384
rect 14701 -25444 14961 -25394
rect 15021 -25444 15031 -25384
rect 14631 -25454 15031 -25444
rect 15087 -25034 15487 -25024
rect 15087 -25094 15097 -25034
rect 15157 -25084 15417 -25034
rect 15157 -25094 15167 -25084
rect 15087 -25104 15167 -25094
rect 15407 -25094 15417 -25084
rect 15477 -25094 15487 -25034
rect 15407 -25104 15487 -25094
rect 15087 -25374 15147 -25104
rect 15227 -25164 15257 -25144
rect 15207 -25204 15257 -25164
rect 15317 -25164 15347 -25144
rect 15317 -25204 15367 -25164
rect 15207 -25274 15367 -25204
rect 15207 -25314 15257 -25274
rect 15227 -25334 15257 -25314
rect 15317 -25314 15367 -25274
rect 15317 -25334 15347 -25314
rect 15427 -25364 15487 -25104
rect 15417 -25374 15487 -25364
rect 15087 -25384 15167 -25374
rect 15087 -25444 15097 -25384
rect 15157 -25394 15167 -25384
rect 15407 -25384 15487 -25374
rect 15407 -25394 15417 -25384
rect 15157 -25444 15417 -25394
rect 15477 -25444 15487 -25384
rect 15087 -25454 15487 -25444
rect 1 -25526 401 -25516
rect 1 -25586 11 -25526
rect 71 -25576 331 -25526
rect 71 -25586 81 -25576
rect 1 -25596 81 -25586
rect 321 -25586 331 -25576
rect 391 -25586 401 -25526
rect 321 -25596 401 -25586
rect 1 -25866 61 -25596
rect 141 -25656 171 -25636
rect 121 -25696 171 -25656
rect 231 -25656 261 -25636
rect 231 -25696 281 -25656
rect 121 -25766 281 -25696
rect 121 -25806 171 -25766
rect 141 -25826 171 -25806
rect 231 -25806 281 -25766
rect 231 -25826 261 -25806
rect 341 -25856 401 -25596
rect 331 -25866 401 -25856
rect 1 -25876 81 -25866
rect 1 -25936 11 -25876
rect 71 -25886 81 -25876
rect 321 -25876 401 -25866
rect 321 -25886 331 -25876
rect 71 -25936 331 -25886
rect 391 -25936 401 -25876
rect 1 -25946 401 -25936
rect 457 -25526 857 -25516
rect 457 -25586 467 -25526
rect 527 -25576 787 -25526
rect 527 -25586 537 -25576
rect 457 -25596 537 -25586
rect 777 -25586 787 -25576
rect 847 -25586 857 -25526
rect 777 -25596 857 -25586
rect 457 -25866 517 -25596
rect 597 -25656 627 -25636
rect 577 -25696 627 -25656
rect 687 -25656 717 -25636
rect 687 -25696 737 -25656
rect 577 -25766 737 -25696
rect 577 -25806 627 -25766
rect 597 -25826 627 -25806
rect 687 -25806 737 -25766
rect 687 -25826 717 -25806
rect 797 -25856 857 -25596
rect 787 -25866 857 -25856
rect 457 -25876 537 -25866
rect 457 -25936 467 -25876
rect 527 -25886 537 -25876
rect 777 -25876 857 -25866
rect 777 -25886 787 -25876
rect 527 -25936 787 -25886
rect 847 -25936 857 -25876
rect 457 -25946 857 -25936
rect 913 -25526 1313 -25516
rect 913 -25586 923 -25526
rect 983 -25576 1243 -25526
rect 983 -25586 993 -25576
rect 913 -25596 993 -25586
rect 1233 -25586 1243 -25576
rect 1303 -25586 1313 -25526
rect 1233 -25596 1313 -25586
rect 913 -25866 973 -25596
rect 1053 -25656 1083 -25636
rect 1033 -25696 1083 -25656
rect 1143 -25656 1173 -25636
rect 1143 -25696 1193 -25656
rect 1033 -25766 1193 -25696
rect 1033 -25806 1083 -25766
rect 1053 -25826 1083 -25806
rect 1143 -25806 1193 -25766
rect 1143 -25826 1173 -25806
rect 1253 -25856 1313 -25596
rect 1243 -25866 1313 -25856
rect 913 -25876 993 -25866
rect 913 -25936 923 -25876
rect 983 -25886 993 -25876
rect 1233 -25876 1313 -25866
rect 1233 -25886 1243 -25876
rect 983 -25936 1243 -25886
rect 1303 -25936 1313 -25876
rect 913 -25946 1313 -25936
rect 1371 -25526 1771 -25516
rect 1371 -25586 1381 -25526
rect 1441 -25576 1701 -25526
rect 1441 -25586 1451 -25576
rect 1371 -25596 1451 -25586
rect 1691 -25586 1701 -25576
rect 1761 -25586 1771 -25526
rect 1691 -25596 1771 -25586
rect 1371 -25866 1431 -25596
rect 1511 -25656 1541 -25636
rect 1491 -25696 1541 -25656
rect 1601 -25656 1631 -25636
rect 1601 -25696 1651 -25656
rect 1491 -25766 1651 -25696
rect 1491 -25806 1541 -25766
rect 1511 -25826 1541 -25806
rect 1601 -25806 1651 -25766
rect 1601 -25826 1631 -25806
rect 1711 -25856 1771 -25596
rect 1701 -25866 1771 -25856
rect 1371 -25876 1451 -25866
rect 1371 -25936 1381 -25876
rect 1441 -25886 1451 -25876
rect 1691 -25876 1771 -25866
rect 1691 -25886 1701 -25876
rect 1441 -25936 1701 -25886
rect 1761 -25936 1771 -25876
rect 1371 -25946 1771 -25936
rect 1827 -25526 2227 -25516
rect 1827 -25586 1837 -25526
rect 1897 -25576 2157 -25526
rect 1897 -25586 1907 -25576
rect 1827 -25596 1907 -25586
rect 2147 -25586 2157 -25576
rect 2217 -25586 2227 -25526
rect 2147 -25596 2227 -25586
rect 1827 -25866 1887 -25596
rect 1967 -25656 1997 -25636
rect 1947 -25696 1997 -25656
rect 2057 -25656 2087 -25636
rect 2057 -25696 2107 -25656
rect 1947 -25766 2107 -25696
rect 1947 -25806 1997 -25766
rect 1967 -25826 1997 -25806
rect 2057 -25806 2107 -25766
rect 2057 -25826 2087 -25806
rect 2167 -25856 2227 -25596
rect 2157 -25866 2227 -25856
rect 1827 -25876 1907 -25866
rect 1827 -25936 1837 -25876
rect 1897 -25886 1907 -25876
rect 2147 -25876 2227 -25866
rect 2147 -25886 2157 -25876
rect 1897 -25936 2157 -25886
rect 2217 -25936 2227 -25876
rect 1827 -25946 2227 -25936
rect 2283 -25526 2683 -25516
rect 2283 -25586 2293 -25526
rect 2353 -25576 2613 -25526
rect 2353 -25586 2363 -25576
rect 2283 -25596 2363 -25586
rect 2603 -25586 2613 -25576
rect 2673 -25586 2683 -25526
rect 2603 -25596 2683 -25586
rect 2283 -25866 2343 -25596
rect 2423 -25656 2453 -25636
rect 2403 -25696 2453 -25656
rect 2513 -25656 2543 -25636
rect 2513 -25696 2563 -25656
rect 2403 -25766 2563 -25696
rect 2403 -25806 2453 -25766
rect 2423 -25826 2453 -25806
rect 2513 -25806 2563 -25766
rect 2513 -25826 2543 -25806
rect 2623 -25856 2683 -25596
rect 2613 -25866 2683 -25856
rect 2283 -25876 2363 -25866
rect 2283 -25936 2293 -25876
rect 2353 -25886 2363 -25876
rect 2603 -25876 2683 -25866
rect 2603 -25886 2613 -25876
rect 2353 -25936 2613 -25886
rect 2673 -25936 2683 -25876
rect 2283 -25946 2683 -25936
rect 2741 -25526 3141 -25516
rect 2741 -25586 2751 -25526
rect 2811 -25576 3071 -25526
rect 2811 -25586 2821 -25576
rect 2741 -25596 2821 -25586
rect 3061 -25586 3071 -25576
rect 3131 -25586 3141 -25526
rect 3061 -25596 3141 -25586
rect 2741 -25866 2801 -25596
rect 2881 -25656 2911 -25636
rect 2861 -25696 2911 -25656
rect 2971 -25656 3001 -25636
rect 2971 -25696 3021 -25656
rect 2861 -25766 3021 -25696
rect 2861 -25806 2911 -25766
rect 2881 -25826 2911 -25806
rect 2971 -25806 3021 -25766
rect 2971 -25826 3001 -25806
rect 3081 -25856 3141 -25596
rect 3071 -25866 3141 -25856
rect 2741 -25876 2821 -25866
rect 2741 -25936 2751 -25876
rect 2811 -25886 2821 -25876
rect 3061 -25876 3141 -25866
rect 3061 -25886 3071 -25876
rect 2811 -25936 3071 -25886
rect 3131 -25936 3141 -25876
rect 2741 -25946 3141 -25936
rect 3197 -25526 3597 -25516
rect 3197 -25586 3207 -25526
rect 3267 -25576 3527 -25526
rect 3267 -25586 3277 -25576
rect 3197 -25596 3277 -25586
rect 3517 -25586 3527 -25576
rect 3587 -25586 3597 -25526
rect 3517 -25596 3597 -25586
rect 3197 -25866 3257 -25596
rect 3337 -25656 3367 -25636
rect 3317 -25696 3367 -25656
rect 3427 -25656 3457 -25636
rect 3427 -25696 3477 -25656
rect 3317 -25766 3477 -25696
rect 3317 -25806 3367 -25766
rect 3337 -25826 3367 -25806
rect 3427 -25806 3477 -25766
rect 3427 -25826 3457 -25806
rect 3537 -25856 3597 -25596
rect 3527 -25866 3597 -25856
rect 3197 -25876 3277 -25866
rect 3197 -25936 3207 -25876
rect 3267 -25886 3277 -25876
rect 3517 -25876 3597 -25866
rect 3517 -25886 3527 -25876
rect 3267 -25936 3527 -25886
rect 3587 -25936 3597 -25876
rect 3197 -25946 3597 -25936
rect 3653 -25526 4053 -25516
rect 3653 -25586 3663 -25526
rect 3723 -25576 3983 -25526
rect 3723 -25586 3733 -25576
rect 3653 -25596 3733 -25586
rect 3973 -25586 3983 -25576
rect 4043 -25586 4053 -25526
rect 3973 -25596 4053 -25586
rect 3653 -25866 3713 -25596
rect 3793 -25656 3823 -25636
rect 3773 -25696 3823 -25656
rect 3883 -25656 3913 -25636
rect 3883 -25696 3933 -25656
rect 3773 -25766 3933 -25696
rect 3773 -25806 3823 -25766
rect 3793 -25826 3823 -25806
rect 3883 -25806 3933 -25766
rect 3883 -25826 3913 -25806
rect 3993 -25856 4053 -25596
rect 3983 -25866 4053 -25856
rect 3653 -25876 3733 -25866
rect 3653 -25936 3663 -25876
rect 3723 -25886 3733 -25876
rect 3973 -25876 4053 -25866
rect 3973 -25886 3983 -25876
rect 3723 -25936 3983 -25886
rect 4043 -25936 4053 -25876
rect 3653 -25946 4053 -25936
rect 4111 -25526 4511 -25516
rect 4111 -25586 4121 -25526
rect 4181 -25576 4441 -25526
rect 4181 -25586 4191 -25576
rect 4111 -25596 4191 -25586
rect 4431 -25586 4441 -25576
rect 4501 -25586 4511 -25526
rect 4431 -25596 4511 -25586
rect 4111 -25866 4171 -25596
rect 4251 -25656 4281 -25636
rect 4231 -25696 4281 -25656
rect 4341 -25656 4371 -25636
rect 4341 -25696 4391 -25656
rect 4231 -25766 4391 -25696
rect 4231 -25806 4281 -25766
rect 4251 -25826 4281 -25806
rect 4341 -25806 4391 -25766
rect 4341 -25826 4371 -25806
rect 4451 -25856 4511 -25596
rect 4441 -25866 4511 -25856
rect 4111 -25876 4191 -25866
rect 4111 -25936 4121 -25876
rect 4181 -25886 4191 -25876
rect 4431 -25876 4511 -25866
rect 4431 -25886 4441 -25876
rect 4181 -25936 4441 -25886
rect 4501 -25936 4511 -25876
rect 4111 -25946 4511 -25936
rect 4567 -25526 4967 -25516
rect 4567 -25586 4577 -25526
rect 4637 -25576 4897 -25526
rect 4637 -25586 4647 -25576
rect 4567 -25596 4647 -25586
rect 4887 -25586 4897 -25576
rect 4957 -25586 4967 -25526
rect 4887 -25596 4967 -25586
rect 4567 -25866 4627 -25596
rect 4707 -25656 4737 -25636
rect 4687 -25696 4737 -25656
rect 4797 -25656 4827 -25636
rect 4797 -25696 4847 -25656
rect 4687 -25766 4847 -25696
rect 4687 -25806 4737 -25766
rect 4707 -25826 4737 -25806
rect 4797 -25806 4847 -25766
rect 4797 -25826 4827 -25806
rect 4907 -25856 4967 -25596
rect 4897 -25866 4967 -25856
rect 4567 -25876 4647 -25866
rect 4567 -25936 4577 -25876
rect 4637 -25886 4647 -25876
rect 4887 -25876 4967 -25866
rect 4887 -25886 4897 -25876
rect 4637 -25936 4897 -25886
rect 4957 -25936 4967 -25876
rect 4567 -25946 4967 -25936
rect 5023 -25526 5423 -25516
rect 5023 -25586 5033 -25526
rect 5093 -25576 5353 -25526
rect 5093 -25586 5103 -25576
rect 5023 -25596 5103 -25586
rect 5343 -25586 5353 -25576
rect 5413 -25586 5423 -25526
rect 5343 -25596 5423 -25586
rect 5023 -25866 5083 -25596
rect 5163 -25656 5193 -25636
rect 5143 -25696 5193 -25656
rect 5253 -25656 5283 -25636
rect 5253 -25696 5303 -25656
rect 5143 -25766 5303 -25696
rect 5143 -25806 5193 -25766
rect 5163 -25826 5193 -25806
rect 5253 -25806 5303 -25766
rect 5253 -25826 5283 -25806
rect 5363 -25856 5423 -25596
rect 5353 -25866 5423 -25856
rect 5023 -25876 5103 -25866
rect 5023 -25936 5033 -25876
rect 5093 -25886 5103 -25876
rect 5343 -25876 5423 -25866
rect 5343 -25886 5353 -25876
rect 5093 -25936 5353 -25886
rect 5413 -25936 5423 -25876
rect 5023 -25946 5423 -25936
rect 5481 -25526 5881 -25516
rect 5481 -25586 5491 -25526
rect 5551 -25576 5811 -25526
rect 5551 -25586 5561 -25576
rect 5481 -25596 5561 -25586
rect 5801 -25586 5811 -25576
rect 5871 -25586 5881 -25526
rect 5801 -25596 5881 -25586
rect 5481 -25866 5541 -25596
rect 5621 -25656 5651 -25636
rect 5601 -25696 5651 -25656
rect 5711 -25656 5741 -25636
rect 5711 -25696 5761 -25656
rect 5601 -25766 5761 -25696
rect 5601 -25806 5651 -25766
rect 5621 -25826 5651 -25806
rect 5711 -25806 5761 -25766
rect 5711 -25826 5741 -25806
rect 5821 -25856 5881 -25596
rect 5811 -25866 5881 -25856
rect 5481 -25876 5561 -25866
rect 5481 -25936 5491 -25876
rect 5551 -25886 5561 -25876
rect 5801 -25876 5881 -25866
rect 5801 -25886 5811 -25876
rect 5551 -25936 5811 -25886
rect 5871 -25936 5881 -25876
rect 5481 -25946 5881 -25936
rect 5937 -25526 6337 -25516
rect 5937 -25586 5947 -25526
rect 6007 -25576 6267 -25526
rect 6007 -25586 6017 -25576
rect 5937 -25596 6017 -25586
rect 6257 -25586 6267 -25576
rect 6327 -25586 6337 -25526
rect 6257 -25596 6337 -25586
rect 5937 -25866 5997 -25596
rect 6077 -25656 6107 -25636
rect 6057 -25696 6107 -25656
rect 6167 -25656 6197 -25636
rect 6167 -25696 6217 -25656
rect 6057 -25766 6217 -25696
rect 6057 -25806 6107 -25766
rect 6077 -25826 6107 -25806
rect 6167 -25806 6217 -25766
rect 6167 -25826 6197 -25806
rect 6277 -25856 6337 -25596
rect 6267 -25866 6337 -25856
rect 5937 -25876 6017 -25866
rect 5937 -25936 5947 -25876
rect 6007 -25886 6017 -25876
rect 6257 -25876 6337 -25866
rect 6257 -25886 6267 -25876
rect 6007 -25936 6267 -25886
rect 6327 -25936 6337 -25876
rect 5937 -25946 6337 -25936
rect 6393 -25526 6793 -25516
rect 6393 -25586 6403 -25526
rect 6463 -25576 6723 -25526
rect 6463 -25586 6473 -25576
rect 6393 -25596 6473 -25586
rect 6713 -25586 6723 -25576
rect 6783 -25586 6793 -25526
rect 6713 -25596 6793 -25586
rect 6393 -25866 6453 -25596
rect 6533 -25656 6563 -25636
rect 6513 -25696 6563 -25656
rect 6623 -25656 6653 -25636
rect 6623 -25696 6673 -25656
rect 6513 -25766 6673 -25696
rect 6513 -25806 6563 -25766
rect 6533 -25826 6563 -25806
rect 6623 -25806 6673 -25766
rect 6623 -25826 6653 -25806
rect 6733 -25856 6793 -25596
rect 6723 -25866 6793 -25856
rect 6393 -25876 6473 -25866
rect 6393 -25936 6403 -25876
rect 6463 -25886 6473 -25876
rect 6713 -25876 6793 -25866
rect 6713 -25886 6723 -25876
rect 6463 -25936 6723 -25886
rect 6783 -25936 6793 -25876
rect 6393 -25946 6793 -25936
rect 6851 -25526 7251 -25516
rect 6851 -25586 6861 -25526
rect 6921 -25576 7181 -25526
rect 6921 -25586 6931 -25576
rect 6851 -25596 6931 -25586
rect 7171 -25586 7181 -25576
rect 7241 -25586 7251 -25526
rect 7171 -25596 7251 -25586
rect 6851 -25866 6911 -25596
rect 6991 -25656 7021 -25636
rect 6971 -25696 7021 -25656
rect 7081 -25656 7111 -25636
rect 7081 -25696 7131 -25656
rect 6971 -25766 7131 -25696
rect 6971 -25806 7021 -25766
rect 6991 -25826 7021 -25806
rect 7081 -25806 7131 -25766
rect 7081 -25826 7111 -25806
rect 7191 -25856 7251 -25596
rect 7181 -25866 7251 -25856
rect 6851 -25876 6931 -25866
rect 6851 -25936 6861 -25876
rect 6921 -25886 6931 -25876
rect 7171 -25876 7251 -25866
rect 7171 -25886 7181 -25876
rect 6921 -25936 7181 -25886
rect 7241 -25936 7251 -25876
rect 6851 -25946 7251 -25936
rect 7307 -25526 7707 -25516
rect 7307 -25586 7317 -25526
rect 7377 -25576 7637 -25526
rect 7377 -25586 7387 -25576
rect 7307 -25596 7387 -25586
rect 7627 -25586 7637 -25576
rect 7697 -25586 7707 -25526
rect 7627 -25596 7707 -25586
rect 7307 -25866 7367 -25596
rect 7447 -25656 7477 -25636
rect 7427 -25696 7477 -25656
rect 7537 -25656 7567 -25636
rect 7537 -25696 7587 -25656
rect 7427 -25766 7587 -25696
rect 7427 -25806 7477 -25766
rect 7447 -25826 7477 -25806
rect 7537 -25806 7587 -25766
rect 7537 -25826 7567 -25806
rect 7647 -25856 7707 -25596
rect 7637 -25866 7707 -25856
rect 7307 -25876 7387 -25866
rect 7307 -25936 7317 -25876
rect 7377 -25886 7387 -25876
rect 7627 -25876 7707 -25866
rect 7627 -25886 7637 -25876
rect 7377 -25936 7637 -25886
rect 7697 -25936 7707 -25876
rect 7307 -25946 7707 -25936
rect 7763 -25526 8163 -25516
rect 7763 -25586 7773 -25526
rect 7833 -25576 8093 -25526
rect 7833 -25586 7843 -25576
rect 7763 -25596 7843 -25586
rect 8083 -25586 8093 -25576
rect 8153 -25586 8163 -25526
rect 8083 -25596 8163 -25586
rect 7763 -25866 7823 -25596
rect 7903 -25656 7933 -25636
rect 7883 -25696 7933 -25656
rect 7993 -25656 8023 -25636
rect 7993 -25696 8043 -25656
rect 7883 -25766 8043 -25696
rect 7883 -25806 7933 -25766
rect 7903 -25826 7933 -25806
rect 7993 -25806 8043 -25766
rect 7993 -25826 8023 -25806
rect 8103 -25856 8163 -25596
rect 8093 -25866 8163 -25856
rect 7763 -25876 7843 -25866
rect 7763 -25936 7773 -25876
rect 7833 -25886 7843 -25876
rect 8083 -25876 8163 -25866
rect 8083 -25886 8093 -25876
rect 7833 -25936 8093 -25886
rect 8153 -25936 8163 -25876
rect 7763 -25946 8163 -25936
rect 8237 -25526 8637 -25516
rect 8237 -25586 8247 -25526
rect 8307 -25576 8567 -25526
rect 8307 -25586 8317 -25576
rect 8237 -25596 8317 -25586
rect 8557 -25586 8567 -25576
rect 8627 -25586 8637 -25526
rect 8557 -25596 8637 -25586
rect 8237 -25866 8297 -25596
rect 8377 -25656 8407 -25636
rect 8357 -25696 8407 -25656
rect 8467 -25656 8497 -25636
rect 8467 -25696 8517 -25656
rect 8357 -25766 8517 -25696
rect 8357 -25806 8407 -25766
rect 8377 -25826 8407 -25806
rect 8467 -25806 8517 -25766
rect 8467 -25826 8497 -25806
rect 8577 -25856 8637 -25596
rect 8567 -25866 8637 -25856
rect 8237 -25876 8317 -25866
rect 8237 -25936 8247 -25876
rect 8307 -25886 8317 -25876
rect 8557 -25876 8637 -25866
rect 8557 -25886 8567 -25876
rect 8307 -25936 8567 -25886
rect 8627 -25936 8637 -25876
rect 8237 -25946 8637 -25936
rect 8693 -25526 9093 -25516
rect 8693 -25586 8703 -25526
rect 8763 -25576 9023 -25526
rect 8763 -25586 8773 -25576
rect 8693 -25596 8773 -25586
rect 9013 -25586 9023 -25576
rect 9083 -25586 9093 -25526
rect 9013 -25596 9093 -25586
rect 8693 -25866 8753 -25596
rect 8833 -25656 8863 -25636
rect 8813 -25696 8863 -25656
rect 8923 -25656 8953 -25636
rect 8923 -25696 8973 -25656
rect 8813 -25766 8973 -25696
rect 8813 -25806 8863 -25766
rect 8833 -25826 8863 -25806
rect 8923 -25806 8973 -25766
rect 8923 -25826 8953 -25806
rect 9033 -25856 9093 -25596
rect 9023 -25866 9093 -25856
rect 8693 -25876 8773 -25866
rect 8693 -25936 8703 -25876
rect 8763 -25886 8773 -25876
rect 9013 -25876 9093 -25866
rect 9013 -25886 9023 -25876
rect 8763 -25936 9023 -25886
rect 9083 -25936 9093 -25876
rect 8693 -25946 9093 -25936
rect 9151 -25526 9551 -25516
rect 9151 -25586 9161 -25526
rect 9221 -25576 9481 -25526
rect 9221 -25586 9231 -25576
rect 9151 -25596 9231 -25586
rect 9471 -25586 9481 -25576
rect 9541 -25586 9551 -25526
rect 9471 -25596 9551 -25586
rect 9151 -25866 9211 -25596
rect 9291 -25656 9321 -25636
rect 9271 -25696 9321 -25656
rect 9381 -25656 9411 -25636
rect 9381 -25696 9431 -25656
rect 9271 -25766 9431 -25696
rect 9271 -25806 9321 -25766
rect 9291 -25826 9321 -25806
rect 9381 -25806 9431 -25766
rect 9381 -25826 9411 -25806
rect 9491 -25856 9551 -25596
rect 9481 -25866 9551 -25856
rect 9151 -25876 9231 -25866
rect 9151 -25936 9161 -25876
rect 9221 -25886 9231 -25876
rect 9471 -25876 9551 -25866
rect 9471 -25886 9481 -25876
rect 9221 -25936 9481 -25886
rect 9541 -25936 9551 -25876
rect 9151 -25946 9551 -25936
rect 9607 -25526 10007 -25516
rect 9607 -25586 9617 -25526
rect 9677 -25576 9937 -25526
rect 9677 -25586 9687 -25576
rect 9607 -25596 9687 -25586
rect 9927 -25586 9937 -25576
rect 9997 -25586 10007 -25526
rect 9927 -25596 10007 -25586
rect 9607 -25866 9667 -25596
rect 9747 -25656 9777 -25636
rect 9727 -25696 9777 -25656
rect 9837 -25656 9867 -25636
rect 9837 -25696 9887 -25656
rect 9727 -25766 9887 -25696
rect 9727 -25806 9777 -25766
rect 9747 -25826 9777 -25806
rect 9837 -25806 9887 -25766
rect 9837 -25826 9867 -25806
rect 9947 -25856 10007 -25596
rect 9937 -25866 10007 -25856
rect 9607 -25876 9687 -25866
rect 9607 -25936 9617 -25876
rect 9677 -25886 9687 -25876
rect 9927 -25876 10007 -25866
rect 9927 -25886 9937 -25876
rect 9677 -25936 9937 -25886
rect 9997 -25936 10007 -25876
rect 9607 -25946 10007 -25936
rect 10063 -25526 10463 -25516
rect 10063 -25586 10073 -25526
rect 10133 -25576 10393 -25526
rect 10133 -25586 10143 -25576
rect 10063 -25596 10143 -25586
rect 10383 -25586 10393 -25576
rect 10453 -25586 10463 -25526
rect 10383 -25596 10463 -25586
rect 10063 -25866 10123 -25596
rect 10203 -25656 10233 -25636
rect 10183 -25696 10233 -25656
rect 10293 -25656 10323 -25636
rect 10293 -25696 10343 -25656
rect 10183 -25766 10343 -25696
rect 10183 -25806 10233 -25766
rect 10203 -25826 10233 -25806
rect 10293 -25806 10343 -25766
rect 10293 -25826 10323 -25806
rect 10403 -25856 10463 -25596
rect 10393 -25866 10463 -25856
rect 10063 -25876 10143 -25866
rect 10063 -25936 10073 -25876
rect 10133 -25886 10143 -25876
rect 10383 -25876 10463 -25866
rect 10383 -25886 10393 -25876
rect 10133 -25936 10393 -25886
rect 10453 -25936 10463 -25876
rect 10063 -25946 10463 -25936
rect 10521 -25526 10921 -25516
rect 10521 -25586 10531 -25526
rect 10591 -25576 10851 -25526
rect 10591 -25586 10601 -25576
rect 10521 -25596 10601 -25586
rect 10841 -25586 10851 -25576
rect 10911 -25586 10921 -25526
rect 10841 -25596 10921 -25586
rect 10521 -25866 10581 -25596
rect 10661 -25656 10691 -25636
rect 10641 -25696 10691 -25656
rect 10751 -25656 10781 -25636
rect 10751 -25696 10801 -25656
rect 10641 -25766 10801 -25696
rect 10641 -25806 10691 -25766
rect 10661 -25826 10691 -25806
rect 10751 -25806 10801 -25766
rect 10751 -25826 10781 -25806
rect 10861 -25856 10921 -25596
rect 10851 -25866 10921 -25856
rect 10521 -25876 10601 -25866
rect 10521 -25936 10531 -25876
rect 10591 -25886 10601 -25876
rect 10841 -25876 10921 -25866
rect 10841 -25886 10851 -25876
rect 10591 -25936 10851 -25886
rect 10911 -25936 10921 -25876
rect 10521 -25946 10921 -25936
rect 10977 -25526 11377 -25516
rect 10977 -25586 10987 -25526
rect 11047 -25576 11307 -25526
rect 11047 -25586 11057 -25576
rect 10977 -25596 11057 -25586
rect 11297 -25586 11307 -25576
rect 11367 -25586 11377 -25526
rect 11297 -25596 11377 -25586
rect 10977 -25866 11037 -25596
rect 11117 -25656 11147 -25636
rect 11097 -25696 11147 -25656
rect 11207 -25656 11237 -25636
rect 11207 -25696 11257 -25656
rect 11097 -25766 11257 -25696
rect 11097 -25806 11147 -25766
rect 11117 -25826 11147 -25806
rect 11207 -25806 11257 -25766
rect 11207 -25826 11237 -25806
rect 11317 -25856 11377 -25596
rect 11307 -25866 11377 -25856
rect 10977 -25876 11057 -25866
rect 10977 -25936 10987 -25876
rect 11047 -25886 11057 -25876
rect 11297 -25876 11377 -25866
rect 11297 -25886 11307 -25876
rect 11047 -25936 11307 -25886
rect 11367 -25936 11377 -25876
rect 10977 -25946 11377 -25936
rect 11433 -25526 11833 -25516
rect 11433 -25586 11443 -25526
rect 11503 -25576 11763 -25526
rect 11503 -25586 11513 -25576
rect 11433 -25596 11513 -25586
rect 11753 -25586 11763 -25576
rect 11823 -25586 11833 -25526
rect 11753 -25596 11833 -25586
rect 11433 -25866 11493 -25596
rect 11573 -25656 11603 -25636
rect 11553 -25696 11603 -25656
rect 11663 -25656 11693 -25636
rect 11663 -25696 11713 -25656
rect 11553 -25766 11713 -25696
rect 11553 -25806 11603 -25766
rect 11573 -25826 11603 -25806
rect 11663 -25806 11713 -25766
rect 11663 -25826 11693 -25806
rect 11773 -25856 11833 -25596
rect 11763 -25866 11833 -25856
rect 11433 -25876 11513 -25866
rect 11433 -25936 11443 -25876
rect 11503 -25886 11513 -25876
rect 11753 -25876 11833 -25866
rect 11753 -25886 11763 -25876
rect 11503 -25936 11763 -25886
rect 11823 -25936 11833 -25876
rect 11433 -25946 11833 -25936
rect 11891 -25526 12291 -25516
rect 11891 -25586 11901 -25526
rect 11961 -25576 12221 -25526
rect 11961 -25586 11971 -25576
rect 11891 -25596 11971 -25586
rect 12211 -25586 12221 -25576
rect 12281 -25586 12291 -25526
rect 12211 -25596 12291 -25586
rect 11891 -25866 11951 -25596
rect 12031 -25656 12061 -25636
rect 12011 -25696 12061 -25656
rect 12121 -25656 12151 -25636
rect 12121 -25696 12171 -25656
rect 12011 -25766 12171 -25696
rect 12011 -25806 12061 -25766
rect 12031 -25826 12061 -25806
rect 12121 -25806 12171 -25766
rect 12121 -25826 12151 -25806
rect 12231 -25856 12291 -25596
rect 12221 -25866 12291 -25856
rect 11891 -25876 11971 -25866
rect 11891 -25936 11901 -25876
rect 11961 -25886 11971 -25876
rect 12211 -25876 12291 -25866
rect 12211 -25886 12221 -25876
rect 11961 -25936 12221 -25886
rect 12281 -25936 12291 -25876
rect 11891 -25946 12291 -25936
rect 12347 -25526 12747 -25516
rect 12347 -25586 12357 -25526
rect 12417 -25576 12677 -25526
rect 12417 -25586 12427 -25576
rect 12347 -25596 12427 -25586
rect 12667 -25586 12677 -25576
rect 12737 -25586 12747 -25526
rect 12667 -25596 12747 -25586
rect 12347 -25866 12407 -25596
rect 12487 -25656 12517 -25636
rect 12467 -25696 12517 -25656
rect 12577 -25656 12607 -25636
rect 12577 -25696 12627 -25656
rect 12467 -25766 12627 -25696
rect 12467 -25806 12517 -25766
rect 12487 -25826 12517 -25806
rect 12577 -25806 12627 -25766
rect 12577 -25826 12607 -25806
rect 12687 -25856 12747 -25596
rect 12677 -25866 12747 -25856
rect 12347 -25876 12427 -25866
rect 12347 -25936 12357 -25876
rect 12417 -25886 12427 -25876
rect 12667 -25876 12747 -25866
rect 12667 -25886 12677 -25876
rect 12417 -25936 12677 -25886
rect 12737 -25936 12747 -25876
rect 12347 -25946 12747 -25936
rect 12803 -25526 13203 -25516
rect 12803 -25586 12813 -25526
rect 12873 -25576 13133 -25526
rect 12873 -25586 12883 -25576
rect 12803 -25596 12883 -25586
rect 13123 -25586 13133 -25576
rect 13193 -25586 13203 -25526
rect 13123 -25596 13203 -25586
rect 12803 -25866 12863 -25596
rect 12943 -25656 12973 -25636
rect 12923 -25696 12973 -25656
rect 13033 -25656 13063 -25636
rect 13033 -25696 13083 -25656
rect 12923 -25766 13083 -25696
rect 12923 -25806 12973 -25766
rect 12943 -25826 12973 -25806
rect 13033 -25806 13083 -25766
rect 13033 -25826 13063 -25806
rect 13143 -25856 13203 -25596
rect 13133 -25866 13203 -25856
rect 12803 -25876 12883 -25866
rect 12803 -25936 12813 -25876
rect 12873 -25886 12883 -25876
rect 13123 -25876 13203 -25866
rect 13123 -25886 13133 -25876
rect 12873 -25936 13133 -25886
rect 13193 -25936 13203 -25876
rect 12803 -25946 13203 -25936
rect 13261 -25526 13661 -25516
rect 13261 -25586 13271 -25526
rect 13331 -25576 13591 -25526
rect 13331 -25586 13341 -25576
rect 13261 -25596 13341 -25586
rect 13581 -25586 13591 -25576
rect 13651 -25586 13661 -25526
rect 13581 -25596 13661 -25586
rect 13261 -25866 13321 -25596
rect 13401 -25656 13431 -25636
rect 13381 -25696 13431 -25656
rect 13491 -25656 13521 -25636
rect 13491 -25696 13541 -25656
rect 13381 -25766 13541 -25696
rect 13381 -25806 13431 -25766
rect 13401 -25826 13431 -25806
rect 13491 -25806 13541 -25766
rect 13491 -25826 13521 -25806
rect 13601 -25856 13661 -25596
rect 13591 -25866 13661 -25856
rect 13261 -25876 13341 -25866
rect 13261 -25936 13271 -25876
rect 13331 -25886 13341 -25876
rect 13581 -25876 13661 -25866
rect 13581 -25886 13591 -25876
rect 13331 -25936 13591 -25886
rect 13651 -25936 13661 -25876
rect 13261 -25946 13661 -25936
rect 13717 -25526 14117 -25516
rect 13717 -25586 13727 -25526
rect 13787 -25576 14047 -25526
rect 13787 -25586 13797 -25576
rect 13717 -25596 13797 -25586
rect 14037 -25586 14047 -25576
rect 14107 -25586 14117 -25526
rect 14037 -25596 14117 -25586
rect 13717 -25866 13777 -25596
rect 13857 -25656 13887 -25636
rect 13837 -25696 13887 -25656
rect 13947 -25656 13977 -25636
rect 13947 -25696 13997 -25656
rect 13837 -25766 13997 -25696
rect 13837 -25806 13887 -25766
rect 13857 -25826 13887 -25806
rect 13947 -25806 13997 -25766
rect 13947 -25826 13977 -25806
rect 14057 -25856 14117 -25596
rect 14047 -25866 14117 -25856
rect 13717 -25876 13797 -25866
rect 13717 -25936 13727 -25876
rect 13787 -25886 13797 -25876
rect 14037 -25876 14117 -25866
rect 14037 -25886 14047 -25876
rect 13787 -25936 14047 -25886
rect 14107 -25936 14117 -25876
rect 13717 -25946 14117 -25936
rect 14173 -25526 14573 -25516
rect 14173 -25586 14183 -25526
rect 14243 -25576 14503 -25526
rect 14243 -25586 14253 -25576
rect 14173 -25596 14253 -25586
rect 14493 -25586 14503 -25576
rect 14563 -25586 14573 -25526
rect 14493 -25596 14573 -25586
rect 14173 -25866 14233 -25596
rect 14313 -25656 14343 -25636
rect 14293 -25696 14343 -25656
rect 14403 -25656 14433 -25636
rect 14403 -25696 14453 -25656
rect 14293 -25766 14453 -25696
rect 14293 -25806 14343 -25766
rect 14313 -25826 14343 -25806
rect 14403 -25806 14453 -25766
rect 14403 -25826 14433 -25806
rect 14513 -25856 14573 -25596
rect 14503 -25866 14573 -25856
rect 14173 -25876 14253 -25866
rect 14173 -25936 14183 -25876
rect 14243 -25886 14253 -25876
rect 14493 -25876 14573 -25866
rect 14493 -25886 14503 -25876
rect 14243 -25936 14503 -25886
rect 14563 -25936 14573 -25876
rect 14173 -25946 14573 -25936
rect 14631 -25526 15031 -25516
rect 14631 -25586 14641 -25526
rect 14701 -25576 14961 -25526
rect 14701 -25586 14711 -25576
rect 14631 -25596 14711 -25586
rect 14951 -25586 14961 -25576
rect 15021 -25586 15031 -25526
rect 14951 -25596 15031 -25586
rect 14631 -25866 14691 -25596
rect 14771 -25656 14801 -25636
rect 14751 -25696 14801 -25656
rect 14861 -25656 14891 -25636
rect 14861 -25696 14911 -25656
rect 14751 -25766 14911 -25696
rect 14751 -25806 14801 -25766
rect 14771 -25826 14801 -25806
rect 14861 -25806 14911 -25766
rect 14861 -25826 14891 -25806
rect 14971 -25856 15031 -25596
rect 14961 -25866 15031 -25856
rect 14631 -25876 14711 -25866
rect 14631 -25936 14641 -25876
rect 14701 -25886 14711 -25876
rect 14951 -25876 15031 -25866
rect 14951 -25886 14961 -25876
rect 14701 -25936 14961 -25886
rect 15021 -25936 15031 -25876
rect 14631 -25946 15031 -25936
rect 15087 -25526 15487 -25516
rect 15087 -25586 15097 -25526
rect 15157 -25576 15417 -25526
rect 15157 -25586 15167 -25576
rect 15087 -25596 15167 -25586
rect 15407 -25586 15417 -25576
rect 15477 -25586 15487 -25526
rect 15407 -25596 15487 -25586
rect 15087 -25866 15147 -25596
rect 15227 -25656 15257 -25636
rect 15207 -25696 15257 -25656
rect 15317 -25656 15347 -25636
rect 15317 -25696 15367 -25656
rect 15207 -25766 15367 -25696
rect 15207 -25806 15257 -25766
rect 15227 -25826 15257 -25806
rect 15317 -25806 15367 -25766
rect 15317 -25826 15347 -25806
rect 15427 -25856 15487 -25596
rect 15417 -25866 15487 -25856
rect 15087 -25876 15167 -25866
rect 15087 -25936 15097 -25876
rect 15157 -25886 15167 -25876
rect 15407 -25876 15487 -25866
rect 15407 -25886 15417 -25876
rect 15157 -25936 15417 -25886
rect 15477 -25936 15487 -25876
rect 15087 -25946 15487 -25936
rect 0 -26023 400 -26013
rect 0 -26083 10 -26023
rect 70 -26073 330 -26023
rect 70 -26083 80 -26073
rect 0 -26093 80 -26083
rect 320 -26083 330 -26073
rect 390 -26083 400 -26023
rect 320 -26093 400 -26083
rect 0 -26363 60 -26093
rect 140 -26153 170 -26133
rect 120 -26193 170 -26153
rect 230 -26153 260 -26133
rect 230 -26193 280 -26153
rect 120 -26263 280 -26193
rect 120 -26303 170 -26263
rect 140 -26323 170 -26303
rect 230 -26303 280 -26263
rect 230 -26323 260 -26303
rect 340 -26353 400 -26093
rect 330 -26363 400 -26353
rect 0 -26373 80 -26363
rect 0 -26433 10 -26373
rect 70 -26383 80 -26373
rect 320 -26373 400 -26363
rect 320 -26383 330 -26373
rect 70 -26433 330 -26383
rect 390 -26433 400 -26373
rect 0 -26443 400 -26433
rect 456 -26023 856 -26013
rect 456 -26083 466 -26023
rect 526 -26073 786 -26023
rect 526 -26083 536 -26073
rect 456 -26093 536 -26083
rect 776 -26083 786 -26073
rect 846 -26083 856 -26023
rect 776 -26093 856 -26083
rect 456 -26363 516 -26093
rect 596 -26153 626 -26133
rect 576 -26193 626 -26153
rect 686 -26153 716 -26133
rect 686 -26193 736 -26153
rect 576 -26263 736 -26193
rect 576 -26303 626 -26263
rect 596 -26323 626 -26303
rect 686 -26303 736 -26263
rect 686 -26323 716 -26303
rect 796 -26353 856 -26093
rect 786 -26363 856 -26353
rect 456 -26373 536 -26363
rect 456 -26433 466 -26373
rect 526 -26383 536 -26373
rect 776 -26373 856 -26363
rect 776 -26383 786 -26373
rect 526 -26433 786 -26383
rect 846 -26433 856 -26373
rect 456 -26443 856 -26433
rect 912 -26023 1312 -26013
rect 912 -26083 922 -26023
rect 982 -26073 1242 -26023
rect 982 -26083 992 -26073
rect 912 -26093 992 -26083
rect 1232 -26083 1242 -26073
rect 1302 -26083 1312 -26023
rect 1232 -26093 1312 -26083
rect 912 -26363 972 -26093
rect 1052 -26153 1082 -26133
rect 1032 -26193 1082 -26153
rect 1142 -26153 1172 -26133
rect 1142 -26193 1192 -26153
rect 1032 -26263 1192 -26193
rect 1032 -26303 1082 -26263
rect 1052 -26323 1082 -26303
rect 1142 -26303 1192 -26263
rect 1142 -26323 1172 -26303
rect 1252 -26353 1312 -26093
rect 1242 -26363 1312 -26353
rect 912 -26373 992 -26363
rect 912 -26433 922 -26373
rect 982 -26383 992 -26373
rect 1232 -26373 1312 -26363
rect 1232 -26383 1242 -26373
rect 982 -26433 1242 -26383
rect 1302 -26433 1312 -26373
rect 912 -26443 1312 -26433
rect 1370 -26023 1770 -26013
rect 1370 -26083 1380 -26023
rect 1440 -26073 1700 -26023
rect 1440 -26083 1450 -26073
rect 1370 -26093 1450 -26083
rect 1690 -26083 1700 -26073
rect 1760 -26083 1770 -26023
rect 1690 -26093 1770 -26083
rect 1370 -26363 1430 -26093
rect 1510 -26153 1540 -26133
rect 1490 -26193 1540 -26153
rect 1600 -26153 1630 -26133
rect 1600 -26193 1650 -26153
rect 1490 -26263 1650 -26193
rect 1490 -26303 1540 -26263
rect 1510 -26323 1540 -26303
rect 1600 -26303 1650 -26263
rect 1600 -26323 1630 -26303
rect 1710 -26353 1770 -26093
rect 1700 -26363 1770 -26353
rect 1370 -26373 1450 -26363
rect 1370 -26433 1380 -26373
rect 1440 -26383 1450 -26373
rect 1690 -26373 1770 -26363
rect 1690 -26383 1700 -26373
rect 1440 -26433 1700 -26383
rect 1760 -26433 1770 -26373
rect 1370 -26443 1770 -26433
rect 1826 -26023 2226 -26013
rect 1826 -26083 1836 -26023
rect 1896 -26073 2156 -26023
rect 1896 -26083 1906 -26073
rect 1826 -26093 1906 -26083
rect 2146 -26083 2156 -26073
rect 2216 -26083 2226 -26023
rect 2146 -26093 2226 -26083
rect 1826 -26363 1886 -26093
rect 1966 -26153 1996 -26133
rect 1946 -26193 1996 -26153
rect 2056 -26153 2086 -26133
rect 2056 -26193 2106 -26153
rect 1946 -26263 2106 -26193
rect 1946 -26303 1996 -26263
rect 1966 -26323 1996 -26303
rect 2056 -26303 2106 -26263
rect 2056 -26323 2086 -26303
rect 2166 -26353 2226 -26093
rect 2156 -26363 2226 -26353
rect 1826 -26373 1906 -26363
rect 1826 -26433 1836 -26373
rect 1896 -26383 1906 -26373
rect 2146 -26373 2226 -26363
rect 2146 -26383 2156 -26373
rect 1896 -26433 2156 -26383
rect 2216 -26433 2226 -26373
rect 1826 -26443 2226 -26433
rect 2282 -26023 2682 -26013
rect 2282 -26083 2292 -26023
rect 2352 -26073 2612 -26023
rect 2352 -26083 2362 -26073
rect 2282 -26093 2362 -26083
rect 2602 -26083 2612 -26073
rect 2672 -26083 2682 -26023
rect 2602 -26093 2682 -26083
rect 2282 -26363 2342 -26093
rect 2422 -26153 2452 -26133
rect 2402 -26193 2452 -26153
rect 2512 -26153 2542 -26133
rect 2512 -26193 2562 -26153
rect 2402 -26263 2562 -26193
rect 2402 -26303 2452 -26263
rect 2422 -26323 2452 -26303
rect 2512 -26303 2562 -26263
rect 2512 -26323 2542 -26303
rect 2622 -26353 2682 -26093
rect 2612 -26363 2682 -26353
rect 2282 -26373 2362 -26363
rect 2282 -26433 2292 -26373
rect 2352 -26383 2362 -26373
rect 2602 -26373 2682 -26363
rect 2602 -26383 2612 -26373
rect 2352 -26433 2612 -26383
rect 2672 -26433 2682 -26373
rect 2282 -26443 2682 -26433
rect 2740 -26023 3140 -26013
rect 2740 -26083 2750 -26023
rect 2810 -26073 3070 -26023
rect 2810 -26083 2820 -26073
rect 2740 -26093 2820 -26083
rect 3060 -26083 3070 -26073
rect 3130 -26083 3140 -26023
rect 3060 -26093 3140 -26083
rect 2740 -26363 2800 -26093
rect 2880 -26153 2910 -26133
rect 2860 -26193 2910 -26153
rect 2970 -26153 3000 -26133
rect 2970 -26193 3020 -26153
rect 2860 -26263 3020 -26193
rect 2860 -26303 2910 -26263
rect 2880 -26323 2910 -26303
rect 2970 -26303 3020 -26263
rect 2970 -26323 3000 -26303
rect 3080 -26353 3140 -26093
rect 3070 -26363 3140 -26353
rect 2740 -26373 2820 -26363
rect 2740 -26433 2750 -26373
rect 2810 -26383 2820 -26373
rect 3060 -26373 3140 -26363
rect 3060 -26383 3070 -26373
rect 2810 -26433 3070 -26383
rect 3130 -26433 3140 -26373
rect 2740 -26443 3140 -26433
rect 3196 -26023 3596 -26013
rect 3196 -26083 3206 -26023
rect 3266 -26073 3526 -26023
rect 3266 -26083 3276 -26073
rect 3196 -26093 3276 -26083
rect 3516 -26083 3526 -26073
rect 3586 -26083 3596 -26023
rect 3516 -26093 3596 -26083
rect 3196 -26363 3256 -26093
rect 3336 -26153 3366 -26133
rect 3316 -26193 3366 -26153
rect 3426 -26153 3456 -26133
rect 3426 -26193 3476 -26153
rect 3316 -26263 3476 -26193
rect 3316 -26303 3366 -26263
rect 3336 -26323 3366 -26303
rect 3426 -26303 3476 -26263
rect 3426 -26323 3456 -26303
rect 3536 -26353 3596 -26093
rect 3526 -26363 3596 -26353
rect 3196 -26373 3276 -26363
rect 3196 -26433 3206 -26373
rect 3266 -26383 3276 -26373
rect 3516 -26373 3596 -26363
rect 3516 -26383 3526 -26373
rect 3266 -26433 3526 -26383
rect 3586 -26433 3596 -26373
rect 3196 -26443 3596 -26433
rect 3652 -26023 4052 -26013
rect 3652 -26083 3662 -26023
rect 3722 -26073 3982 -26023
rect 3722 -26083 3732 -26073
rect 3652 -26093 3732 -26083
rect 3972 -26083 3982 -26073
rect 4042 -26083 4052 -26023
rect 3972 -26093 4052 -26083
rect 3652 -26363 3712 -26093
rect 3792 -26153 3822 -26133
rect 3772 -26193 3822 -26153
rect 3882 -26153 3912 -26133
rect 3882 -26193 3932 -26153
rect 3772 -26263 3932 -26193
rect 3772 -26303 3822 -26263
rect 3792 -26323 3822 -26303
rect 3882 -26303 3932 -26263
rect 3882 -26323 3912 -26303
rect 3992 -26353 4052 -26093
rect 3982 -26363 4052 -26353
rect 3652 -26373 3732 -26363
rect 3652 -26433 3662 -26373
rect 3722 -26383 3732 -26373
rect 3972 -26373 4052 -26363
rect 3972 -26383 3982 -26373
rect 3722 -26433 3982 -26383
rect 4042 -26433 4052 -26373
rect 3652 -26443 4052 -26433
rect 4110 -26023 4510 -26013
rect 4110 -26083 4120 -26023
rect 4180 -26073 4440 -26023
rect 4180 -26083 4190 -26073
rect 4110 -26093 4190 -26083
rect 4430 -26083 4440 -26073
rect 4500 -26083 4510 -26023
rect 4430 -26093 4510 -26083
rect 4110 -26363 4170 -26093
rect 4250 -26153 4280 -26133
rect 4230 -26193 4280 -26153
rect 4340 -26153 4370 -26133
rect 4340 -26193 4390 -26153
rect 4230 -26263 4390 -26193
rect 4230 -26303 4280 -26263
rect 4250 -26323 4280 -26303
rect 4340 -26303 4390 -26263
rect 4340 -26323 4370 -26303
rect 4450 -26353 4510 -26093
rect 4440 -26363 4510 -26353
rect 4110 -26373 4190 -26363
rect 4110 -26433 4120 -26373
rect 4180 -26383 4190 -26373
rect 4430 -26373 4510 -26363
rect 4430 -26383 4440 -26373
rect 4180 -26433 4440 -26383
rect 4500 -26433 4510 -26373
rect 4110 -26443 4510 -26433
rect 4566 -26023 4966 -26013
rect 4566 -26083 4576 -26023
rect 4636 -26073 4896 -26023
rect 4636 -26083 4646 -26073
rect 4566 -26093 4646 -26083
rect 4886 -26083 4896 -26073
rect 4956 -26083 4966 -26023
rect 4886 -26093 4966 -26083
rect 4566 -26363 4626 -26093
rect 4706 -26153 4736 -26133
rect 4686 -26193 4736 -26153
rect 4796 -26153 4826 -26133
rect 4796 -26193 4846 -26153
rect 4686 -26263 4846 -26193
rect 4686 -26303 4736 -26263
rect 4706 -26323 4736 -26303
rect 4796 -26303 4846 -26263
rect 4796 -26323 4826 -26303
rect 4906 -26353 4966 -26093
rect 4896 -26363 4966 -26353
rect 4566 -26373 4646 -26363
rect 4566 -26433 4576 -26373
rect 4636 -26383 4646 -26373
rect 4886 -26373 4966 -26363
rect 4886 -26383 4896 -26373
rect 4636 -26433 4896 -26383
rect 4956 -26433 4966 -26373
rect 4566 -26443 4966 -26433
rect 5022 -26023 5422 -26013
rect 5022 -26083 5032 -26023
rect 5092 -26073 5352 -26023
rect 5092 -26083 5102 -26073
rect 5022 -26093 5102 -26083
rect 5342 -26083 5352 -26073
rect 5412 -26083 5422 -26023
rect 5342 -26093 5422 -26083
rect 5022 -26363 5082 -26093
rect 5162 -26153 5192 -26133
rect 5142 -26193 5192 -26153
rect 5252 -26153 5282 -26133
rect 5252 -26193 5302 -26153
rect 5142 -26263 5302 -26193
rect 5142 -26303 5192 -26263
rect 5162 -26323 5192 -26303
rect 5252 -26303 5302 -26263
rect 5252 -26323 5282 -26303
rect 5362 -26353 5422 -26093
rect 5352 -26363 5422 -26353
rect 5022 -26373 5102 -26363
rect 5022 -26433 5032 -26373
rect 5092 -26383 5102 -26373
rect 5342 -26373 5422 -26363
rect 5342 -26383 5352 -26373
rect 5092 -26433 5352 -26383
rect 5412 -26433 5422 -26373
rect 5022 -26443 5422 -26433
rect 5480 -26023 5880 -26013
rect 5480 -26083 5490 -26023
rect 5550 -26073 5810 -26023
rect 5550 -26083 5560 -26073
rect 5480 -26093 5560 -26083
rect 5800 -26083 5810 -26073
rect 5870 -26083 5880 -26023
rect 5800 -26093 5880 -26083
rect 5480 -26363 5540 -26093
rect 5620 -26153 5650 -26133
rect 5600 -26193 5650 -26153
rect 5710 -26153 5740 -26133
rect 5710 -26193 5760 -26153
rect 5600 -26263 5760 -26193
rect 5600 -26303 5650 -26263
rect 5620 -26323 5650 -26303
rect 5710 -26303 5760 -26263
rect 5710 -26323 5740 -26303
rect 5820 -26353 5880 -26093
rect 5810 -26363 5880 -26353
rect 5480 -26373 5560 -26363
rect 5480 -26433 5490 -26373
rect 5550 -26383 5560 -26373
rect 5800 -26373 5880 -26363
rect 5800 -26383 5810 -26373
rect 5550 -26433 5810 -26383
rect 5870 -26433 5880 -26373
rect 5480 -26443 5880 -26433
rect 5936 -26023 6336 -26013
rect 5936 -26083 5946 -26023
rect 6006 -26073 6266 -26023
rect 6006 -26083 6016 -26073
rect 5936 -26093 6016 -26083
rect 6256 -26083 6266 -26073
rect 6326 -26083 6336 -26023
rect 6256 -26093 6336 -26083
rect 5936 -26363 5996 -26093
rect 6076 -26153 6106 -26133
rect 6056 -26193 6106 -26153
rect 6166 -26153 6196 -26133
rect 6166 -26193 6216 -26153
rect 6056 -26263 6216 -26193
rect 6056 -26303 6106 -26263
rect 6076 -26323 6106 -26303
rect 6166 -26303 6216 -26263
rect 6166 -26323 6196 -26303
rect 6276 -26353 6336 -26093
rect 6266 -26363 6336 -26353
rect 5936 -26373 6016 -26363
rect 5936 -26433 5946 -26373
rect 6006 -26383 6016 -26373
rect 6256 -26373 6336 -26363
rect 6256 -26383 6266 -26373
rect 6006 -26433 6266 -26383
rect 6326 -26433 6336 -26373
rect 5936 -26443 6336 -26433
rect 6392 -26023 6792 -26013
rect 6392 -26083 6402 -26023
rect 6462 -26073 6722 -26023
rect 6462 -26083 6472 -26073
rect 6392 -26093 6472 -26083
rect 6712 -26083 6722 -26073
rect 6782 -26083 6792 -26023
rect 6712 -26093 6792 -26083
rect 6392 -26363 6452 -26093
rect 6532 -26153 6562 -26133
rect 6512 -26193 6562 -26153
rect 6622 -26153 6652 -26133
rect 6622 -26193 6672 -26153
rect 6512 -26263 6672 -26193
rect 6512 -26303 6562 -26263
rect 6532 -26323 6562 -26303
rect 6622 -26303 6672 -26263
rect 6622 -26323 6652 -26303
rect 6732 -26353 6792 -26093
rect 6722 -26363 6792 -26353
rect 6392 -26373 6472 -26363
rect 6392 -26433 6402 -26373
rect 6462 -26383 6472 -26373
rect 6712 -26373 6792 -26363
rect 6712 -26383 6722 -26373
rect 6462 -26433 6722 -26383
rect 6782 -26433 6792 -26373
rect 6392 -26443 6792 -26433
rect 6850 -26023 7250 -26013
rect 6850 -26083 6860 -26023
rect 6920 -26073 7180 -26023
rect 6920 -26083 6930 -26073
rect 6850 -26093 6930 -26083
rect 7170 -26083 7180 -26073
rect 7240 -26083 7250 -26023
rect 7170 -26093 7250 -26083
rect 6850 -26363 6910 -26093
rect 6990 -26153 7020 -26133
rect 6970 -26193 7020 -26153
rect 7080 -26153 7110 -26133
rect 7080 -26193 7130 -26153
rect 6970 -26263 7130 -26193
rect 6970 -26303 7020 -26263
rect 6990 -26323 7020 -26303
rect 7080 -26303 7130 -26263
rect 7080 -26323 7110 -26303
rect 7190 -26353 7250 -26093
rect 7180 -26363 7250 -26353
rect 6850 -26373 6930 -26363
rect 6850 -26433 6860 -26373
rect 6920 -26383 6930 -26373
rect 7170 -26373 7250 -26363
rect 7170 -26383 7180 -26373
rect 6920 -26433 7180 -26383
rect 7240 -26433 7250 -26373
rect 6850 -26443 7250 -26433
rect 7306 -26023 7706 -26013
rect 7306 -26083 7316 -26023
rect 7376 -26073 7636 -26023
rect 7376 -26083 7386 -26073
rect 7306 -26093 7386 -26083
rect 7626 -26083 7636 -26073
rect 7696 -26083 7706 -26023
rect 7626 -26093 7706 -26083
rect 7306 -26363 7366 -26093
rect 7446 -26153 7476 -26133
rect 7426 -26193 7476 -26153
rect 7536 -26153 7566 -26133
rect 7536 -26193 7586 -26153
rect 7426 -26263 7586 -26193
rect 7426 -26303 7476 -26263
rect 7446 -26323 7476 -26303
rect 7536 -26303 7586 -26263
rect 7536 -26323 7566 -26303
rect 7646 -26353 7706 -26093
rect 7636 -26363 7706 -26353
rect 7306 -26373 7386 -26363
rect 7306 -26433 7316 -26373
rect 7376 -26383 7386 -26373
rect 7626 -26373 7706 -26363
rect 7626 -26383 7636 -26373
rect 7376 -26433 7636 -26383
rect 7696 -26433 7706 -26373
rect 7306 -26443 7706 -26433
rect 7762 -26023 8162 -26013
rect 7762 -26083 7772 -26023
rect 7832 -26073 8092 -26023
rect 7832 -26083 7842 -26073
rect 7762 -26093 7842 -26083
rect 8082 -26083 8092 -26073
rect 8152 -26083 8162 -26023
rect 8082 -26093 8162 -26083
rect 7762 -26363 7822 -26093
rect 7902 -26153 7932 -26133
rect 7882 -26193 7932 -26153
rect 7992 -26153 8022 -26133
rect 7992 -26193 8042 -26153
rect 7882 -26263 8042 -26193
rect 7882 -26303 7932 -26263
rect 7902 -26323 7932 -26303
rect 7992 -26303 8042 -26263
rect 7992 -26323 8022 -26303
rect 8102 -26353 8162 -26093
rect 8092 -26363 8162 -26353
rect 7762 -26373 7842 -26363
rect 7762 -26433 7772 -26373
rect 7832 -26383 7842 -26373
rect 8082 -26373 8162 -26363
rect 8082 -26383 8092 -26373
rect 7832 -26433 8092 -26383
rect 8152 -26433 8162 -26373
rect 7762 -26443 8162 -26433
rect 8236 -26023 8636 -26013
rect 8236 -26083 8246 -26023
rect 8306 -26073 8566 -26023
rect 8306 -26083 8316 -26073
rect 8236 -26093 8316 -26083
rect 8556 -26083 8566 -26073
rect 8626 -26083 8636 -26023
rect 8556 -26093 8636 -26083
rect 8236 -26363 8296 -26093
rect 8376 -26153 8406 -26133
rect 8356 -26193 8406 -26153
rect 8466 -26153 8496 -26133
rect 8466 -26193 8516 -26153
rect 8356 -26263 8516 -26193
rect 8356 -26303 8406 -26263
rect 8376 -26323 8406 -26303
rect 8466 -26303 8516 -26263
rect 8466 -26323 8496 -26303
rect 8576 -26353 8636 -26093
rect 8566 -26363 8636 -26353
rect 8236 -26373 8316 -26363
rect 8236 -26433 8246 -26373
rect 8306 -26383 8316 -26373
rect 8556 -26373 8636 -26363
rect 8556 -26383 8566 -26373
rect 8306 -26433 8566 -26383
rect 8626 -26433 8636 -26373
rect 8236 -26443 8636 -26433
rect 8692 -26023 9092 -26013
rect 8692 -26083 8702 -26023
rect 8762 -26073 9022 -26023
rect 8762 -26083 8772 -26073
rect 8692 -26093 8772 -26083
rect 9012 -26083 9022 -26073
rect 9082 -26083 9092 -26023
rect 9012 -26093 9092 -26083
rect 8692 -26363 8752 -26093
rect 8832 -26153 8862 -26133
rect 8812 -26193 8862 -26153
rect 8922 -26153 8952 -26133
rect 8922 -26193 8972 -26153
rect 8812 -26263 8972 -26193
rect 8812 -26303 8862 -26263
rect 8832 -26323 8862 -26303
rect 8922 -26303 8972 -26263
rect 8922 -26323 8952 -26303
rect 9032 -26353 9092 -26093
rect 9022 -26363 9092 -26353
rect 8692 -26373 8772 -26363
rect 8692 -26433 8702 -26373
rect 8762 -26383 8772 -26373
rect 9012 -26373 9092 -26363
rect 9012 -26383 9022 -26373
rect 8762 -26433 9022 -26383
rect 9082 -26433 9092 -26373
rect 8692 -26443 9092 -26433
rect 9150 -26023 9550 -26013
rect 9150 -26083 9160 -26023
rect 9220 -26073 9480 -26023
rect 9220 -26083 9230 -26073
rect 9150 -26093 9230 -26083
rect 9470 -26083 9480 -26073
rect 9540 -26083 9550 -26023
rect 9470 -26093 9550 -26083
rect 9150 -26363 9210 -26093
rect 9290 -26153 9320 -26133
rect 9270 -26193 9320 -26153
rect 9380 -26153 9410 -26133
rect 9380 -26193 9430 -26153
rect 9270 -26263 9430 -26193
rect 9270 -26303 9320 -26263
rect 9290 -26323 9320 -26303
rect 9380 -26303 9430 -26263
rect 9380 -26323 9410 -26303
rect 9490 -26353 9550 -26093
rect 9480 -26363 9550 -26353
rect 9150 -26373 9230 -26363
rect 9150 -26433 9160 -26373
rect 9220 -26383 9230 -26373
rect 9470 -26373 9550 -26363
rect 9470 -26383 9480 -26373
rect 9220 -26433 9480 -26383
rect 9540 -26433 9550 -26373
rect 9150 -26443 9550 -26433
rect 9606 -26023 10006 -26013
rect 9606 -26083 9616 -26023
rect 9676 -26073 9936 -26023
rect 9676 -26083 9686 -26073
rect 9606 -26093 9686 -26083
rect 9926 -26083 9936 -26073
rect 9996 -26083 10006 -26023
rect 9926 -26093 10006 -26083
rect 9606 -26363 9666 -26093
rect 9746 -26153 9776 -26133
rect 9726 -26193 9776 -26153
rect 9836 -26153 9866 -26133
rect 9836 -26193 9886 -26153
rect 9726 -26263 9886 -26193
rect 9726 -26303 9776 -26263
rect 9746 -26323 9776 -26303
rect 9836 -26303 9886 -26263
rect 9836 -26323 9866 -26303
rect 9946 -26353 10006 -26093
rect 9936 -26363 10006 -26353
rect 9606 -26373 9686 -26363
rect 9606 -26433 9616 -26373
rect 9676 -26383 9686 -26373
rect 9926 -26373 10006 -26363
rect 9926 -26383 9936 -26373
rect 9676 -26433 9936 -26383
rect 9996 -26433 10006 -26373
rect 9606 -26443 10006 -26433
rect 10062 -26023 10462 -26013
rect 10062 -26083 10072 -26023
rect 10132 -26073 10392 -26023
rect 10132 -26083 10142 -26073
rect 10062 -26093 10142 -26083
rect 10382 -26083 10392 -26073
rect 10452 -26083 10462 -26023
rect 10382 -26093 10462 -26083
rect 10062 -26363 10122 -26093
rect 10202 -26153 10232 -26133
rect 10182 -26193 10232 -26153
rect 10292 -26153 10322 -26133
rect 10292 -26193 10342 -26153
rect 10182 -26263 10342 -26193
rect 10182 -26303 10232 -26263
rect 10202 -26323 10232 -26303
rect 10292 -26303 10342 -26263
rect 10292 -26323 10322 -26303
rect 10402 -26353 10462 -26093
rect 10392 -26363 10462 -26353
rect 10062 -26373 10142 -26363
rect 10062 -26433 10072 -26373
rect 10132 -26383 10142 -26373
rect 10382 -26373 10462 -26363
rect 10382 -26383 10392 -26373
rect 10132 -26433 10392 -26383
rect 10452 -26433 10462 -26373
rect 10062 -26443 10462 -26433
rect 10520 -26023 10920 -26013
rect 10520 -26083 10530 -26023
rect 10590 -26073 10850 -26023
rect 10590 -26083 10600 -26073
rect 10520 -26093 10600 -26083
rect 10840 -26083 10850 -26073
rect 10910 -26083 10920 -26023
rect 10840 -26093 10920 -26083
rect 10520 -26363 10580 -26093
rect 10660 -26153 10690 -26133
rect 10640 -26193 10690 -26153
rect 10750 -26153 10780 -26133
rect 10750 -26193 10800 -26153
rect 10640 -26263 10800 -26193
rect 10640 -26303 10690 -26263
rect 10660 -26323 10690 -26303
rect 10750 -26303 10800 -26263
rect 10750 -26323 10780 -26303
rect 10860 -26353 10920 -26093
rect 10850 -26363 10920 -26353
rect 10520 -26373 10600 -26363
rect 10520 -26433 10530 -26373
rect 10590 -26383 10600 -26373
rect 10840 -26373 10920 -26363
rect 10840 -26383 10850 -26373
rect 10590 -26433 10850 -26383
rect 10910 -26433 10920 -26373
rect 10520 -26443 10920 -26433
rect 10976 -26023 11376 -26013
rect 10976 -26083 10986 -26023
rect 11046 -26073 11306 -26023
rect 11046 -26083 11056 -26073
rect 10976 -26093 11056 -26083
rect 11296 -26083 11306 -26073
rect 11366 -26083 11376 -26023
rect 11296 -26093 11376 -26083
rect 10976 -26363 11036 -26093
rect 11116 -26153 11146 -26133
rect 11096 -26193 11146 -26153
rect 11206 -26153 11236 -26133
rect 11206 -26193 11256 -26153
rect 11096 -26263 11256 -26193
rect 11096 -26303 11146 -26263
rect 11116 -26323 11146 -26303
rect 11206 -26303 11256 -26263
rect 11206 -26323 11236 -26303
rect 11316 -26353 11376 -26093
rect 11306 -26363 11376 -26353
rect 10976 -26373 11056 -26363
rect 10976 -26433 10986 -26373
rect 11046 -26383 11056 -26373
rect 11296 -26373 11376 -26363
rect 11296 -26383 11306 -26373
rect 11046 -26433 11306 -26383
rect 11366 -26433 11376 -26373
rect 10976 -26443 11376 -26433
rect 11432 -26023 11832 -26013
rect 11432 -26083 11442 -26023
rect 11502 -26073 11762 -26023
rect 11502 -26083 11512 -26073
rect 11432 -26093 11512 -26083
rect 11752 -26083 11762 -26073
rect 11822 -26083 11832 -26023
rect 11752 -26093 11832 -26083
rect 11432 -26363 11492 -26093
rect 11572 -26153 11602 -26133
rect 11552 -26193 11602 -26153
rect 11662 -26153 11692 -26133
rect 11662 -26193 11712 -26153
rect 11552 -26263 11712 -26193
rect 11552 -26303 11602 -26263
rect 11572 -26323 11602 -26303
rect 11662 -26303 11712 -26263
rect 11662 -26323 11692 -26303
rect 11772 -26353 11832 -26093
rect 11762 -26363 11832 -26353
rect 11432 -26373 11512 -26363
rect 11432 -26433 11442 -26373
rect 11502 -26383 11512 -26373
rect 11752 -26373 11832 -26363
rect 11752 -26383 11762 -26373
rect 11502 -26433 11762 -26383
rect 11822 -26433 11832 -26373
rect 11432 -26443 11832 -26433
rect 11890 -26023 12290 -26013
rect 11890 -26083 11900 -26023
rect 11960 -26073 12220 -26023
rect 11960 -26083 11970 -26073
rect 11890 -26093 11970 -26083
rect 12210 -26083 12220 -26073
rect 12280 -26083 12290 -26023
rect 12210 -26093 12290 -26083
rect 11890 -26363 11950 -26093
rect 12030 -26153 12060 -26133
rect 12010 -26193 12060 -26153
rect 12120 -26153 12150 -26133
rect 12120 -26193 12170 -26153
rect 12010 -26263 12170 -26193
rect 12010 -26303 12060 -26263
rect 12030 -26323 12060 -26303
rect 12120 -26303 12170 -26263
rect 12120 -26323 12150 -26303
rect 12230 -26353 12290 -26093
rect 12220 -26363 12290 -26353
rect 11890 -26373 11970 -26363
rect 11890 -26433 11900 -26373
rect 11960 -26383 11970 -26373
rect 12210 -26373 12290 -26363
rect 12210 -26383 12220 -26373
rect 11960 -26433 12220 -26383
rect 12280 -26433 12290 -26373
rect 11890 -26443 12290 -26433
rect 12346 -26023 12746 -26013
rect 12346 -26083 12356 -26023
rect 12416 -26073 12676 -26023
rect 12416 -26083 12426 -26073
rect 12346 -26093 12426 -26083
rect 12666 -26083 12676 -26073
rect 12736 -26083 12746 -26023
rect 12666 -26093 12746 -26083
rect 12346 -26363 12406 -26093
rect 12486 -26153 12516 -26133
rect 12466 -26193 12516 -26153
rect 12576 -26153 12606 -26133
rect 12576 -26193 12626 -26153
rect 12466 -26263 12626 -26193
rect 12466 -26303 12516 -26263
rect 12486 -26323 12516 -26303
rect 12576 -26303 12626 -26263
rect 12576 -26323 12606 -26303
rect 12686 -26353 12746 -26093
rect 12676 -26363 12746 -26353
rect 12346 -26373 12426 -26363
rect 12346 -26433 12356 -26373
rect 12416 -26383 12426 -26373
rect 12666 -26373 12746 -26363
rect 12666 -26383 12676 -26373
rect 12416 -26433 12676 -26383
rect 12736 -26433 12746 -26373
rect 12346 -26443 12746 -26433
rect 12802 -26023 13202 -26013
rect 12802 -26083 12812 -26023
rect 12872 -26073 13132 -26023
rect 12872 -26083 12882 -26073
rect 12802 -26093 12882 -26083
rect 13122 -26083 13132 -26073
rect 13192 -26083 13202 -26023
rect 13122 -26093 13202 -26083
rect 12802 -26363 12862 -26093
rect 12942 -26153 12972 -26133
rect 12922 -26193 12972 -26153
rect 13032 -26153 13062 -26133
rect 13032 -26193 13082 -26153
rect 12922 -26263 13082 -26193
rect 12922 -26303 12972 -26263
rect 12942 -26323 12972 -26303
rect 13032 -26303 13082 -26263
rect 13032 -26323 13062 -26303
rect 13142 -26353 13202 -26093
rect 13132 -26363 13202 -26353
rect 12802 -26373 12882 -26363
rect 12802 -26433 12812 -26373
rect 12872 -26383 12882 -26373
rect 13122 -26373 13202 -26363
rect 13122 -26383 13132 -26373
rect 12872 -26433 13132 -26383
rect 13192 -26433 13202 -26373
rect 12802 -26443 13202 -26433
rect 13260 -26023 13660 -26013
rect 13260 -26083 13270 -26023
rect 13330 -26073 13590 -26023
rect 13330 -26083 13340 -26073
rect 13260 -26093 13340 -26083
rect 13580 -26083 13590 -26073
rect 13650 -26083 13660 -26023
rect 13580 -26093 13660 -26083
rect 13260 -26363 13320 -26093
rect 13400 -26153 13430 -26133
rect 13380 -26193 13430 -26153
rect 13490 -26153 13520 -26133
rect 13490 -26193 13540 -26153
rect 13380 -26263 13540 -26193
rect 13380 -26303 13430 -26263
rect 13400 -26323 13430 -26303
rect 13490 -26303 13540 -26263
rect 13490 -26323 13520 -26303
rect 13600 -26353 13660 -26093
rect 13590 -26363 13660 -26353
rect 13260 -26373 13340 -26363
rect 13260 -26433 13270 -26373
rect 13330 -26383 13340 -26373
rect 13580 -26373 13660 -26363
rect 13580 -26383 13590 -26373
rect 13330 -26433 13590 -26383
rect 13650 -26433 13660 -26373
rect 13260 -26443 13660 -26433
rect 13716 -26023 14116 -26013
rect 13716 -26083 13726 -26023
rect 13786 -26073 14046 -26023
rect 13786 -26083 13796 -26073
rect 13716 -26093 13796 -26083
rect 14036 -26083 14046 -26073
rect 14106 -26083 14116 -26023
rect 14036 -26093 14116 -26083
rect 13716 -26363 13776 -26093
rect 13856 -26153 13886 -26133
rect 13836 -26193 13886 -26153
rect 13946 -26153 13976 -26133
rect 13946 -26193 13996 -26153
rect 13836 -26263 13996 -26193
rect 13836 -26303 13886 -26263
rect 13856 -26323 13886 -26303
rect 13946 -26303 13996 -26263
rect 13946 -26323 13976 -26303
rect 14056 -26353 14116 -26093
rect 14046 -26363 14116 -26353
rect 13716 -26373 13796 -26363
rect 13716 -26433 13726 -26373
rect 13786 -26383 13796 -26373
rect 14036 -26373 14116 -26363
rect 14036 -26383 14046 -26373
rect 13786 -26433 14046 -26383
rect 14106 -26433 14116 -26373
rect 13716 -26443 14116 -26433
rect 14172 -26023 14572 -26013
rect 14172 -26083 14182 -26023
rect 14242 -26073 14502 -26023
rect 14242 -26083 14252 -26073
rect 14172 -26093 14252 -26083
rect 14492 -26083 14502 -26073
rect 14562 -26083 14572 -26023
rect 14492 -26093 14572 -26083
rect 14172 -26363 14232 -26093
rect 14312 -26153 14342 -26133
rect 14292 -26193 14342 -26153
rect 14402 -26153 14432 -26133
rect 14402 -26193 14452 -26153
rect 14292 -26263 14452 -26193
rect 14292 -26303 14342 -26263
rect 14312 -26323 14342 -26303
rect 14402 -26303 14452 -26263
rect 14402 -26323 14432 -26303
rect 14512 -26353 14572 -26093
rect 14502 -26363 14572 -26353
rect 14172 -26373 14252 -26363
rect 14172 -26433 14182 -26373
rect 14242 -26383 14252 -26373
rect 14492 -26373 14572 -26363
rect 14492 -26383 14502 -26373
rect 14242 -26433 14502 -26383
rect 14562 -26433 14572 -26373
rect 14172 -26443 14572 -26433
rect 14630 -26023 15030 -26013
rect 14630 -26083 14640 -26023
rect 14700 -26073 14960 -26023
rect 14700 -26083 14710 -26073
rect 14630 -26093 14710 -26083
rect 14950 -26083 14960 -26073
rect 15020 -26083 15030 -26023
rect 14950 -26093 15030 -26083
rect 14630 -26363 14690 -26093
rect 14770 -26153 14800 -26133
rect 14750 -26193 14800 -26153
rect 14860 -26153 14890 -26133
rect 14860 -26193 14910 -26153
rect 14750 -26263 14910 -26193
rect 14750 -26303 14800 -26263
rect 14770 -26323 14800 -26303
rect 14860 -26303 14910 -26263
rect 14860 -26323 14890 -26303
rect 14970 -26353 15030 -26093
rect 14960 -26363 15030 -26353
rect 14630 -26373 14710 -26363
rect 14630 -26433 14640 -26373
rect 14700 -26383 14710 -26373
rect 14950 -26373 15030 -26363
rect 14950 -26383 14960 -26373
rect 14700 -26433 14960 -26383
rect 15020 -26433 15030 -26373
rect 14630 -26443 15030 -26433
rect 15086 -26023 15486 -26013
rect 15086 -26083 15096 -26023
rect 15156 -26073 15416 -26023
rect 15156 -26083 15166 -26073
rect 15086 -26093 15166 -26083
rect 15406 -26083 15416 -26073
rect 15476 -26083 15486 -26023
rect 15406 -26093 15486 -26083
rect 15086 -26363 15146 -26093
rect 15226 -26153 15256 -26133
rect 15206 -26193 15256 -26153
rect 15316 -26153 15346 -26133
rect 15316 -26193 15366 -26153
rect 15206 -26263 15366 -26193
rect 15206 -26303 15256 -26263
rect 15226 -26323 15256 -26303
rect 15316 -26303 15366 -26263
rect 15316 -26323 15346 -26303
rect 15426 -26353 15486 -26093
rect 15416 -26363 15486 -26353
rect 15086 -26373 15166 -26363
rect 15086 -26433 15096 -26373
rect 15156 -26383 15166 -26373
rect 15406 -26373 15486 -26363
rect 15406 -26383 15416 -26373
rect 15156 -26433 15416 -26383
rect 15476 -26433 15486 -26373
rect 15086 -26443 15486 -26433
rect 0 -26515 400 -26505
rect 0 -26575 10 -26515
rect 70 -26565 330 -26515
rect 70 -26575 80 -26565
rect 0 -26585 80 -26575
rect 320 -26575 330 -26565
rect 390 -26575 400 -26515
rect 320 -26585 400 -26575
rect 0 -26855 60 -26585
rect 140 -26645 170 -26625
rect 120 -26685 170 -26645
rect 230 -26645 260 -26625
rect 230 -26685 280 -26645
rect 120 -26755 280 -26685
rect 120 -26795 170 -26755
rect 140 -26815 170 -26795
rect 230 -26795 280 -26755
rect 230 -26815 260 -26795
rect 340 -26845 400 -26585
rect 330 -26855 400 -26845
rect 0 -26865 80 -26855
rect 0 -26925 10 -26865
rect 70 -26875 80 -26865
rect 320 -26865 400 -26855
rect 320 -26875 330 -26865
rect 70 -26925 330 -26875
rect 390 -26925 400 -26865
rect 0 -26935 400 -26925
rect 456 -26515 856 -26505
rect 456 -26575 466 -26515
rect 526 -26565 786 -26515
rect 526 -26575 536 -26565
rect 456 -26585 536 -26575
rect 776 -26575 786 -26565
rect 846 -26575 856 -26515
rect 776 -26585 856 -26575
rect 456 -26855 516 -26585
rect 596 -26645 626 -26625
rect 576 -26685 626 -26645
rect 686 -26645 716 -26625
rect 686 -26685 736 -26645
rect 576 -26755 736 -26685
rect 576 -26795 626 -26755
rect 596 -26815 626 -26795
rect 686 -26795 736 -26755
rect 686 -26815 716 -26795
rect 796 -26845 856 -26585
rect 786 -26855 856 -26845
rect 456 -26865 536 -26855
rect 456 -26925 466 -26865
rect 526 -26875 536 -26865
rect 776 -26865 856 -26855
rect 776 -26875 786 -26865
rect 526 -26925 786 -26875
rect 846 -26925 856 -26865
rect 456 -26935 856 -26925
rect 912 -26515 1312 -26505
rect 912 -26575 922 -26515
rect 982 -26565 1242 -26515
rect 982 -26575 992 -26565
rect 912 -26585 992 -26575
rect 1232 -26575 1242 -26565
rect 1302 -26575 1312 -26515
rect 1232 -26585 1312 -26575
rect 912 -26855 972 -26585
rect 1052 -26645 1082 -26625
rect 1032 -26685 1082 -26645
rect 1142 -26645 1172 -26625
rect 1142 -26685 1192 -26645
rect 1032 -26755 1192 -26685
rect 1032 -26795 1082 -26755
rect 1052 -26815 1082 -26795
rect 1142 -26795 1192 -26755
rect 1142 -26815 1172 -26795
rect 1252 -26845 1312 -26585
rect 1242 -26855 1312 -26845
rect 912 -26865 992 -26855
rect 912 -26925 922 -26865
rect 982 -26875 992 -26865
rect 1232 -26865 1312 -26855
rect 1232 -26875 1242 -26865
rect 982 -26925 1242 -26875
rect 1302 -26925 1312 -26865
rect 912 -26935 1312 -26925
rect 1370 -26515 1770 -26505
rect 1370 -26575 1380 -26515
rect 1440 -26565 1700 -26515
rect 1440 -26575 1450 -26565
rect 1370 -26585 1450 -26575
rect 1690 -26575 1700 -26565
rect 1760 -26575 1770 -26515
rect 1690 -26585 1770 -26575
rect 1370 -26855 1430 -26585
rect 1510 -26645 1540 -26625
rect 1490 -26685 1540 -26645
rect 1600 -26645 1630 -26625
rect 1600 -26685 1650 -26645
rect 1490 -26755 1650 -26685
rect 1490 -26795 1540 -26755
rect 1510 -26815 1540 -26795
rect 1600 -26795 1650 -26755
rect 1600 -26815 1630 -26795
rect 1710 -26845 1770 -26585
rect 1700 -26855 1770 -26845
rect 1370 -26865 1450 -26855
rect 1370 -26925 1380 -26865
rect 1440 -26875 1450 -26865
rect 1690 -26865 1770 -26855
rect 1690 -26875 1700 -26865
rect 1440 -26925 1700 -26875
rect 1760 -26925 1770 -26865
rect 1370 -26935 1770 -26925
rect 1826 -26515 2226 -26505
rect 1826 -26575 1836 -26515
rect 1896 -26565 2156 -26515
rect 1896 -26575 1906 -26565
rect 1826 -26585 1906 -26575
rect 2146 -26575 2156 -26565
rect 2216 -26575 2226 -26515
rect 2146 -26585 2226 -26575
rect 1826 -26855 1886 -26585
rect 1966 -26645 1996 -26625
rect 1946 -26685 1996 -26645
rect 2056 -26645 2086 -26625
rect 2056 -26685 2106 -26645
rect 1946 -26755 2106 -26685
rect 1946 -26795 1996 -26755
rect 1966 -26815 1996 -26795
rect 2056 -26795 2106 -26755
rect 2056 -26815 2086 -26795
rect 2166 -26845 2226 -26585
rect 2156 -26855 2226 -26845
rect 1826 -26865 1906 -26855
rect 1826 -26925 1836 -26865
rect 1896 -26875 1906 -26865
rect 2146 -26865 2226 -26855
rect 2146 -26875 2156 -26865
rect 1896 -26925 2156 -26875
rect 2216 -26925 2226 -26865
rect 1826 -26935 2226 -26925
rect 2282 -26515 2682 -26505
rect 2282 -26575 2292 -26515
rect 2352 -26565 2612 -26515
rect 2352 -26575 2362 -26565
rect 2282 -26585 2362 -26575
rect 2602 -26575 2612 -26565
rect 2672 -26575 2682 -26515
rect 2602 -26585 2682 -26575
rect 2282 -26855 2342 -26585
rect 2422 -26645 2452 -26625
rect 2402 -26685 2452 -26645
rect 2512 -26645 2542 -26625
rect 2512 -26685 2562 -26645
rect 2402 -26755 2562 -26685
rect 2402 -26795 2452 -26755
rect 2422 -26815 2452 -26795
rect 2512 -26795 2562 -26755
rect 2512 -26815 2542 -26795
rect 2622 -26845 2682 -26585
rect 2612 -26855 2682 -26845
rect 2282 -26865 2362 -26855
rect 2282 -26925 2292 -26865
rect 2352 -26875 2362 -26865
rect 2602 -26865 2682 -26855
rect 2602 -26875 2612 -26865
rect 2352 -26925 2612 -26875
rect 2672 -26925 2682 -26865
rect 2282 -26935 2682 -26925
rect 2740 -26515 3140 -26505
rect 2740 -26575 2750 -26515
rect 2810 -26565 3070 -26515
rect 2810 -26575 2820 -26565
rect 2740 -26585 2820 -26575
rect 3060 -26575 3070 -26565
rect 3130 -26575 3140 -26515
rect 3060 -26585 3140 -26575
rect 2740 -26855 2800 -26585
rect 2880 -26645 2910 -26625
rect 2860 -26685 2910 -26645
rect 2970 -26645 3000 -26625
rect 2970 -26685 3020 -26645
rect 2860 -26755 3020 -26685
rect 2860 -26795 2910 -26755
rect 2880 -26815 2910 -26795
rect 2970 -26795 3020 -26755
rect 2970 -26815 3000 -26795
rect 3080 -26845 3140 -26585
rect 3070 -26855 3140 -26845
rect 2740 -26865 2820 -26855
rect 2740 -26925 2750 -26865
rect 2810 -26875 2820 -26865
rect 3060 -26865 3140 -26855
rect 3060 -26875 3070 -26865
rect 2810 -26925 3070 -26875
rect 3130 -26925 3140 -26865
rect 2740 -26935 3140 -26925
rect 3196 -26515 3596 -26505
rect 3196 -26575 3206 -26515
rect 3266 -26565 3526 -26515
rect 3266 -26575 3276 -26565
rect 3196 -26585 3276 -26575
rect 3516 -26575 3526 -26565
rect 3586 -26575 3596 -26515
rect 3516 -26585 3596 -26575
rect 3196 -26855 3256 -26585
rect 3336 -26645 3366 -26625
rect 3316 -26685 3366 -26645
rect 3426 -26645 3456 -26625
rect 3426 -26685 3476 -26645
rect 3316 -26755 3476 -26685
rect 3316 -26795 3366 -26755
rect 3336 -26815 3366 -26795
rect 3426 -26795 3476 -26755
rect 3426 -26815 3456 -26795
rect 3536 -26845 3596 -26585
rect 3526 -26855 3596 -26845
rect 3196 -26865 3276 -26855
rect 3196 -26925 3206 -26865
rect 3266 -26875 3276 -26865
rect 3516 -26865 3596 -26855
rect 3516 -26875 3526 -26865
rect 3266 -26925 3526 -26875
rect 3586 -26925 3596 -26865
rect 3196 -26935 3596 -26925
rect 3652 -26515 4052 -26505
rect 3652 -26575 3662 -26515
rect 3722 -26565 3982 -26515
rect 3722 -26575 3732 -26565
rect 3652 -26585 3732 -26575
rect 3972 -26575 3982 -26565
rect 4042 -26575 4052 -26515
rect 3972 -26585 4052 -26575
rect 3652 -26855 3712 -26585
rect 3792 -26645 3822 -26625
rect 3772 -26685 3822 -26645
rect 3882 -26645 3912 -26625
rect 3882 -26685 3932 -26645
rect 3772 -26755 3932 -26685
rect 3772 -26795 3822 -26755
rect 3792 -26815 3822 -26795
rect 3882 -26795 3932 -26755
rect 3882 -26815 3912 -26795
rect 3992 -26845 4052 -26585
rect 3982 -26855 4052 -26845
rect 3652 -26865 3732 -26855
rect 3652 -26925 3662 -26865
rect 3722 -26875 3732 -26865
rect 3972 -26865 4052 -26855
rect 3972 -26875 3982 -26865
rect 3722 -26925 3982 -26875
rect 4042 -26925 4052 -26865
rect 3652 -26935 4052 -26925
rect 4110 -26515 4510 -26505
rect 4110 -26575 4120 -26515
rect 4180 -26565 4440 -26515
rect 4180 -26575 4190 -26565
rect 4110 -26585 4190 -26575
rect 4430 -26575 4440 -26565
rect 4500 -26575 4510 -26515
rect 4430 -26585 4510 -26575
rect 4110 -26855 4170 -26585
rect 4250 -26645 4280 -26625
rect 4230 -26685 4280 -26645
rect 4340 -26645 4370 -26625
rect 4340 -26685 4390 -26645
rect 4230 -26755 4390 -26685
rect 4230 -26795 4280 -26755
rect 4250 -26815 4280 -26795
rect 4340 -26795 4390 -26755
rect 4340 -26815 4370 -26795
rect 4450 -26845 4510 -26585
rect 4440 -26855 4510 -26845
rect 4110 -26865 4190 -26855
rect 4110 -26925 4120 -26865
rect 4180 -26875 4190 -26865
rect 4430 -26865 4510 -26855
rect 4430 -26875 4440 -26865
rect 4180 -26925 4440 -26875
rect 4500 -26925 4510 -26865
rect 4110 -26935 4510 -26925
rect 4566 -26515 4966 -26505
rect 4566 -26575 4576 -26515
rect 4636 -26565 4896 -26515
rect 4636 -26575 4646 -26565
rect 4566 -26585 4646 -26575
rect 4886 -26575 4896 -26565
rect 4956 -26575 4966 -26515
rect 4886 -26585 4966 -26575
rect 4566 -26855 4626 -26585
rect 4706 -26645 4736 -26625
rect 4686 -26685 4736 -26645
rect 4796 -26645 4826 -26625
rect 4796 -26685 4846 -26645
rect 4686 -26755 4846 -26685
rect 4686 -26795 4736 -26755
rect 4706 -26815 4736 -26795
rect 4796 -26795 4846 -26755
rect 4796 -26815 4826 -26795
rect 4906 -26845 4966 -26585
rect 4896 -26855 4966 -26845
rect 4566 -26865 4646 -26855
rect 4566 -26925 4576 -26865
rect 4636 -26875 4646 -26865
rect 4886 -26865 4966 -26855
rect 4886 -26875 4896 -26865
rect 4636 -26925 4896 -26875
rect 4956 -26925 4966 -26865
rect 4566 -26935 4966 -26925
rect 5022 -26515 5422 -26505
rect 5022 -26575 5032 -26515
rect 5092 -26565 5352 -26515
rect 5092 -26575 5102 -26565
rect 5022 -26585 5102 -26575
rect 5342 -26575 5352 -26565
rect 5412 -26575 5422 -26515
rect 5342 -26585 5422 -26575
rect 5022 -26855 5082 -26585
rect 5162 -26645 5192 -26625
rect 5142 -26685 5192 -26645
rect 5252 -26645 5282 -26625
rect 5252 -26685 5302 -26645
rect 5142 -26755 5302 -26685
rect 5142 -26795 5192 -26755
rect 5162 -26815 5192 -26795
rect 5252 -26795 5302 -26755
rect 5252 -26815 5282 -26795
rect 5362 -26845 5422 -26585
rect 5352 -26855 5422 -26845
rect 5022 -26865 5102 -26855
rect 5022 -26925 5032 -26865
rect 5092 -26875 5102 -26865
rect 5342 -26865 5422 -26855
rect 5342 -26875 5352 -26865
rect 5092 -26925 5352 -26875
rect 5412 -26925 5422 -26865
rect 5022 -26935 5422 -26925
rect 5480 -26515 5880 -26505
rect 5480 -26575 5490 -26515
rect 5550 -26565 5810 -26515
rect 5550 -26575 5560 -26565
rect 5480 -26585 5560 -26575
rect 5800 -26575 5810 -26565
rect 5870 -26575 5880 -26515
rect 5800 -26585 5880 -26575
rect 5480 -26855 5540 -26585
rect 5620 -26645 5650 -26625
rect 5600 -26685 5650 -26645
rect 5710 -26645 5740 -26625
rect 5710 -26685 5760 -26645
rect 5600 -26755 5760 -26685
rect 5600 -26795 5650 -26755
rect 5620 -26815 5650 -26795
rect 5710 -26795 5760 -26755
rect 5710 -26815 5740 -26795
rect 5820 -26845 5880 -26585
rect 5810 -26855 5880 -26845
rect 5480 -26865 5560 -26855
rect 5480 -26925 5490 -26865
rect 5550 -26875 5560 -26865
rect 5800 -26865 5880 -26855
rect 5800 -26875 5810 -26865
rect 5550 -26925 5810 -26875
rect 5870 -26925 5880 -26865
rect 5480 -26935 5880 -26925
rect 5936 -26515 6336 -26505
rect 5936 -26575 5946 -26515
rect 6006 -26565 6266 -26515
rect 6006 -26575 6016 -26565
rect 5936 -26585 6016 -26575
rect 6256 -26575 6266 -26565
rect 6326 -26575 6336 -26515
rect 6256 -26585 6336 -26575
rect 5936 -26855 5996 -26585
rect 6076 -26645 6106 -26625
rect 6056 -26685 6106 -26645
rect 6166 -26645 6196 -26625
rect 6166 -26685 6216 -26645
rect 6056 -26755 6216 -26685
rect 6056 -26795 6106 -26755
rect 6076 -26815 6106 -26795
rect 6166 -26795 6216 -26755
rect 6166 -26815 6196 -26795
rect 6276 -26845 6336 -26585
rect 6266 -26855 6336 -26845
rect 5936 -26865 6016 -26855
rect 5936 -26925 5946 -26865
rect 6006 -26875 6016 -26865
rect 6256 -26865 6336 -26855
rect 6256 -26875 6266 -26865
rect 6006 -26925 6266 -26875
rect 6326 -26925 6336 -26865
rect 5936 -26935 6336 -26925
rect 6392 -26515 6792 -26505
rect 6392 -26575 6402 -26515
rect 6462 -26565 6722 -26515
rect 6462 -26575 6472 -26565
rect 6392 -26585 6472 -26575
rect 6712 -26575 6722 -26565
rect 6782 -26575 6792 -26515
rect 6712 -26585 6792 -26575
rect 6392 -26855 6452 -26585
rect 6532 -26645 6562 -26625
rect 6512 -26685 6562 -26645
rect 6622 -26645 6652 -26625
rect 6622 -26685 6672 -26645
rect 6512 -26755 6672 -26685
rect 6512 -26795 6562 -26755
rect 6532 -26815 6562 -26795
rect 6622 -26795 6672 -26755
rect 6622 -26815 6652 -26795
rect 6732 -26845 6792 -26585
rect 6722 -26855 6792 -26845
rect 6392 -26865 6472 -26855
rect 6392 -26925 6402 -26865
rect 6462 -26875 6472 -26865
rect 6712 -26865 6792 -26855
rect 6712 -26875 6722 -26865
rect 6462 -26925 6722 -26875
rect 6782 -26925 6792 -26865
rect 6392 -26935 6792 -26925
rect 6850 -26515 7250 -26505
rect 6850 -26575 6860 -26515
rect 6920 -26565 7180 -26515
rect 6920 -26575 6930 -26565
rect 6850 -26585 6930 -26575
rect 7170 -26575 7180 -26565
rect 7240 -26575 7250 -26515
rect 7170 -26585 7250 -26575
rect 6850 -26855 6910 -26585
rect 6990 -26645 7020 -26625
rect 6970 -26685 7020 -26645
rect 7080 -26645 7110 -26625
rect 7080 -26685 7130 -26645
rect 6970 -26755 7130 -26685
rect 6970 -26795 7020 -26755
rect 6990 -26815 7020 -26795
rect 7080 -26795 7130 -26755
rect 7080 -26815 7110 -26795
rect 7190 -26845 7250 -26585
rect 7180 -26855 7250 -26845
rect 6850 -26865 6930 -26855
rect 6850 -26925 6860 -26865
rect 6920 -26875 6930 -26865
rect 7170 -26865 7250 -26855
rect 7170 -26875 7180 -26865
rect 6920 -26925 7180 -26875
rect 7240 -26925 7250 -26865
rect 6850 -26935 7250 -26925
rect 7306 -26515 7706 -26505
rect 7306 -26575 7316 -26515
rect 7376 -26565 7636 -26515
rect 7376 -26575 7386 -26565
rect 7306 -26585 7386 -26575
rect 7626 -26575 7636 -26565
rect 7696 -26575 7706 -26515
rect 7626 -26585 7706 -26575
rect 7306 -26855 7366 -26585
rect 7446 -26645 7476 -26625
rect 7426 -26685 7476 -26645
rect 7536 -26645 7566 -26625
rect 7536 -26685 7586 -26645
rect 7426 -26755 7586 -26685
rect 7426 -26795 7476 -26755
rect 7446 -26815 7476 -26795
rect 7536 -26795 7586 -26755
rect 7536 -26815 7566 -26795
rect 7646 -26845 7706 -26585
rect 7636 -26855 7706 -26845
rect 7306 -26865 7386 -26855
rect 7306 -26925 7316 -26865
rect 7376 -26875 7386 -26865
rect 7626 -26865 7706 -26855
rect 7626 -26875 7636 -26865
rect 7376 -26925 7636 -26875
rect 7696 -26925 7706 -26865
rect 7306 -26935 7706 -26925
rect 7762 -26515 8162 -26505
rect 7762 -26575 7772 -26515
rect 7832 -26565 8092 -26515
rect 7832 -26575 7842 -26565
rect 7762 -26585 7842 -26575
rect 8082 -26575 8092 -26565
rect 8152 -26575 8162 -26515
rect 8082 -26585 8162 -26575
rect 7762 -26855 7822 -26585
rect 7902 -26645 7932 -26625
rect 7882 -26685 7932 -26645
rect 7992 -26645 8022 -26625
rect 7992 -26685 8042 -26645
rect 7882 -26755 8042 -26685
rect 7882 -26795 7932 -26755
rect 7902 -26815 7932 -26795
rect 7992 -26795 8042 -26755
rect 7992 -26815 8022 -26795
rect 8102 -26845 8162 -26585
rect 8092 -26855 8162 -26845
rect 7762 -26865 7842 -26855
rect 7762 -26925 7772 -26865
rect 7832 -26875 7842 -26865
rect 8082 -26865 8162 -26855
rect 8082 -26875 8092 -26865
rect 7832 -26925 8092 -26875
rect 8152 -26925 8162 -26865
rect 7762 -26935 8162 -26925
rect 8236 -26515 8636 -26505
rect 8236 -26575 8246 -26515
rect 8306 -26565 8566 -26515
rect 8306 -26575 8316 -26565
rect 8236 -26585 8316 -26575
rect 8556 -26575 8566 -26565
rect 8626 -26575 8636 -26515
rect 8556 -26585 8636 -26575
rect 8236 -26855 8296 -26585
rect 8376 -26645 8406 -26625
rect 8356 -26685 8406 -26645
rect 8466 -26645 8496 -26625
rect 8466 -26685 8516 -26645
rect 8356 -26755 8516 -26685
rect 8356 -26795 8406 -26755
rect 8376 -26815 8406 -26795
rect 8466 -26795 8516 -26755
rect 8466 -26815 8496 -26795
rect 8576 -26845 8636 -26585
rect 8566 -26855 8636 -26845
rect 8236 -26865 8316 -26855
rect 8236 -26925 8246 -26865
rect 8306 -26875 8316 -26865
rect 8556 -26865 8636 -26855
rect 8556 -26875 8566 -26865
rect 8306 -26925 8566 -26875
rect 8626 -26925 8636 -26865
rect 8236 -26935 8636 -26925
rect 8692 -26515 9092 -26505
rect 8692 -26575 8702 -26515
rect 8762 -26565 9022 -26515
rect 8762 -26575 8772 -26565
rect 8692 -26585 8772 -26575
rect 9012 -26575 9022 -26565
rect 9082 -26575 9092 -26515
rect 9012 -26585 9092 -26575
rect 8692 -26855 8752 -26585
rect 8832 -26645 8862 -26625
rect 8812 -26685 8862 -26645
rect 8922 -26645 8952 -26625
rect 8922 -26685 8972 -26645
rect 8812 -26755 8972 -26685
rect 8812 -26795 8862 -26755
rect 8832 -26815 8862 -26795
rect 8922 -26795 8972 -26755
rect 8922 -26815 8952 -26795
rect 9032 -26845 9092 -26585
rect 9022 -26855 9092 -26845
rect 8692 -26865 8772 -26855
rect 8692 -26925 8702 -26865
rect 8762 -26875 8772 -26865
rect 9012 -26865 9092 -26855
rect 9012 -26875 9022 -26865
rect 8762 -26925 9022 -26875
rect 9082 -26925 9092 -26865
rect 8692 -26935 9092 -26925
rect 9150 -26515 9550 -26505
rect 9150 -26575 9160 -26515
rect 9220 -26565 9480 -26515
rect 9220 -26575 9230 -26565
rect 9150 -26585 9230 -26575
rect 9470 -26575 9480 -26565
rect 9540 -26575 9550 -26515
rect 9470 -26585 9550 -26575
rect 9150 -26855 9210 -26585
rect 9290 -26645 9320 -26625
rect 9270 -26685 9320 -26645
rect 9380 -26645 9410 -26625
rect 9380 -26685 9430 -26645
rect 9270 -26755 9430 -26685
rect 9270 -26795 9320 -26755
rect 9290 -26815 9320 -26795
rect 9380 -26795 9430 -26755
rect 9380 -26815 9410 -26795
rect 9490 -26845 9550 -26585
rect 9480 -26855 9550 -26845
rect 9150 -26865 9230 -26855
rect 9150 -26925 9160 -26865
rect 9220 -26875 9230 -26865
rect 9470 -26865 9550 -26855
rect 9470 -26875 9480 -26865
rect 9220 -26925 9480 -26875
rect 9540 -26925 9550 -26865
rect 9150 -26935 9550 -26925
rect 9606 -26515 10006 -26505
rect 9606 -26575 9616 -26515
rect 9676 -26565 9936 -26515
rect 9676 -26575 9686 -26565
rect 9606 -26585 9686 -26575
rect 9926 -26575 9936 -26565
rect 9996 -26575 10006 -26515
rect 9926 -26585 10006 -26575
rect 9606 -26855 9666 -26585
rect 9746 -26645 9776 -26625
rect 9726 -26685 9776 -26645
rect 9836 -26645 9866 -26625
rect 9836 -26685 9886 -26645
rect 9726 -26755 9886 -26685
rect 9726 -26795 9776 -26755
rect 9746 -26815 9776 -26795
rect 9836 -26795 9886 -26755
rect 9836 -26815 9866 -26795
rect 9946 -26845 10006 -26585
rect 9936 -26855 10006 -26845
rect 9606 -26865 9686 -26855
rect 9606 -26925 9616 -26865
rect 9676 -26875 9686 -26865
rect 9926 -26865 10006 -26855
rect 9926 -26875 9936 -26865
rect 9676 -26925 9936 -26875
rect 9996 -26925 10006 -26865
rect 9606 -26935 10006 -26925
rect 10062 -26515 10462 -26505
rect 10062 -26575 10072 -26515
rect 10132 -26565 10392 -26515
rect 10132 -26575 10142 -26565
rect 10062 -26585 10142 -26575
rect 10382 -26575 10392 -26565
rect 10452 -26575 10462 -26515
rect 10382 -26585 10462 -26575
rect 10062 -26855 10122 -26585
rect 10202 -26645 10232 -26625
rect 10182 -26685 10232 -26645
rect 10292 -26645 10322 -26625
rect 10292 -26685 10342 -26645
rect 10182 -26755 10342 -26685
rect 10182 -26795 10232 -26755
rect 10202 -26815 10232 -26795
rect 10292 -26795 10342 -26755
rect 10292 -26815 10322 -26795
rect 10402 -26845 10462 -26585
rect 10392 -26855 10462 -26845
rect 10062 -26865 10142 -26855
rect 10062 -26925 10072 -26865
rect 10132 -26875 10142 -26865
rect 10382 -26865 10462 -26855
rect 10382 -26875 10392 -26865
rect 10132 -26925 10392 -26875
rect 10452 -26925 10462 -26865
rect 10062 -26935 10462 -26925
rect 10520 -26515 10920 -26505
rect 10520 -26575 10530 -26515
rect 10590 -26565 10850 -26515
rect 10590 -26575 10600 -26565
rect 10520 -26585 10600 -26575
rect 10840 -26575 10850 -26565
rect 10910 -26575 10920 -26515
rect 10840 -26585 10920 -26575
rect 10520 -26855 10580 -26585
rect 10660 -26645 10690 -26625
rect 10640 -26685 10690 -26645
rect 10750 -26645 10780 -26625
rect 10750 -26685 10800 -26645
rect 10640 -26755 10800 -26685
rect 10640 -26795 10690 -26755
rect 10660 -26815 10690 -26795
rect 10750 -26795 10800 -26755
rect 10750 -26815 10780 -26795
rect 10860 -26845 10920 -26585
rect 10850 -26855 10920 -26845
rect 10520 -26865 10600 -26855
rect 10520 -26925 10530 -26865
rect 10590 -26875 10600 -26865
rect 10840 -26865 10920 -26855
rect 10840 -26875 10850 -26865
rect 10590 -26925 10850 -26875
rect 10910 -26925 10920 -26865
rect 10520 -26935 10920 -26925
rect 10976 -26515 11376 -26505
rect 10976 -26575 10986 -26515
rect 11046 -26565 11306 -26515
rect 11046 -26575 11056 -26565
rect 10976 -26585 11056 -26575
rect 11296 -26575 11306 -26565
rect 11366 -26575 11376 -26515
rect 11296 -26585 11376 -26575
rect 10976 -26855 11036 -26585
rect 11116 -26645 11146 -26625
rect 11096 -26685 11146 -26645
rect 11206 -26645 11236 -26625
rect 11206 -26685 11256 -26645
rect 11096 -26755 11256 -26685
rect 11096 -26795 11146 -26755
rect 11116 -26815 11146 -26795
rect 11206 -26795 11256 -26755
rect 11206 -26815 11236 -26795
rect 11316 -26845 11376 -26585
rect 11306 -26855 11376 -26845
rect 10976 -26865 11056 -26855
rect 10976 -26925 10986 -26865
rect 11046 -26875 11056 -26865
rect 11296 -26865 11376 -26855
rect 11296 -26875 11306 -26865
rect 11046 -26925 11306 -26875
rect 11366 -26925 11376 -26865
rect 10976 -26935 11376 -26925
rect 11432 -26515 11832 -26505
rect 11432 -26575 11442 -26515
rect 11502 -26565 11762 -26515
rect 11502 -26575 11512 -26565
rect 11432 -26585 11512 -26575
rect 11752 -26575 11762 -26565
rect 11822 -26575 11832 -26515
rect 11752 -26585 11832 -26575
rect 11432 -26855 11492 -26585
rect 11572 -26645 11602 -26625
rect 11552 -26685 11602 -26645
rect 11662 -26645 11692 -26625
rect 11662 -26685 11712 -26645
rect 11552 -26755 11712 -26685
rect 11552 -26795 11602 -26755
rect 11572 -26815 11602 -26795
rect 11662 -26795 11712 -26755
rect 11662 -26815 11692 -26795
rect 11772 -26845 11832 -26585
rect 11762 -26855 11832 -26845
rect 11432 -26865 11512 -26855
rect 11432 -26925 11442 -26865
rect 11502 -26875 11512 -26865
rect 11752 -26865 11832 -26855
rect 11752 -26875 11762 -26865
rect 11502 -26925 11762 -26875
rect 11822 -26925 11832 -26865
rect 11432 -26935 11832 -26925
rect 11890 -26515 12290 -26505
rect 11890 -26575 11900 -26515
rect 11960 -26565 12220 -26515
rect 11960 -26575 11970 -26565
rect 11890 -26585 11970 -26575
rect 12210 -26575 12220 -26565
rect 12280 -26575 12290 -26515
rect 12210 -26585 12290 -26575
rect 11890 -26855 11950 -26585
rect 12030 -26645 12060 -26625
rect 12010 -26685 12060 -26645
rect 12120 -26645 12150 -26625
rect 12120 -26685 12170 -26645
rect 12010 -26755 12170 -26685
rect 12010 -26795 12060 -26755
rect 12030 -26815 12060 -26795
rect 12120 -26795 12170 -26755
rect 12120 -26815 12150 -26795
rect 12230 -26845 12290 -26585
rect 12220 -26855 12290 -26845
rect 11890 -26865 11970 -26855
rect 11890 -26925 11900 -26865
rect 11960 -26875 11970 -26865
rect 12210 -26865 12290 -26855
rect 12210 -26875 12220 -26865
rect 11960 -26925 12220 -26875
rect 12280 -26925 12290 -26865
rect 11890 -26935 12290 -26925
rect 12346 -26515 12746 -26505
rect 12346 -26575 12356 -26515
rect 12416 -26565 12676 -26515
rect 12416 -26575 12426 -26565
rect 12346 -26585 12426 -26575
rect 12666 -26575 12676 -26565
rect 12736 -26575 12746 -26515
rect 12666 -26585 12746 -26575
rect 12346 -26855 12406 -26585
rect 12486 -26645 12516 -26625
rect 12466 -26685 12516 -26645
rect 12576 -26645 12606 -26625
rect 12576 -26685 12626 -26645
rect 12466 -26755 12626 -26685
rect 12466 -26795 12516 -26755
rect 12486 -26815 12516 -26795
rect 12576 -26795 12626 -26755
rect 12576 -26815 12606 -26795
rect 12686 -26845 12746 -26585
rect 12676 -26855 12746 -26845
rect 12346 -26865 12426 -26855
rect 12346 -26925 12356 -26865
rect 12416 -26875 12426 -26865
rect 12666 -26865 12746 -26855
rect 12666 -26875 12676 -26865
rect 12416 -26925 12676 -26875
rect 12736 -26925 12746 -26865
rect 12346 -26935 12746 -26925
rect 12802 -26515 13202 -26505
rect 12802 -26575 12812 -26515
rect 12872 -26565 13132 -26515
rect 12872 -26575 12882 -26565
rect 12802 -26585 12882 -26575
rect 13122 -26575 13132 -26565
rect 13192 -26575 13202 -26515
rect 13122 -26585 13202 -26575
rect 12802 -26855 12862 -26585
rect 12942 -26645 12972 -26625
rect 12922 -26685 12972 -26645
rect 13032 -26645 13062 -26625
rect 13032 -26685 13082 -26645
rect 12922 -26755 13082 -26685
rect 12922 -26795 12972 -26755
rect 12942 -26815 12972 -26795
rect 13032 -26795 13082 -26755
rect 13032 -26815 13062 -26795
rect 13142 -26845 13202 -26585
rect 13132 -26855 13202 -26845
rect 12802 -26865 12882 -26855
rect 12802 -26925 12812 -26865
rect 12872 -26875 12882 -26865
rect 13122 -26865 13202 -26855
rect 13122 -26875 13132 -26865
rect 12872 -26925 13132 -26875
rect 13192 -26925 13202 -26865
rect 12802 -26935 13202 -26925
rect 13260 -26515 13660 -26505
rect 13260 -26575 13270 -26515
rect 13330 -26565 13590 -26515
rect 13330 -26575 13340 -26565
rect 13260 -26585 13340 -26575
rect 13580 -26575 13590 -26565
rect 13650 -26575 13660 -26515
rect 13580 -26585 13660 -26575
rect 13260 -26855 13320 -26585
rect 13400 -26645 13430 -26625
rect 13380 -26685 13430 -26645
rect 13490 -26645 13520 -26625
rect 13490 -26685 13540 -26645
rect 13380 -26755 13540 -26685
rect 13380 -26795 13430 -26755
rect 13400 -26815 13430 -26795
rect 13490 -26795 13540 -26755
rect 13490 -26815 13520 -26795
rect 13600 -26845 13660 -26585
rect 13590 -26855 13660 -26845
rect 13260 -26865 13340 -26855
rect 13260 -26925 13270 -26865
rect 13330 -26875 13340 -26865
rect 13580 -26865 13660 -26855
rect 13580 -26875 13590 -26865
rect 13330 -26925 13590 -26875
rect 13650 -26925 13660 -26865
rect 13260 -26935 13660 -26925
rect 13716 -26515 14116 -26505
rect 13716 -26575 13726 -26515
rect 13786 -26565 14046 -26515
rect 13786 -26575 13796 -26565
rect 13716 -26585 13796 -26575
rect 14036 -26575 14046 -26565
rect 14106 -26575 14116 -26515
rect 14036 -26585 14116 -26575
rect 13716 -26855 13776 -26585
rect 13856 -26645 13886 -26625
rect 13836 -26685 13886 -26645
rect 13946 -26645 13976 -26625
rect 13946 -26685 13996 -26645
rect 13836 -26755 13996 -26685
rect 13836 -26795 13886 -26755
rect 13856 -26815 13886 -26795
rect 13946 -26795 13996 -26755
rect 13946 -26815 13976 -26795
rect 14056 -26845 14116 -26585
rect 14046 -26855 14116 -26845
rect 13716 -26865 13796 -26855
rect 13716 -26925 13726 -26865
rect 13786 -26875 13796 -26865
rect 14036 -26865 14116 -26855
rect 14036 -26875 14046 -26865
rect 13786 -26925 14046 -26875
rect 14106 -26925 14116 -26865
rect 13716 -26935 14116 -26925
rect 14172 -26515 14572 -26505
rect 14172 -26575 14182 -26515
rect 14242 -26565 14502 -26515
rect 14242 -26575 14252 -26565
rect 14172 -26585 14252 -26575
rect 14492 -26575 14502 -26565
rect 14562 -26575 14572 -26515
rect 14492 -26585 14572 -26575
rect 14172 -26855 14232 -26585
rect 14312 -26645 14342 -26625
rect 14292 -26685 14342 -26645
rect 14402 -26645 14432 -26625
rect 14402 -26685 14452 -26645
rect 14292 -26755 14452 -26685
rect 14292 -26795 14342 -26755
rect 14312 -26815 14342 -26795
rect 14402 -26795 14452 -26755
rect 14402 -26815 14432 -26795
rect 14512 -26845 14572 -26585
rect 14502 -26855 14572 -26845
rect 14172 -26865 14252 -26855
rect 14172 -26925 14182 -26865
rect 14242 -26875 14252 -26865
rect 14492 -26865 14572 -26855
rect 14492 -26875 14502 -26865
rect 14242 -26925 14502 -26875
rect 14562 -26925 14572 -26865
rect 14172 -26935 14572 -26925
rect 14630 -26515 15030 -26505
rect 14630 -26575 14640 -26515
rect 14700 -26565 14960 -26515
rect 14700 -26575 14710 -26565
rect 14630 -26585 14710 -26575
rect 14950 -26575 14960 -26565
rect 15020 -26575 15030 -26515
rect 14950 -26585 15030 -26575
rect 14630 -26855 14690 -26585
rect 14770 -26645 14800 -26625
rect 14750 -26685 14800 -26645
rect 14860 -26645 14890 -26625
rect 14860 -26685 14910 -26645
rect 14750 -26755 14910 -26685
rect 14750 -26795 14800 -26755
rect 14770 -26815 14800 -26795
rect 14860 -26795 14910 -26755
rect 14860 -26815 14890 -26795
rect 14970 -26845 15030 -26585
rect 14960 -26855 15030 -26845
rect 14630 -26865 14710 -26855
rect 14630 -26925 14640 -26865
rect 14700 -26875 14710 -26865
rect 14950 -26865 15030 -26855
rect 14950 -26875 14960 -26865
rect 14700 -26925 14960 -26875
rect 15020 -26925 15030 -26865
rect 14630 -26935 15030 -26925
rect 15086 -26515 15486 -26505
rect 15086 -26575 15096 -26515
rect 15156 -26565 15416 -26515
rect 15156 -26575 15166 -26565
rect 15086 -26585 15166 -26575
rect 15406 -26575 15416 -26565
rect 15476 -26575 15486 -26515
rect 15406 -26585 15486 -26575
rect 15086 -26855 15146 -26585
rect 15226 -26645 15256 -26625
rect 15206 -26685 15256 -26645
rect 15316 -26645 15346 -26625
rect 15316 -26685 15366 -26645
rect 15206 -26755 15366 -26685
rect 15206 -26795 15256 -26755
rect 15226 -26815 15256 -26795
rect 15316 -26795 15366 -26755
rect 15316 -26815 15346 -26795
rect 15426 -26845 15486 -26585
rect 15416 -26855 15486 -26845
rect 15086 -26865 15166 -26855
rect 15086 -26925 15096 -26865
rect 15156 -26875 15166 -26865
rect 15406 -26865 15486 -26855
rect 15406 -26875 15416 -26865
rect 15156 -26925 15416 -26875
rect 15476 -26925 15486 -26865
rect 15086 -26935 15486 -26925
rect 0 -27017 400 -27007
rect 0 -27077 10 -27017
rect 70 -27067 330 -27017
rect 70 -27077 80 -27067
rect 0 -27087 80 -27077
rect 320 -27077 330 -27067
rect 390 -27077 400 -27017
rect 320 -27087 400 -27077
rect 0 -27357 60 -27087
rect 140 -27147 170 -27127
rect 120 -27187 170 -27147
rect 230 -27147 260 -27127
rect 230 -27187 280 -27147
rect 120 -27257 280 -27187
rect 120 -27297 170 -27257
rect 140 -27317 170 -27297
rect 230 -27297 280 -27257
rect 230 -27317 260 -27297
rect 340 -27347 400 -27087
rect 330 -27357 400 -27347
rect 0 -27367 80 -27357
rect 0 -27427 10 -27367
rect 70 -27377 80 -27367
rect 320 -27367 400 -27357
rect 320 -27377 330 -27367
rect 70 -27427 330 -27377
rect 390 -27427 400 -27367
rect 0 -27437 400 -27427
rect 456 -27017 856 -27007
rect 456 -27077 466 -27017
rect 526 -27067 786 -27017
rect 526 -27077 536 -27067
rect 456 -27087 536 -27077
rect 776 -27077 786 -27067
rect 846 -27077 856 -27017
rect 776 -27087 856 -27077
rect 456 -27357 516 -27087
rect 596 -27147 626 -27127
rect 576 -27187 626 -27147
rect 686 -27147 716 -27127
rect 686 -27187 736 -27147
rect 576 -27257 736 -27187
rect 576 -27297 626 -27257
rect 596 -27317 626 -27297
rect 686 -27297 736 -27257
rect 686 -27317 716 -27297
rect 796 -27347 856 -27087
rect 786 -27357 856 -27347
rect 456 -27367 536 -27357
rect 456 -27427 466 -27367
rect 526 -27377 536 -27367
rect 776 -27367 856 -27357
rect 776 -27377 786 -27367
rect 526 -27427 786 -27377
rect 846 -27427 856 -27367
rect 456 -27437 856 -27427
rect 912 -27017 1312 -27007
rect 912 -27077 922 -27017
rect 982 -27067 1242 -27017
rect 982 -27077 992 -27067
rect 912 -27087 992 -27077
rect 1232 -27077 1242 -27067
rect 1302 -27077 1312 -27017
rect 1232 -27087 1312 -27077
rect 912 -27357 972 -27087
rect 1052 -27147 1082 -27127
rect 1032 -27187 1082 -27147
rect 1142 -27147 1172 -27127
rect 1142 -27187 1192 -27147
rect 1032 -27257 1192 -27187
rect 1032 -27297 1082 -27257
rect 1052 -27317 1082 -27297
rect 1142 -27297 1192 -27257
rect 1142 -27317 1172 -27297
rect 1252 -27347 1312 -27087
rect 1242 -27357 1312 -27347
rect 912 -27367 992 -27357
rect 912 -27427 922 -27367
rect 982 -27377 992 -27367
rect 1232 -27367 1312 -27357
rect 1232 -27377 1242 -27367
rect 982 -27427 1242 -27377
rect 1302 -27427 1312 -27367
rect 912 -27437 1312 -27427
rect 1370 -27017 1770 -27007
rect 1370 -27077 1380 -27017
rect 1440 -27067 1700 -27017
rect 1440 -27077 1450 -27067
rect 1370 -27087 1450 -27077
rect 1690 -27077 1700 -27067
rect 1760 -27077 1770 -27017
rect 1690 -27087 1770 -27077
rect 1370 -27357 1430 -27087
rect 1510 -27147 1540 -27127
rect 1490 -27187 1540 -27147
rect 1600 -27147 1630 -27127
rect 1600 -27187 1650 -27147
rect 1490 -27257 1650 -27187
rect 1490 -27297 1540 -27257
rect 1510 -27317 1540 -27297
rect 1600 -27297 1650 -27257
rect 1600 -27317 1630 -27297
rect 1710 -27347 1770 -27087
rect 1700 -27357 1770 -27347
rect 1370 -27367 1450 -27357
rect 1370 -27427 1380 -27367
rect 1440 -27377 1450 -27367
rect 1690 -27367 1770 -27357
rect 1690 -27377 1700 -27367
rect 1440 -27427 1700 -27377
rect 1760 -27427 1770 -27367
rect 1370 -27437 1770 -27427
rect 1826 -27017 2226 -27007
rect 1826 -27077 1836 -27017
rect 1896 -27067 2156 -27017
rect 1896 -27077 1906 -27067
rect 1826 -27087 1906 -27077
rect 2146 -27077 2156 -27067
rect 2216 -27077 2226 -27017
rect 2146 -27087 2226 -27077
rect 1826 -27357 1886 -27087
rect 1966 -27147 1996 -27127
rect 1946 -27187 1996 -27147
rect 2056 -27147 2086 -27127
rect 2056 -27187 2106 -27147
rect 1946 -27257 2106 -27187
rect 1946 -27297 1996 -27257
rect 1966 -27317 1996 -27297
rect 2056 -27297 2106 -27257
rect 2056 -27317 2086 -27297
rect 2166 -27347 2226 -27087
rect 2156 -27357 2226 -27347
rect 1826 -27367 1906 -27357
rect 1826 -27427 1836 -27367
rect 1896 -27377 1906 -27367
rect 2146 -27367 2226 -27357
rect 2146 -27377 2156 -27367
rect 1896 -27427 2156 -27377
rect 2216 -27427 2226 -27367
rect 1826 -27437 2226 -27427
rect 2282 -27017 2682 -27007
rect 2282 -27077 2292 -27017
rect 2352 -27067 2612 -27017
rect 2352 -27077 2362 -27067
rect 2282 -27087 2362 -27077
rect 2602 -27077 2612 -27067
rect 2672 -27077 2682 -27017
rect 2602 -27087 2682 -27077
rect 2282 -27357 2342 -27087
rect 2422 -27147 2452 -27127
rect 2402 -27187 2452 -27147
rect 2512 -27147 2542 -27127
rect 2512 -27187 2562 -27147
rect 2402 -27257 2562 -27187
rect 2402 -27297 2452 -27257
rect 2422 -27317 2452 -27297
rect 2512 -27297 2562 -27257
rect 2512 -27317 2542 -27297
rect 2622 -27347 2682 -27087
rect 2612 -27357 2682 -27347
rect 2282 -27367 2362 -27357
rect 2282 -27427 2292 -27367
rect 2352 -27377 2362 -27367
rect 2602 -27367 2682 -27357
rect 2602 -27377 2612 -27367
rect 2352 -27427 2612 -27377
rect 2672 -27427 2682 -27367
rect 2282 -27437 2682 -27427
rect 2740 -27017 3140 -27007
rect 2740 -27077 2750 -27017
rect 2810 -27067 3070 -27017
rect 2810 -27077 2820 -27067
rect 2740 -27087 2820 -27077
rect 3060 -27077 3070 -27067
rect 3130 -27077 3140 -27017
rect 3060 -27087 3140 -27077
rect 2740 -27357 2800 -27087
rect 2880 -27147 2910 -27127
rect 2860 -27187 2910 -27147
rect 2970 -27147 3000 -27127
rect 2970 -27187 3020 -27147
rect 2860 -27257 3020 -27187
rect 2860 -27297 2910 -27257
rect 2880 -27317 2910 -27297
rect 2970 -27297 3020 -27257
rect 2970 -27317 3000 -27297
rect 3080 -27347 3140 -27087
rect 3070 -27357 3140 -27347
rect 2740 -27367 2820 -27357
rect 2740 -27427 2750 -27367
rect 2810 -27377 2820 -27367
rect 3060 -27367 3140 -27357
rect 3060 -27377 3070 -27367
rect 2810 -27427 3070 -27377
rect 3130 -27427 3140 -27367
rect 2740 -27437 3140 -27427
rect 3196 -27017 3596 -27007
rect 3196 -27077 3206 -27017
rect 3266 -27067 3526 -27017
rect 3266 -27077 3276 -27067
rect 3196 -27087 3276 -27077
rect 3516 -27077 3526 -27067
rect 3586 -27077 3596 -27017
rect 3516 -27087 3596 -27077
rect 3196 -27357 3256 -27087
rect 3336 -27147 3366 -27127
rect 3316 -27187 3366 -27147
rect 3426 -27147 3456 -27127
rect 3426 -27187 3476 -27147
rect 3316 -27257 3476 -27187
rect 3316 -27297 3366 -27257
rect 3336 -27317 3366 -27297
rect 3426 -27297 3476 -27257
rect 3426 -27317 3456 -27297
rect 3536 -27347 3596 -27087
rect 3526 -27357 3596 -27347
rect 3196 -27367 3276 -27357
rect 3196 -27427 3206 -27367
rect 3266 -27377 3276 -27367
rect 3516 -27367 3596 -27357
rect 3516 -27377 3526 -27367
rect 3266 -27427 3526 -27377
rect 3586 -27427 3596 -27367
rect 3196 -27437 3596 -27427
rect 3652 -27017 4052 -27007
rect 3652 -27077 3662 -27017
rect 3722 -27067 3982 -27017
rect 3722 -27077 3732 -27067
rect 3652 -27087 3732 -27077
rect 3972 -27077 3982 -27067
rect 4042 -27077 4052 -27017
rect 3972 -27087 4052 -27077
rect 3652 -27357 3712 -27087
rect 3792 -27147 3822 -27127
rect 3772 -27187 3822 -27147
rect 3882 -27147 3912 -27127
rect 3882 -27187 3932 -27147
rect 3772 -27257 3932 -27187
rect 3772 -27297 3822 -27257
rect 3792 -27317 3822 -27297
rect 3882 -27297 3932 -27257
rect 3882 -27317 3912 -27297
rect 3992 -27347 4052 -27087
rect 3982 -27357 4052 -27347
rect 3652 -27367 3732 -27357
rect 3652 -27427 3662 -27367
rect 3722 -27377 3732 -27367
rect 3972 -27367 4052 -27357
rect 3972 -27377 3982 -27367
rect 3722 -27427 3982 -27377
rect 4042 -27427 4052 -27367
rect 3652 -27437 4052 -27427
rect 4110 -27017 4510 -27007
rect 4110 -27077 4120 -27017
rect 4180 -27067 4440 -27017
rect 4180 -27077 4190 -27067
rect 4110 -27087 4190 -27077
rect 4430 -27077 4440 -27067
rect 4500 -27077 4510 -27017
rect 4430 -27087 4510 -27077
rect 4110 -27357 4170 -27087
rect 4250 -27147 4280 -27127
rect 4230 -27187 4280 -27147
rect 4340 -27147 4370 -27127
rect 4340 -27187 4390 -27147
rect 4230 -27257 4390 -27187
rect 4230 -27297 4280 -27257
rect 4250 -27317 4280 -27297
rect 4340 -27297 4390 -27257
rect 4340 -27317 4370 -27297
rect 4450 -27347 4510 -27087
rect 4440 -27357 4510 -27347
rect 4110 -27367 4190 -27357
rect 4110 -27427 4120 -27367
rect 4180 -27377 4190 -27367
rect 4430 -27367 4510 -27357
rect 4430 -27377 4440 -27367
rect 4180 -27427 4440 -27377
rect 4500 -27427 4510 -27367
rect 4110 -27437 4510 -27427
rect 4566 -27017 4966 -27007
rect 4566 -27077 4576 -27017
rect 4636 -27067 4896 -27017
rect 4636 -27077 4646 -27067
rect 4566 -27087 4646 -27077
rect 4886 -27077 4896 -27067
rect 4956 -27077 4966 -27017
rect 4886 -27087 4966 -27077
rect 4566 -27357 4626 -27087
rect 4706 -27147 4736 -27127
rect 4686 -27187 4736 -27147
rect 4796 -27147 4826 -27127
rect 4796 -27187 4846 -27147
rect 4686 -27257 4846 -27187
rect 4686 -27297 4736 -27257
rect 4706 -27317 4736 -27297
rect 4796 -27297 4846 -27257
rect 4796 -27317 4826 -27297
rect 4906 -27347 4966 -27087
rect 4896 -27357 4966 -27347
rect 4566 -27367 4646 -27357
rect 4566 -27427 4576 -27367
rect 4636 -27377 4646 -27367
rect 4886 -27367 4966 -27357
rect 4886 -27377 4896 -27367
rect 4636 -27427 4896 -27377
rect 4956 -27427 4966 -27367
rect 4566 -27437 4966 -27427
rect 5022 -27017 5422 -27007
rect 5022 -27077 5032 -27017
rect 5092 -27067 5352 -27017
rect 5092 -27077 5102 -27067
rect 5022 -27087 5102 -27077
rect 5342 -27077 5352 -27067
rect 5412 -27077 5422 -27017
rect 5342 -27087 5422 -27077
rect 5022 -27357 5082 -27087
rect 5162 -27147 5192 -27127
rect 5142 -27187 5192 -27147
rect 5252 -27147 5282 -27127
rect 5252 -27187 5302 -27147
rect 5142 -27257 5302 -27187
rect 5142 -27297 5192 -27257
rect 5162 -27317 5192 -27297
rect 5252 -27297 5302 -27257
rect 5252 -27317 5282 -27297
rect 5362 -27347 5422 -27087
rect 5352 -27357 5422 -27347
rect 5022 -27367 5102 -27357
rect 5022 -27427 5032 -27367
rect 5092 -27377 5102 -27367
rect 5342 -27367 5422 -27357
rect 5342 -27377 5352 -27367
rect 5092 -27427 5352 -27377
rect 5412 -27427 5422 -27367
rect 5022 -27437 5422 -27427
rect 5480 -27017 5880 -27007
rect 5480 -27077 5490 -27017
rect 5550 -27067 5810 -27017
rect 5550 -27077 5560 -27067
rect 5480 -27087 5560 -27077
rect 5800 -27077 5810 -27067
rect 5870 -27077 5880 -27017
rect 5800 -27087 5880 -27077
rect 5480 -27357 5540 -27087
rect 5620 -27147 5650 -27127
rect 5600 -27187 5650 -27147
rect 5710 -27147 5740 -27127
rect 5710 -27187 5760 -27147
rect 5600 -27257 5760 -27187
rect 5600 -27297 5650 -27257
rect 5620 -27317 5650 -27297
rect 5710 -27297 5760 -27257
rect 5710 -27317 5740 -27297
rect 5820 -27347 5880 -27087
rect 5810 -27357 5880 -27347
rect 5480 -27367 5560 -27357
rect 5480 -27427 5490 -27367
rect 5550 -27377 5560 -27367
rect 5800 -27367 5880 -27357
rect 5800 -27377 5810 -27367
rect 5550 -27427 5810 -27377
rect 5870 -27427 5880 -27367
rect 5480 -27437 5880 -27427
rect 5936 -27017 6336 -27007
rect 5936 -27077 5946 -27017
rect 6006 -27067 6266 -27017
rect 6006 -27077 6016 -27067
rect 5936 -27087 6016 -27077
rect 6256 -27077 6266 -27067
rect 6326 -27077 6336 -27017
rect 6256 -27087 6336 -27077
rect 5936 -27357 5996 -27087
rect 6076 -27147 6106 -27127
rect 6056 -27187 6106 -27147
rect 6166 -27147 6196 -27127
rect 6166 -27187 6216 -27147
rect 6056 -27257 6216 -27187
rect 6056 -27297 6106 -27257
rect 6076 -27317 6106 -27297
rect 6166 -27297 6216 -27257
rect 6166 -27317 6196 -27297
rect 6276 -27347 6336 -27087
rect 6266 -27357 6336 -27347
rect 5936 -27367 6016 -27357
rect 5936 -27427 5946 -27367
rect 6006 -27377 6016 -27367
rect 6256 -27367 6336 -27357
rect 6256 -27377 6266 -27367
rect 6006 -27427 6266 -27377
rect 6326 -27427 6336 -27367
rect 5936 -27437 6336 -27427
rect 6392 -27017 6792 -27007
rect 6392 -27077 6402 -27017
rect 6462 -27067 6722 -27017
rect 6462 -27077 6472 -27067
rect 6392 -27087 6472 -27077
rect 6712 -27077 6722 -27067
rect 6782 -27077 6792 -27017
rect 6712 -27087 6792 -27077
rect 6392 -27357 6452 -27087
rect 6532 -27147 6562 -27127
rect 6512 -27187 6562 -27147
rect 6622 -27147 6652 -27127
rect 6622 -27187 6672 -27147
rect 6512 -27257 6672 -27187
rect 6512 -27297 6562 -27257
rect 6532 -27317 6562 -27297
rect 6622 -27297 6672 -27257
rect 6622 -27317 6652 -27297
rect 6732 -27347 6792 -27087
rect 6722 -27357 6792 -27347
rect 6392 -27367 6472 -27357
rect 6392 -27427 6402 -27367
rect 6462 -27377 6472 -27367
rect 6712 -27367 6792 -27357
rect 6712 -27377 6722 -27367
rect 6462 -27427 6722 -27377
rect 6782 -27427 6792 -27367
rect 6392 -27437 6792 -27427
rect 6850 -27017 7250 -27007
rect 6850 -27077 6860 -27017
rect 6920 -27067 7180 -27017
rect 6920 -27077 6930 -27067
rect 6850 -27087 6930 -27077
rect 7170 -27077 7180 -27067
rect 7240 -27077 7250 -27017
rect 7170 -27087 7250 -27077
rect 6850 -27357 6910 -27087
rect 6990 -27147 7020 -27127
rect 6970 -27187 7020 -27147
rect 7080 -27147 7110 -27127
rect 7080 -27187 7130 -27147
rect 6970 -27257 7130 -27187
rect 6970 -27297 7020 -27257
rect 6990 -27317 7020 -27297
rect 7080 -27297 7130 -27257
rect 7080 -27317 7110 -27297
rect 7190 -27347 7250 -27087
rect 7180 -27357 7250 -27347
rect 6850 -27367 6930 -27357
rect 6850 -27427 6860 -27367
rect 6920 -27377 6930 -27367
rect 7170 -27367 7250 -27357
rect 7170 -27377 7180 -27367
rect 6920 -27427 7180 -27377
rect 7240 -27427 7250 -27367
rect 6850 -27437 7250 -27427
rect 7306 -27017 7706 -27007
rect 7306 -27077 7316 -27017
rect 7376 -27067 7636 -27017
rect 7376 -27077 7386 -27067
rect 7306 -27087 7386 -27077
rect 7626 -27077 7636 -27067
rect 7696 -27077 7706 -27017
rect 7626 -27087 7706 -27077
rect 7306 -27357 7366 -27087
rect 7446 -27147 7476 -27127
rect 7426 -27187 7476 -27147
rect 7536 -27147 7566 -27127
rect 7536 -27187 7586 -27147
rect 7426 -27257 7586 -27187
rect 7426 -27297 7476 -27257
rect 7446 -27317 7476 -27297
rect 7536 -27297 7586 -27257
rect 7536 -27317 7566 -27297
rect 7646 -27347 7706 -27087
rect 7636 -27357 7706 -27347
rect 7306 -27367 7386 -27357
rect 7306 -27427 7316 -27367
rect 7376 -27377 7386 -27367
rect 7626 -27367 7706 -27357
rect 7626 -27377 7636 -27367
rect 7376 -27427 7636 -27377
rect 7696 -27427 7706 -27367
rect 7306 -27437 7706 -27427
rect 7762 -27017 8162 -27007
rect 7762 -27077 7772 -27017
rect 7832 -27067 8092 -27017
rect 7832 -27077 7842 -27067
rect 7762 -27087 7842 -27077
rect 8082 -27077 8092 -27067
rect 8152 -27077 8162 -27017
rect 8082 -27087 8162 -27077
rect 7762 -27357 7822 -27087
rect 7902 -27147 7932 -27127
rect 7882 -27187 7932 -27147
rect 7992 -27147 8022 -27127
rect 7992 -27187 8042 -27147
rect 7882 -27257 8042 -27187
rect 7882 -27297 7932 -27257
rect 7902 -27317 7932 -27297
rect 7992 -27297 8042 -27257
rect 7992 -27317 8022 -27297
rect 8102 -27347 8162 -27087
rect 8092 -27357 8162 -27347
rect 7762 -27367 7842 -27357
rect 7762 -27427 7772 -27367
rect 7832 -27377 7842 -27367
rect 8082 -27367 8162 -27357
rect 8082 -27377 8092 -27367
rect 7832 -27427 8092 -27377
rect 8152 -27427 8162 -27367
rect 7762 -27437 8162 -27427
rect 8236 -27017 8636 -27007
rect 8236 -27077 8246 -27017
rect 8306 -27067 8566 -27017
rect 8306 -27077 8316 -27067
rect 8236 -27087 8316 -27077
rect 8556 -27077 8566 -27067
rect 8626 -27077 8636 -27017
rect 8556 -27087 8636 -27077
rect 8236 -27357 8296 -27087
rect 8376 -27147 8406 -27127
rect 8356 -27187 8406 -27147
rect 8466 -27147 8496 -27127
rect 8466 -27187 8516 -27147
rect 8356 -27257 8516 -27187
rect 8356 -27297 8406 -27257
rect 8376 -27317 8406 -27297
rect 8466 -27297 8516 -27257
rect 8466 -27317 8496 -27297
rect 8576 -27347 8636 -27087
rect 8566 -27357 8636 -27347
rect 8236 -27367 8316 -27357
rect 8236 -27427 8246 -27367
rect 8306 -27377 8316 -27367
rect 8556 -27367 8636 -27357
rect 8556 -27377 8566 -27367
rect 8306 -27427 8566 -27377
rect 8626 -27427 8636 -27367
rect 8236 -27437 8636 -27427
rect 8692 -27017 9092 -27007
rect 8692 -27077 8702 -27017
rect 8762 -27067 9022 -27017
rect 8762 -27077 8772 -27067
rect 8692 -27087 8772 -27077
rect 9012 -27077 9022 -27067
rect 9082 -27077 9092 -27017
rect 9012 -27087 9092 -27077
rect 8692 -27357 8752 -27087
rect 8832 -27147 8862 -27127
rect 8812 -27187 8862 -27147
rect 8922 -27147 8952 -27127
rect 8922 -27187 8972 -27147
rect 8812 -27257 8972 -27187
rect 8812 -27297 8862 -27257
rect 8832 -27317 8862 -27297
rect 8922 -27297 8972 -27257
rect 8922 -27317 8952 -27297
rect 9032 -27347 9092 -27087
rect 9022 -27357 9092 -27347
rect 8692 -27367 8772 -27357
rect 8692 -27427 8702 -27367
rect 8762 -27377 8772 -27367
rect 9012 -27367 9092 -27357
rect 9012 -27377 9022 -27367
rect 8762 -27427 9022 -27377
rect 9082 -27427 9092 -27367
rect 8692 -27437 9092 -27427
rect 9150 -27017 9550 -27007
rect 9150 -27077 9160 -27017
rect 9220 -27067 9480 -27017
rect 9220 -27077 9230 -27067
rect 9150 -27087 9230 -27077
rect 9470 -27077 9480 -27067
rect 9540 -27077 9550 -27017
rect 9470 -27087 9550 -27077
rect 9150 -27357 9210 -27087
rect 9290 -27147 9320 -27127
rect 9270 -27187 9320 -27147
rect 9380 -27147 9410 -27127
rect 9380 -27187 9430 -27147
rect 9270 -27257 9430 -27187
rect 9270 -27297 9320 -27257
rect 9290 -27317 9320 -27297
rect 9380 -27297 9430 -27257
rect 9380 -27317 9410 -27297
rect 9490 -27347 9550 -27087
rect 9480 -27357 9550 -27347
rect 9150 -27367 9230 -27357
rect 9150 -27427 9160 -27367
rect 9220 -27377 9230 -27367
rect 9470 -27367 9550 -27357
rect 9470 -27377 9480 -27367
rect 9220 -27427 9480 -27377
rect 9540 -27427 9550 -27367
rect 9150 -27437 9550 -27427
rect 9606 -27017 10006 -27007
rect 9606 -27077 9616 -27017
rect 9676 -27067 9936 -27017
rect 9676 -27077 9686 -27067
rect 9606 -27087 9686 -27077
rect 9926 -27077 9936 -27067
rect 9996 -27077 10006 -27017
rect 9926 -27087 10006 -27077
rect 9606 -27357 9666 -27087
rect 9746 -27147 9776 -27127
rect 9726 -27187 9776 -27147
rect 9836 -27147 9866 -27127
rect 9836 -27187 9886 -27147
rect 9726 -27257 9886 -27187
rect 9726 -27297 9776 -27257
rect 9746 -27317 9776 -27297
rect 9836 -27297 9886 -27257
rect 9836 -27317 9866 -27297
rect 9946 -27347 10006 -27087
rect 9936 -27357 10006 -27347
rect 9606 -27367 9686 -27357
rect 9606 -27427 9616 -27367
rect 9676 -27377 9686 -27367
rect 9926 -27367 10006 -27357
rect 9926 -27377 9936 -27367
rect 9676 -27427 9936 -27377
rect 9996 -27427 10006 -27367
rect 9606 -27437 10006 -27427
rect 10062 -27017 10462 -27007
rect 10062 -27077 10072 -27017
rect 10132 -27067 10392 -27017
rect 10132 -27077 10142 -27067
rect 10062 -27087 10142 -27077
rect 10382 -27077 10392 -27067
rect 10452 -27077 10462 -27017
rect 10382 -27087 10462 -27077
rect 10062 -27357 10122 -27087
rect 10202 -27147 10232 -27127
rect 10182 -27187 10232 -27147
rect 10292 -27147 10322 -27127
rect 10292 -27187 10342 -27147
rect 10182 -27257 10342 -27187
rect 10182 -27297 10232 -27257
rect 10202 -27317 10232 -27297
rect 10292 -27297 10342 -27257
rect 10292 -27317 10322 -27297
rect 10402 -27347 10462 -27087
rect 10392 -27357 10462 -27347
rect 10062 -27367 10142 -27357
rect 10062 -27427 10072 -27367
rect 10132 -27377 10142 -27367
rect 10382 -27367 10462 -27357
rect 10382 -27377 10392 -27367
rect 10132 -27427 10392 -27377
rect 10452 -27427 10462 -27367
rect 10062 -27437 10462 -27427
rect 10520 -27017 10920 -27007
rect 10520 -27077 10530 -27017
rect 10590 -27067 10850 -27017
rect 10590 -27077 10600 -27067
rect 10520 -27087 10600 -27077
rect 10840 -27077 10850 -27067
rect 10910 -27077 10920 -27017
rect 10840 -27087 10920 -27077
rect 10520 -27357 10580 -27087
rect 10660 -27147 10690 -27127
rect 10640 -27187 10690 -27147
rect 10750 -27147 10780 -27127
rect 10750 -27187 10800 -27147
rect 10640 -27257 10800 -27187
rect 10640 -27297 10690 -27257
rect 10660 -27317 10690 -27297
rect 10750 -27297 10800 -27257
rect 10750 -27317 10780 -27297
rect 10860 -27347 10920 -27087
rect 10850 -27357 10920 -27347
rect 10520 -27367 10600 -27357
rect 10520 -27427 10530 -27367
rect 10590 -27377 10600 -27367
rect 10840 -27367 10920 -27357
rect 10840 -27377 10850 -27367
rect 10590 -27427 10850 -27377
rect 10910 -27427 10920 -27367
rect 10520 -27437 10920 -27427
rect 10976 -27017 11376 -27007
rect 10976 -27077 10986 -27017
rect 11046 -27067 11306 -27017
rect 11046 -27077 11056 -27067
rect 10976 -27087 11056 -27077
rect 11296 -27077 11306 -27067
rect 11366 -27077 11376 -27017
rect 11296 -27087 11376 -27077
rect 10976 -27357 11036 -27087
rect 11116 -27147 11146 -27127
rect 11096 -27187 11146 -27147
rect 11206 -27147 11236 -27127
rect 11206 -27187 11256 -27147
rect 11096 -27257 11256 -27187
rect 11096 -27297 11146 -27257
rect 11116 -27317 11146 -27297
rect 11206 -27297 11256 -27257
rect 11206 -27317 11236 -27297
rect 11316 -27347 11376 -27087
rect 11306 -27357 11376 -27347
rect 10976 -27367 11056 -27357
rect 10976 -27427 10986 -27367
rect 11046 -27377 11056 -27367
rect 11296 -27367 11376 -27357
rect 11296 -27377 11306 -27367
rect 11046 -27427 11306 -27377
rect 11366 -27427 11376 -27367
rect 10976 -27437 11376 -27427
rect 11432 -27017 11832 -27007
rect 11432 -27077 11442 -27017
rect 11502 -27067 11762 -27017
rect 11502 -27077 11512 -27067
rect 11432 -27087 11512 -27077
rect 11752 -27077 11762 -27067
rect 11822 -27077 11832 -27017
rect 11752 -27087 11832 -27077
rect 11432 -27357 11492 -27087
rect 11572 -27147 11602 -27127
rect 11552 -27187 11602 -27147
rect 11662 -27147 11692 -27127
rect 11662 -27187 11712 -27147
rect 11552 -27257 11712 -27187
rect 11552 -27297 11602 -27257
rect 11572 -27317 11602 -27297
rect 11662 -27297 11712 -27257
rect 11662 -27317 11692 -27297
rect 11772 -27347 11832 -27087
rect 11762 -27357 11832 -27347
rect 11432 -27367 11512 -27357
rect 11432 -27427 11442 -27367
rect 11502 -27377 11512 -27367
rect 11752 -27367 11832 -27357
rect 11752 -27377 11762 -27367
rect 11502 -27427 11762 -27377
rect 11822 -27427 11832 -27367
rect 11432 -27437 11832 -27427
rect 11890 -27017 12290 -27007
rect 11890 -27077 11900 -27017
rect 11960 -27067 12220 -27017
rect 11960 -27077 11970 -27067
rect 11890 -27087 11970 -27077
rect 12210 -27077 12220 -27067
rect 12280 -27077 12290 -27017
rect 12210 -27087 12290 -27077
rect 11890 -27357 11950 -27087
rect 12030 -27147 12060 -27127
rect 12010 -27187 12060 -27147
rect 12120 -27147 12150 -27127
rect 12120 -27187 12170 -27147
rect 12010 -27257 12170 -27187
rect 12010 -27297 12060 -27257
rect 12030 -27317 12060 -27297
rect 12120 -27297 12170 -27257
rect 12120 -27317 12150 -27297
rect 12230 -27347 12290 -27087
rect 12220 -27357 12290 -27347
rect 11890 -27367 11970 -27357
rect 11890 -27427 11900 -27367
rect 11960 -27377 11970 -27367
rect 12210 -27367 12290 -27357
rect 12210 -27377 12220 -27367
rect 11960 -27427 12220 -27377
rect 12280 -27427 12290 -27367
rect 11890 -27437 12290 -27427
rect 12346 -27017 12746 -27007
rect 12346 -27077 12356 -27017
rect 12416 -27067 12676 -27017
rect 12416 -27077 12426 -27067
rect 12346 -27087 12426 -27077
rect 12666 -27077 12676 -27067
rect 12736 -27077 12746 -27017
rect 12666 -27087 12746 -27077
rect 12346 -27357 12406 -27087
rect 12486 -27147 12516 -27127
rect 12466 -27187 12516 -27147
rect 12576 -27147 12606 -27127
rect 12576 -27187 12626 -27147
rect 12466 -27257 12626 -27187
rect 12466 -27297 12516 -27257
rect 12486 -27317 12516 -27297
rect 12576 -27297 12626 -27257
rect 12576 -27317 12606 -27297
rect 12686 -27347 12746 -27087
rect 12676 -27357 12746 -27347
rect 12346 -27367 12426 -27357
rect 12346 -27427 12356 -27367
rect 12416 -27377 12426 -27367
rect 12666 -27367 12746 -27357
rect 12666 -27377 12676 -27367
rect 12416 -27427 12676 -27377
rect 12736 -27427 12746 -27367
rect 12346 -27437 12746 -27427
rect 12802 -27017 13202 -27007
rect 12802 -27077 12812 -27017
rect 12872 -27067 13132 -27017
rect 12872 -27077 12882 -27067
rect 12802 -27087 12882 -27077
rect 13122 -27077 13132 -27067
rect 13192 -27077 13202 -27017
rect 13122 -27087 13202 -27077
rect 12802 -27357 12862 -27087
rect 12942 -27147 12972 -27127
rect 12922 -27187 12972 -27147
rect 13032 -27147 13062 -27127
rect 13032 -27187 13082 -27147
rect 12922 -27257 13082 -27187
rect 12922 -27297 12972 -27257
rect 12942 -27317 12972 -27297
rect 13032 -27297 13082 -27257
rect 13032 -27317 13062 -27297
rect 13142 -27347 13202 -27087
rect 13132 -27357 13202 -27347
rect 12802 -27367 12882 -27357
rect 12802 -27427 12812 -27367
rect 12872 -27377 12882 -27367
rect 13122 -27367 13202 -27357
rect 13122 -27377 13132 -27367
rect 12872 -27427 13132 -27377
rect 13192 -27427 13202 -27367
rect 12802 -27437 13202 -27427
rect 13260 -27017 13660 -27007
rect 13260 -27077 13270 -27017
rect 13330 -27067 13590 -27017
rect 13330 -27077 13340 -27067
rect 13260 -27087 13340 -27077
rect 13580 -27077 13590 -27067
rect 13650 -27077 13660 -27017
rect 13580 -27087 13660 -27077
rect 13260 -27357 13320 -27087
rect 13400 -27147 13430 -27127
rect 13380 -27187 13430 -27147
rect 13490 -27147 13520 -27127
rect 13490 -27187 13540 -27147
rect 13380 -27257 13540 -27187
rect 13380 -27297 13430 -27257
rect 13400 -27317 13430 -27297
rect 13490 -27297 13540 -27257
rect 13490 -27317 13520 -27297
rect 13600 -27347 13660 -27087
rect 13590 -27357 13660 -27347
rect 13260 -27367 13340 -27357
rect 13260 -27427 13270 -27367
rect 13330 -27377 13340 -27367
rect 13580 -27367 13660 -27357
rect 13580 -27377 13590 -27367
rect 13330 -27427 13590 -27377
rect 13650 -27427 13660 -27367
rect 13260 -27437 13660 -27427
rect 13716 -27017 14116 -27007
rect 13716 -27077 13726 -27017
rect 13786 -27067 14046 -27017
rect 13786 -27077 13796 -27067
rect 13716 -27087 13796 -27077
rect 14036 -27077 14046 -27067
rect 14106 -27077 14116 -27017
rect 14036 -27087 14116 -27077
rect 13716 -27357 13776 -27087
rect 13856 -27147 13886 -27127
rect 13836 -27187 13886 -27147
rect 13946 -27147 13976 -27127
rect 13946 -27187 13996 -27147
rect 13836 -27257 13996 -27187
rect 13836 -27297 13886 -27257
rect 13856 -27317 13886 -27297
rect 13946 -27297 13996 -27257
rect 13946 -27317 13976 -27297
rect 14056 -27347 14116 -27087
rect 14046 -27357 14116 -27347
rect 13716 -27367 13796 -27357
rect 13716 -27427 13726 -27367
rect 13786 -27377 13796 -27367
rect 14036 -27367 14116 -27357
rect 14036 -27377 14046 -27367
rect 13786 -27427 14046 -27377
rect 14106 -27427 14116 -27367
rect 13716 -27437 14116 -27427
rect 14172 -27017 14572 -27007
rect 14172 -27077 14182 -27017
rect 14242 -27067 14502 -27017
rect 14242 -27077 14252 -27067
rect 14172 -27087 14252 -27077
rect 14492 -27077 14502 -27067
rect 14562 -27077 14572 -27017
rect 14492 -27087 14572 -27077
rect 14172 -27357 14232 -27087
rect 14312 -27147 14342 -27127
rect 14292 -27187 14342 -27147
rect 14402 -27147 14432 -27127
rect 14402 -27187 14452 -27147
rect 14292 -27257 14452 -27187
rect 14292 -27297 14342 -27257
rect 14312 -27317 14342 -27297
rect 14402 -27297 14452 -27257
rect 14402 -27317 14432 -27297
rect 14512 -27347 14572 -27087
rect 14502 -27357 14572 -27347
rect 14172 -27367 14252 -27357
rect 14172 -27427 14182 -27367
rect 14242 -27377 14252 -27367
rect 14492 -27367 14572 -27357
rect 14492 -27377 14502 -27367
rect 14242 -27427 14502 -27377
rect 14562 -27427 14572 -27367
rect 14172 -27437 14572 -27427
rect 14630 -27017 15030 -27007
rect 14630 -27077 14640 -27017
rect 14700 -27067 14960 -27017
rect 14700 -27077 14710 -27067
rect 14630 -27087 14710 -27077
rect 14950 -27077 14960 -27067
rect 15020 -27077 15030 -27017
rect 14950 -27087 15030 -27077
rect 14630 -27357 14690 -27087
rect 14770 -27147 14800 -27127
rect 14750 -27187 14800 -27147
rect 14860 -27147 14890 -27127
rect 14860 -27187 14910 -27147
rect 14750 -27257 14910 -27187
rect 14750 -27297 14800 -27257
rect 14770 -27317 14800 -27297
rect 14860 -27297 14910 -27257
rect 14860 -27317 14890 -27297
rect 14970 -27347 15030 -27087
rect 14960 -27357 15030 -27347
rect 14630 -27367 14710 -27357
rect 14630 -27427 14640 -27367
rect 14700 -27377 14710 -27367
rect 14950 -27367 15030 -27357
rect 14950 -27377 14960 -27367
rect 14700 -27427 14960 -27377
rect 15020 -27427 15030 -27367
rect 14630 -27437 15030 -27427
rect 15086 -27017 15486 -27007
rect 15086 -27077 15096 -27017
rect 15156 -27067 15416 -27017
rect 15156 -27077 15166 -27067
rect 15086 -27087 15166 -27077
rect 15406 -27077 15416 -27067
rect 15476 -27077 15486 -27017
rect 15406 -27087 15486 -27077
rect 15086 -27357 15146 -27087
rect 15226 -27147 15256 -27127
rect 15206 -27187 15256 -27147
rect 15316 -27147 15346 -27127
rect 15316 -27187 15366 -27147
rect 15206 -27257 15366 -27187
rect 15206 -27297 15256 -27257
rect 15226 -27317 15256 -27297
rect 15316 -27297 15366 -27257
rect 15316 -27317 15346 -27297
rect 15426 -27347 15486 -27087
rect 15416 -27357 15486 -27347
rect 15086 -27367 15166 -27357
rect 15086 -27427 15096 -27367
rect 15156 -27377 15166 -27367
rect 15406 -27367 15486 -27357
rect 15406 -27377 15416 -27367
rect 15156 -27427 15416 -27377
rect 15476 -27427 15486 -27367
rect 15086 -27437 15486 -27427
rect 0 -27533 400 -27523
rect 0 -27593 10 -27533
rect 70 -27583 330 -27533
rect 70 -27593 80 -27583
rect 0 -27603 80 -27593
rect 320 -27593 330 -27583
rect 390 -27593 400 -27533
rect 320 -27603 400 -27593
rect 0 -27873 60 -27603
rect 140 -27663 170 -27643
rect 120 -27703 170 -27663
rect 230 -27663 260 -27643
rect 230 -27703 280 -27663
rect 120 -27773 280 -27703
rect 120 -27813 170 -27773
rect 140 -27833 170 -27813
rect 230 -27813 280 -27773
rect 230 -27833 260 -27813
rect 340 -27863 400 -27603
rect 330 -27873 400 -27863
rect 0 -27883 80 -27873
rect 0 -27943 10 -27883
rect 70 -27893 80 -27883
rect 320 -27883 400 -27873
rect 320 -27893 330 -27883
rect 70 -27943 330 -27893
rect 390 -27943 400 -27883
rect 0 -27953 400 -27943
rect 456 -27533 856 -27523
rect 456 -27593 466 -27533
rect 526 -27583 786 -27533
rect 526 -27593 536 -27583
rect 456 -27603 536 -27593
rect 776 -27593 786 -27583
rect 846 -27593 856 -27533
rect 776 -27603 856 -27593
rect 456 -27873 516 -27603
rect 596 -27663 626 -27643
rect 576 -27703 626 -27663
rect 686 -27663 716 -27643
rect 686 -27703 736 -27663
rect 576 -27773 736 -27703
rect 576 -27813 626 -27773
rect 596 -27833 626 -27813
rect 686 -27813 736 -27773
rect 686 -27833 716 -27813
rect 796 -27863 856 -27603
rect 786 -27873 856 -27863
rect 456 -27883 536 -27873
rect 456 -27943 466 -27883
rect 526 -27893 536 -27883
rect 776 -27883 856 -27873
rect 776 -27893 786 -27883
rect 526 -27943 786 -27893
rect 846 -27943 856 -27883
rect 456 -27953 856 -27943
rect 912 -27533 1312 -27523
rect 912 -27593 922 -27533
rect 982 -27583 1242 -27533
rect 982 -27593 992 -27583
rect 912 -27603 992 -27593
rect 1232 -27593 1242 -27583
rect 1302 -27593 1312 -27533
rect 1232 -27603 1312 -27593
rect 912 -27873 972 -27603
rect 1052 -27663 1082 -27643
rect 1032 -27703 1082 -27663
rect 1142 -27663 1172 -27643
rect 1142 -27703 1192 -27663
rect 1032 -27773 1192 -27703
rect 1032 -27813 1082 -27773
rect 1052 -27833 1082 -27813
rect 1142 -27813 1192 -27773
rect 1142 -27833 1172 -27813
rect 1252 -27863 1312 -27603
rect 1242 -27873 1312 -27863
rect 912 -27883 992 -27873
rect 912 -27943 922 -27883
rect 982 -27893 992 -27883
rect 1232 -27883 1312 -27873
rect 1232 -27893 1242 -27883
rect 982 -27943 1242 -27893
rect 1302 -27943 1312 -27883
rect 912 -27953 1312 -27943
rect 1370 -27533 1770 -27523
rect 1370 -27593 1380 -27533
rect 1440 -27583 1700 -27533
rect 1440 -27593 1450 -27583
rect 1370 -27603 1450 -27593
rect 1690 -27593 1700 -27583
rect 1760 -27593 1770 -27533
rect 1690 -27603 1770 -27593
rect 1370 -27873 1430 -27603
rect 1510 -27663 1540 -27643
rect 1490 -27703 1540 -27663
rect 1600 -27663 1630 -27643
rect 1600 -27703 1650 -27663
rect 1490 -27773 1650 -27703
rect 1490 -27813 1540 -27773
rect 1510 -27833 1540 -27813
rect 1600 -27813 1650 -27773
rect 1600 -27833 1630 -27813
rect 1710 -27863 1770 -27603
rect 1700 -27873 1770 -27863
rect 1370 -27883 1450 -27873
rect 1370 -27943 1380 -27883
rect 1440 -27893 1450 -27883
rect 1690 -27883 1770 -27873
rect 1690 -27893 1700 -27883
rect 1440 -27943 1700 -27893
rect 1760 -27943 1770 -27883
rect 1370 -27953 1770 -27943
rect 1826 -27533 2226 -27523
rect 1826 -27593 1836 -27533
rect 1896 -27583 2156 -27533
rect 1896 -27593 1906 -27583
rect 1826 -27603 1906 -27593
rect 2146 -27593 2156 -27583
rect 2216 -27593 2226 -27533
rect 2146 -27603 2226 -27593
rect 1826 -27873 1886 -27603
rect 1966 -27663 1996 -27643
rect 1946 -27703 1996 -27663
rect 2056 -27663 2086 -27643
rect 2056 -27703 2106 -27663
rect 1946 -27773 2106 -27703
rect 1946 -27813 1996 -27773
rect 1966 -27833 1996 -27813
rect 2056 -27813 2106 -27773
rect 2056 -27833 2086 -27813
rect 2166 -27863 2226 -27603
rect 2156 -27873 2226 -27863
rect 1826 -27883 1906 -27873
rect 1826 -27943 1836 -27883
rect 1896 -27893 1906 -27883
rect 2146 -27883 2226 -27873
rect 2146 -27893 2156 -27883
rect 1896 -27943 2156 -27893
rect 2216 -27943 2226 -27883
rect 1826 -27953 2226 -27943
rect 2282 -27533 2682 -27523
rect 2282 -27593 2292 -27533
rect 2352 -27583 2612 -27533
rect 2352 -27593 2362 -27583
rect 2282 -27603 2362 -27593
rect 2602 -27593 2612 -27583
rect 2672 -27593 2682 -27533
rect 2602 -27603 2682 -27593
rect 2282 -27873 2342 -27603
rect 2422 -27663 2452 -27643
rect 2402 -27703 2452 -27663
rect 2512 -27663 2542 -27643
rect 2512 -27703 2562 -27663
rect 2402 -27773 2562 -27703
rect 2402 -27813 2452 -27773
rect 2422 -27833 2452 -27813
rect 2512 -27813 2562 -27773
rect 2512 -27833 2542 -27813
rect 2622 -27863 2682 -27603
rect 2612 -27873 2682 -27863
rect 2282 -27883 2362 -27873
rect 2282 -27943 2292 -27883
rect 2352 -27893 2362 -27883
rect 2602 -27883 2682 -27873
rect 2602 -27893 2612 -27883
rect 2352 -27943 2612 -27893
rect 2672 -27943 2682 -27883
rect 2282 -27953 2682 -27943
rect 2740 -27533 3140 -27523
rect 2740 -27593 2750 -27533
rect 2810 -27583 3070 -27533
rect 2810 -27593 2820 -27583
rect 2740 -27603 2820 -27593
rect 3060 -27593 3070 -27583
rect 3130 -27593 3140 -27533
rect 3060 -27603 3140 -27593
rect 2740 -27873 2800 -27603
rect 2880 -27663 2910 -27643
rect 2860 -27703 2910 -27663
rect 2970 -27663 3000 -27643
rect 2970 -27703 3020 -27663
rect 2860 -27773 3020 -27703
rect 2860 -27813 2910 -27773
rect 2880 -27833 2910 -27813
rect 2970 -27813 3020 -27773
rect 2970 -27833 3000 -27813
rect 3080 -27863 3140 -27603
rect 3070 -27873 3140 -27863
rect 2740 -27883 2820 -27873
rect 2740 -27943 2750 -27883
rect 2810 -27893 2820 -27883
rect 3060 -27883 3140 -27873
rect 3060 -27893 3070 -27883
rect 2810 -27943 3070 -27893
rect 3130 -27943 3140 -27883
rect 2740 -27953 3140 -27943
rect 3196 -27533 3596 -27523
rect 3196 -27593 3206 -27533
rect 3266 -27583 3526 -27533
rect 3266 -27593 3276 -27583
rect 3196 -27603 3276 -27593
rect 3516 -27593 3526 -27583
rect 3586 -27593 3596 -27533
rect 3516 -27603 3596 -27593
rect 3196 -27873 3256 -27603
rect 3336 -27663 3366 -27643
rect 3316 -27703 3366 -27663
rect 3426 -27663 3456 -27643
rect 3426 -27703 3476 -27663
rect 3316 -27773 3476 -27703
rect 3316 -27813 3366 -27773
rect 3336 -27833 3366 -27813
rect 3426 -27813 3476 -27773
rect 3426 -27833 3456 -27813
rect 3536 -27863 3596 -27603
rect 3526 -27873 3596 -27863
rect 3196 -27883 3276 -27873
rect 3196 -27943 3206 -27883
rect 3266 -27893 3276 -27883
rect 3516 -27883 3596 -27873
rect 3516 -27893 3526 -27883
rect 3266 -27943 3526 -27893
rect 3586 -27943 3596 -27883
rect 3196 -27953 3596 -27943
rect 3652 -27533 4052 -27523
rect 3652 -27593 3662 -27533
rect 3722 -27583 3982 -27533
rect 3722 -27593 3732 -27583
rect 3652 -27603 3732 -27593
rect 3972 -27593 3982 -27583
rect 4042 -27593 4052 -27533
rect 3972 -27603 4052 -27593
rect 3652 -27873 3712 -27603
rect 3792 -27663 3822 -27643
rect 3772 -27703 3822 -27663
rect 3882 -27663 3912 -27643
rect 3882 -27703 3932 -27663
rect 3772 -27773 3932 -27703
rect 3772 -27813 3822 -27773
rect 3792 -27833 3822 -27813
rect 3882 -27813 3932 -27773
rect 3882 -27833 3912 -27813
rect 3992 -27863 4052 -27603
rect 3982 -27873 4052 -27863
rect 3652 -27883 3732 -27873
rect 3652 -27943 3662 -27883
rect 3722 -27893 3732 -27883
rect 3972 -27883 4052 -27873
rect 3972 -27893 3982 -27883
rect 3722 -27943 3982 -27893
rect 4042 -27943 4052 -27883
rect 3652 -27953 4052 -27943
rect 4110 -27533 4510 -27523
rect 4110 -27593 4120 -27533
rect 4180 -27583 4440 -27533
rect 4180 -27593 4190 -27583
rect 4110 -27603 4190 -27593
rect 4430 -27593 4440 -27583
rect 4500 -27593 4510 -27533
rect 4430 -27603 4510 -27593
rect 4110 -27873 4170 -27603
rect 4250 -27663 4280 -27643
rect 4230 -27703 4280 -27663
rect 4340 -27663 4370 -27643
rect 4340 -27703 4390 -27663
rect 4230 -27773 4390 -27703
rect 4230 -27813 4280 -27773
rect 4250 -27833 4280 -27813
rect 4340 -27813 4390 -27773
rect 4340 -27833 4370 -27813
rect 4450 -27863 4510 -27603
rect 4440 -27873 4510 -27863
rect 4110 -27883 4190 -27873
rect 4110 -27943 4120 -27883
rect 4180 -27893 4190 -27883
rect 4430 -27883 4510 -27873
rect 4430 -27893 4440 -27883
rect 4180 -27943 4440 -27893
rect 4500 -27943 4510 -27883
rect 4110 -27953 4510 -27943
rect 4566 -27533 4966 -27523
rect 4566 -27593 4576 -27533
rect 4636 -27583 4896 -27533
rect 4636 -27593 4646 -27583
rect 4566 -27603 4646 -27593
rect 4886 -27593 4896 -27583
rect 4956 -27593 4966 -27533
rect 4886 -27603 4966 -27593
rect 4566 -27873 4626 -27603
rect 4706 -27663 4736 -27643
rect 4686 -27703 4736 -27663
rect 4796 -27663 4826 -27643
rect 4796 -27703 4846 -27663
rect 4686 -27773 4846 -27703
rect 4686 -27813 4736 -27773
rect 4706 -27833 4736 -27813
rect 4796 -27813 4846 -27773
rect 4796 -27833 4826 -27813
rect 4906 -27863 4966 -27603
rect 4896 -27873 4966 -27863
rect 4566 -27883 4646 -27873
rect 4566 -27943 4576 -27883
rect 4636 -27893 4646 -27883
rect 4886 -27883 4966 -27873
rect 4886 -27893 4896 -27883
rect 4636 -27943 4896 -27893
rect 4956 -27943 4966 -27883
rect 4566 -27953 4966 -27943
rect 5022 -27533 5422 -27523
rect 5022 -27593 5032 -27533
rect 5092 -27583 5352 -27533
rect 5092 -27593 5102 -27583
rect 5022 -27603 5102 -27593
rect 5342 -27593 5352 -27583
rect 5412 -27593 5422 -27533
rect 5342 -27603 5422 -27593
rect 5022 -27873 5082 -27603
rect 5162 -27663 5192 -27643
rect 5142 -27703 5192 -27663
rect 5252 -27663 5282 -27643
rect 5252 -27703 5302 -27663
rect 5142 -27773 5302 -27703
rect 5142 -27813 5192 -27773
rect 5162 -27833 5192 -27813
rect 5252 -27813 5302 -27773
rect 5252 -27833 5282 -27813
rect 5362 -27863 5422 -27603
rect 5352 -27873 5422 -27863
rect 5022 -27883 5102 -27873
rect 5022 -27943 5032 -27883
rect 5092 -27893 5102 -27883
rect 5342 -27883 5422 -27873
rect 5342 -27893 5352 -27883
rect 5092 -27943 5352 -27893
rect 5412 -27943 5422 -27883
rect 5022 -27953 5422 -27943
rect 5480 -27533 5880 -27523
rect 5480 -27593 5490 -27533
rect 5550 -27583 5810 -27533
rect 5550 -27593 5560 -27583
rect 5480 -27603 5560 -27593
rect 5800 -27593 5810 -27583
rect 5870 -27593 5880 -27533
rect 5800 -27603 5880 -27593
rect 5480 -27873 5540 -27603
rect 5620 -27663 5650 -27643
rect 5600 -27703 5650 -27663
rect 5710 -27663 5740 -27643
rect 5710 -27703 5760 -27663
rect 5600 -27773 5760 -27703
rect 5600 -27813 5650 -27773
rect 5620 -27833 5650 -27813
rect 5710 -27813 5760 -27773
rect 5710 -27833 5740 -27813
rect 5820 -27863 5880 -27603
rect 5810 -27873 5880 -27863
rect 5480 -27883 5560 -27873
rect 5480 -27943 5490 -27883
rect 5550 -27893 5560 -27883
rect 5800 -27883 5880 -27873
rect 5800 -27893 5810 -27883
rect 5550 -27943 5810 -27893
rect 5870 -27943 5880 -27883
rect 5480 -27953 5880 -27943
rect 5936 -27533 6336 -27523
rect 5936 -27593 5946 -27533
rect 6006 -27583 6266 -27533
rect 6006 -27593 6016 -27583
rect 5936 -27603 6016 -27593
rect 6256 -27593 6266 -27583
rect 6326 -27593 6336 -27533
rect 6256 -27603 6336 -27593
rect 5936 -27873 5996 -27603
rect 6076 -27663 6106 -27643
rect 6056 -27703 6106 -27663
rect 6166 -27663 6196 -27643
rect 6166 -27703 6216 -27663
rect 6056 -27773 6216 -27703
rect 6056 -27813 6106 -27773
rect 6076 -27833 6106 -27813
rect 6166 -27813 6216 -27773
rect 6166 -27833 6196 -27813
rect 6276 -27863 6336 -27603
rect 6266 -27873 6336 -27863
rect 5936 -27883 6016 -27873
rect 5936 -27943 5946 -27883
rect 6006 -27893 6016 -27883
rect 6256 -27883 6336 -27873
rect 6256 -27893 6266 -27883
rect 6006 -27943 6266 -27893
rect 6326 -27943 6336 -27883
rect 5936 -27953 6336 -27943
rect 6392 -27533 6792 -27523
rect 6392 -27593 6402 -27533
rect 6462 -27583 6722 -27533
rect 6462 -27593 6472 -27583
rect 6392 -27603 6472 -27593
rect 6712 -27593 6722 -27583
rect 6782 -27593 6792 -27533
rect 6712 -27603 6792 -27593
rect 6392 -27873 6452 -27603
rect 6532 -27663 6562 -27643
rect 6512 -27703 6562 -27663
rect 6622 -27663 6652 -27643
rect 6622 -27703 6672 -27663
rect 6512 -27773 6672 -27703
rect 6512 -27813 6562 -27773
rect 6532 -27833 6562 -27813
rect 6622 -27813 6672 -27773
rect 6622 -27833 6652 -27813
rect 6732 -27863 6792 -27603
rect 6722 -27873 6792 -27863
rect 6392 -27883 6472 -27873
rect 6392 -27943 6402 -27883
rect 6462 -27893 6472 -27883
rect 6712 -27883 6792 -27873
rect 6712 -27893 6722 -27883
rect 6462 -27943 6722 -27893
rect 6782 -27943 6792 -27883
rect 6392 -27953 6792 -27943
rect 6850 -27533 7250 -27523
rect 6850 -27593 6860 -27533
rect 6920 -27583 7180 -27533
rect 6920 -27593 6930 -27583
rect 6850 -27603 6930 -27593
rect 7170 -27593 7180 -27583
rect 7240 -27593 7250 -27533
rect 7170 -27603 7250 -27593
rect 6850 -27873 6910 -27603
rect 6990 -27663 7020 -27643
rect 6970 -27703 7020 -27663
rect 7080 -27663 7110 -27643
rect 7080 -27703 7130 -27663
rect 6970 -27773 7130 -27703
rect 6970 -27813 7020 -27773
rect 6990 -27833 7020 -27813
rect 7080 -27813 7130 -27773
rect 7080 -27833 7110 -27813
rect 7190 -27863 7250 -27603
rect 7180 -27873 7250 -27863
rect 6850 -27883 6930 -27873
rect 6850 -27943 6860 -27883
rect 6920 -27893 6930 -27883
rect 7170 -27883 7250 -27873
rect 7170 -27893 7180 -27883
rect 6920 -27943 7180 -27893
rect 7240 -27943 7250 -27883
rect 6850 -27953 7250 -27943
rect 7306 -27533 7706 -27523
rect 7306 -27593 7316 -27533
rect 7376 -27583 7636 -27533
rect 7376 -27593 7386 -27583
rect 7306 -27603 7386 -27593
rect 7626 -27593 7636 -27583
rect 7696 -27593 7706 -27533
rect 7626 -27603 7706 -27593
rect 7306 -27873 7366 -27603
rect 7446 -27663 7476 -27643
rect 7426 -27703 7476 -27663
rect 7536 -27663 7566 -27643
rect 7536 -27703 7586 -27663
rect 7426 -27773 7586 -27703
rect 7426 -27813 7476 -27773
rect 7446 -27833 7476 -27813
rect 7536 -27813 7586 -27773
rect 7536 -27833 7566 -27813
rect 7646 -27863 7706 -27603
rect 7636 -27873 7706 -27863
rect 7306 -27883 7386 -27873
rect 7306 -27943 7316 -27883
rect 7376 -27893 7386 -27883
rect 7626 -27883 7706 -27873
rect 7626 -27893 7636 -27883
rect 7376 -27943 7636 -27893
rect 7696 -27943 7706 -27883
rect 7306 -27953 7706 -27943
rect 7762 -27533 8162 -27523
rect 7762 -27593 7772 -27533
rect 7832 -27583 8092 -27533
rect 7832 -27593 7842 -27583
rect 7762 -27603 7842 -27593
rect 8082 -27593 8092 -27583
rect 8152 -27593 8162 -27533
rect 8082 -27603 8162 -27593
rect 7762 -27873 7822 -27603
rect 7902 -27663 7932 -27643
rect 7882 -27703 7932 -27663
rect 7992 -27663 8022 -27643
rect 7992 -27703 8042 -27663
rect 7882 -27773 8042 -27703
rect 7882 -27813 7932 -27773
rect 7902 -27833 7932 -27813
rect 7992 -27813 8042 -27773
rect 7992 -27833 8022 -27813
rect 8102 -27863 8162 -27603
rect 8092 -27873 8162 -27863
rect 7762 -27883 7842 -27873
rect 7762 -27943 7772 -27883
rect 7832 -27893 7842 -27883
rect 8082 -27883 8162 -27873
rect 8082 -27893 8092 -27883
rect 7832 -27943 8092 -27893
rect 8152 -27943 8162 -27883
rect 7762 -27953 8162 -27943
rect 8236 -27533 8636 -27523
rect 8236 -27593 8246 -27533
rect 8306 -27583 8566 -27533
rect 8306 -27593 8316 -27583
rect 8236 -27603 8316 -27593
rect 8556 -27593 8566 -27583
rect 8626 -27593 8636 -27533
rect 8556 -27603 8636 -27593
rect 8236 -27873 8296 -27603
rect 8376 -27663 8406 -27643
rect 8356 -27703 8406 -27663
rect 8466 -27663 8496 -27643
rect 8466 -27703 8516 -27663
rect 8356 -27773 8516 -27703
rect 8356 -27813 8406 -27773
rect 8376 -27833 8406 -27813
rect 8466 -27813 8516 -27773
rect 8466 -27833 8496 -27813
rect 8576 -27863 8636 -27603
rect 8566 -27873 8636 -27863
rect 8236 -27883 8316 -27873
rect 8236 -27943 8246 -27883
rect 8306 -27893 8316 -27883
rect 8556 -27883 8636 -27873
rect 8556 -27893 8566 -27883
rect 8306 -27943 8566 -27893
rect 8626 -27943 8636 -27883
rect 8236 -27953 8636 -27943
rect 8692 -27533 9092 -27523
rect 8692 -27593 8702 -27533
rect 8762 -27583 9022 -27533
rect 8762 -27593 8772 -27583
rect 8692 -27603 8772 -27593
rect 9012 -27593 9022 -27583
rect 9082 -27593 9092 -27533
rect 9012 -27603 9092 -27593
rect 8692 -27873 8752 -27603
rect 8832 -27663 8862 -27643
rect 8812 -27703 8862 -27663
rect 8922 -27663 8952 -27643
rect 8922 -27703 8972 -27663
rect 8812 -27773 8972 -27703
rect 8812 -27813 8862 -27773
rect 8832 -27833 8862 -27813
rect 8922 -27813 8972 -27773
rect 8922 -27833 8952 -27813
rect 9032 -27863 9092 -27603
rect 9022 -27873 9092 -27863
rect 8692 -27883 8772 -27873
rect 8692 -27943 8702 -27883
rect 8762 -27893 8772 -27883
rect 9012 -27883 9092 -27873
rect 9012 -27893 9022 -27883
rect 8762 -27943 9022 -27893
rect 9082 -27943 9092 -27883
rect 8692 -27953 9092 -27943
rect 9150 -27533 9550 -27523
rect 9150 -27593 9160 -27533
rect 9220 -27583 9480 -27533
rect 9220 -27593 9230 -27583
rect 9150 -27603 9230 -27593
rect 9470 -27593 9480 -27583
rect 9540 -27593 9550 -27533
rect 9470 -27603 9550 -27593
rect 9150 -27873 9210 -27603
rect 9290 -27663 9320 -27643
rect 9270 -27703 9320 -27663
rect 9380 -27663 9410 -27643
rect 9380 -27703 9430 -27663
rect 9270 -27773 9430 -27703
rect 9270 -27813 9320 -27773
rect 9290 -27833 9320 -27813
rect 9380 -27813 9430 -27773
rect 9380 -27833 9410 -27813
rect 9490 -27863 9550 -27603
rect 9480 -27873 9550 -27863
rect 9150 -27883 9230 -27873
rect 9150 -27943 9160 -27883
rect 9220 -27893 9230 -27883
rect 9470 -27883 9550 -27873
rect 9470 -27893 9480 -27883
rect 9220 -27943 9480 -27893
rect 9540 -27943 9550 -27883
rect 9150 -27953 9550 -27943
rect 9606 -27533 10006 -27523
rect 9606 -27593 9616 -27533
rect 9676 -27583 9936 -27533
rect 9676 -27593 9686 -27583
rect 9606 -27603 9686 -27593
rect 9926 -27593 9936 -27583
rect 9996 -27593 10006 -27533
rect 9926 -27603 10006 -27593
rect 9606 -27873 9666 -27603
rect 9746 -27663 9776 -27643
rect 9726 -27703 9776 -27663
rect 9836 -27663 9866 -27643
rect 9836 -27703 9886 -27663
rect 9726 -27773 9886 -27703
rect 9726 -27813 9776 -27773
rect 9746 -27833 9776 -27813
rect 9836 -27813 9886 -27773
rect 9836 -27833 9866 -27813
rect 9946 -27863 10006 -27603
rect 9936 -27873 10006 -27863
rect 9606 -27883 9686 -27873
rect 9606 -27943 9616 -27883
rect 9676 -27893 9686 -27883
rect 9926 -27883 10006 -27873
rect 9926 -27893 9936 -27883
rect 9676 -27943 9936 -27893
rect 9996 -27943 10006 -27883
rect 9606 -27953 10006 -27943
rect 10062 -27533 10462 -27523
rect 10062 -27593 10072 -27533
rect 10132 -27583 10392 -27533
rect 10132 -27593 10142 -27583
rect 10062 -27603 10142 -27593
rect 10382 -27593 10392 -27583
rect 10452 -27593 10462 -27533
rect 10382 -27603 10462 -27593
rect 10062 -27873 10122 -27603
rect 10202 -27663 10232 -27643
rect 10182 -27703 10232 -27663
rect 10292 -27663 10322 -27643
rect 10292 -27703 10342 -27663
rect 10182 -27773 10342 -27703
rect 10182 -27813 10232 -27773
rect 10202 -27833 10232 -27813
rect 10292 -27813 10342 -27773
rect 10292 -27833 10322 -27813
rect 10402 -27863 10462 -27603
rect 10392 -27873 10462 -27863
rect 10062 -27883 10142 -27873
rect 10062 -27943 10072 -27883
rect 10132 -27893 10142 -27883
rect 10382 -27883 10462 -27873
rect 10382 -27893 10392 -27883
rect 10132 -27943 10392 -27893
rect 10452 -27943 10462 -27883
rect 10062 -27953 10462 -27943
rect 10520 -27533 10920 -27523
rect 10520 -27593 10530 -27533
rect 10590 -27583 10850 -27533
rect 10590 -27593 10600 -27583
rect 10520 -27603 10600 -27593
rect 10840 -27593 10850 -27583
rect 10910 -27593 10920 -27533
rect 10840 -27603 10920 -27593
rect 10520 -27873 10580 -27603
rect 10660 -27663 10690 -27643
rect 10640 -27703 10690 -27663
rect 10750 -27663 10780 -27643
rect 10750 -27703 10800 -27663
rect 10640 -27773 10800 -27703
rect 10640 -27813 10690 -27773
rect 10660 -27833 10690 -27813
rect 10750 -27813 10800 -27773
rect 10750 -27833 10780 -27813
rect 10860 -27863 10920 -27603
rect 10850 -27873 10920 -27863
rect 10520 -27883 10600 -27873
rect 10520 -27943 10530 -27883
rect 10590 -27893 10600 -27883
rect 10840 -27883 10920 -27873
rect 10840 -27893 10850 -27883
rect 10590 -27943 10850 -27893
rect 10910 -27943 10920 -27883
rect 10520 -27953 10920 -27943
rect 10976 -27533 11376 -27523
rect 10976 -27593 10986 -27533
rect 11046 -27583 11306 -27533
rect 11046 -27593 11056 -27583
rect 10976 -27603 11056 -27593
rect 11296 -27593 11306 -27583
rect 11366 -27593 11376 -27533
rect 11296 -27603 11376 -27593
rect 10976 -27873 11036 -27603
rect 11116 -27663 11146 -27643
rect 11096 -27703 11146 -27663
rect 11206 -27663 11236 -27643
rect 11206 -27703 11256 -27663
rect 11096 -27773 11256 -27703
rect 11096 -27813 11146 -27773
rect 11116 -27833 11146 -27813
rect 11206 -27813 11256 -27773
rect 11206 -27833 11236 -27813
rect 11316 -27863 11376 -27603
rect 11306 -27873 11376 -27863
rect 10976 -27883 11056 -27873
rect 10976 -27943 10986 -27883
rect 11046 -27893 11056 -27883
rect 11296 -27883 11376 -27873
rect 11296 -27893 11306 -27883
rect 11046 -27943 11306 -27893
rect 11366 -27943 11376 -27883
rect 10976 -27953 11376 -27943
rect 11432 -27533 11832 -27523
rect 11432 -27593 11442 -27533
rect 11502 -27583 11762 -27533
rect 11502 -27593 11512 -27583
rect 11432 -27603 11512 -27593
rect 11752 -27593 11762 -27583
rect 11822 -27593 11832 -27533
rect 11752 -27603 11832 -27593
rect 11432 -27873 11492 -27603
rect 11572 -27663 11602 -27643
rect 11552 -27703 11602 -27663
rect 11662 -27663 11692 -27643
rect 11662 -27703 11712 -27663
rect 11552 -27773 11712 -27703
rect 11552 -27813 11602 -27773
rect 11572 -27833 11602 -27813
rect 11662 -27813 11712 -27773
rect 11662 -27833 11692 -27813
rect 11772 -27863 11832 -27603
rect 11762 -27873 11832 -27863
rect 11432 -27883 11512 -27873
rect 11432 -27943 11442 -27883
rect 11502 -27893 11512 -27883
rect 11752 -27883 11832 -27873
rect 11752 -27893 11762 -27883
rect 11502 -27943 11762 -27893
rect 11822 -27943 11832 -27883
rect 11432 -27953 11832 -27943
rect 11890 -27533 12290 -27523
rect 11890 -27593 11900 -27533
rect 11960 -27583 12220 -27533
rect 11960 -27593 11970 -27583
rect 11890 -27603 11970 -27593
rect 12210 -27593 12220 -27583
rect 12280 -27593 12290 -27533
rect 12210 -27603 12290 -27593
rect 11890 -27873 11950 -27603
rect 12030 -27663 12060 -27643
rect 12010 -27703 12060 -27663
rect 12120 -27663 12150 -27643
rect 12120 -27703 12170 -27663
rect 12010 -27773 12170 -27703
rect 12010 -27813 12060 -27773
rect 12030 -27833 12060 -27813
rect 12120 -27813 12170 -27773
rect 12120 -27833 12150 -27813
rect 12230 -27863 12290 -27603
rect 12220 -27873 12290 -27863
rect 11890 -27883 11970 -27873
rect 11890 -27943 11900 -27883
rect 11960 -27893 11970 -27883
rect 12210 -27883 12290 -27873
rect 12210 -27893 12220 -27883
rect 11960 -27943 12220 -27893
rect 12280 -27943 12290 -27883
rect 11890 -27953 12290 -27943
rect 12346 -27533 12746 -27523
rect 12346 -27593 12356 -27533
rect 12416 -27583 12676 -27533
rect 12416 -27593 12426 -27583
rect 12346 -27603 12426 -27593
rect 12666 -27593 12676 -27583
rect 12736 -27593 12746 -27533
rect 12666 -27603 12746 -27593
rect 12346 -27873 12406 -27603
rect 12486 -27663 12516 -27643
rect 12466 -27703 12516 -27663
rect 12576 -27663 12606 -27643
rect 12576 -27703 12626 -27663
rect 12466 -27773 12626 -27703
rect 12466 -27813 12516 -27773
rect 12486 -27833 12516 -27813
rect 12576 -27813 12626 -27773
rect 12576 -27833 12606 -27813
rect 12686 -27863 12746 -27603
rect 12676 -27873 12746 -27863
rect 12346 -27883 12426 -27873
rect 12346 -27943 12356 -27883
rect 12416 -27893 12426 -27883
rect 12666 -27883 12746 -27873
rect 12666 -27893 12676 -27883
rect 12416 -27943 12676 -27893
rect 12736 -27943 12746 -27883
rect 12346 -27953 12746 -27943
rect 12802 -27533 13202 -27523
rect 12802 -27593 12812 -27533
rect 12872 -27583 13132 -27533
rect 12872 -27593 12882 -27583
rect 12802 -27603 12882 -27593
rect 13122 -27593 13132 -27583
rect 13192 -27593 13202 -27533
rect 13122 -27603 13202 -27593
rect 12802 -27873 12862 -27603
rect 12942 -27663 12972 -27643
rect 12922 -27703 12972 -27663
rect 13032 -27663 13062 -27643
rect 13032 -27703 13082 -27663
rect 12922 -27773 13082 -27703
rect 12922 -27813 12972 -27773
rect 12942 -27833 12972 -27813
rect 13032 -27813 13082 -27773
rect 13032 -27833 13062 -27813
rect 13142 -27863 13202 -27603
rect 13132 -27873 13202 -27863
rect 12802 -27883 12882 -27873
rect 12802 -27943 12812 -27883
rect 12872 -27893 12882 -27883
rect 13122 -27883 13202 -27873
rect 13122 -27893 13132 -27883
rect 12872 -27943 13132 -27893
rect 13192 -27943 13202 -27883
rect 12802 -27953 13202 -27943
rect 13260 -27533 13660 -27523
rect 13260 -27593 13270 -27533
rect 13330 -27583 13590 -27533
rect 13330 -27593 13340 -27583
rect 13260 -27603 13340 -27593
rect 13580 -27593 13590 -27583
rect 13650 -27593 13660 -27533
rect 13580 -27603 13660 -27593
rect 13260 -27873 13320 -27603
rect 13400 -27663 13430 -27643
rect 13380 -27703 13430 -27663
rect 13490 -27663 13520 -27643
rect 13490 -27703 13540 -27663
rect 13380 -27773 13540 -27703
rect 13380 -27813 13430 -27773
rect 13400 -27833 13430 -27813
rect 13490 -27813 13540 -27773
rect 13490 -27833 13520 -27813
rect 13600 -27863 13660 -27603
rect 13590 -27873 13660 -27863
rect 13260 -27883 13340 -27873
rect 13260 -27943 13270 -27883
rect 13330 -27893 13340 -27883
rect 13580 -27883 13660 -27873
rect 13580 -27893 13590 -27883
rect 13330 -27943 13590 -27893
rect 13650 -27943 13660 -27883
rect 13260 -27953 13660 -27943
rect 13716 -27533 14116 -27523
rect 13716 -27593 13726 -27533
rect 13786 -27583 14046 -27533
rect 13786 -27593 13796 -27583
rect 13716 -27603 13796 -27593
rect 14036 -27593 14046 -27583
rect 14106 -27593 14116 -27533
rect 14036 -27603 14116 -27593
rect 13716 -27873 13776 -27603
rect 13856 -27663 13886 -27643
rect 13836 -27703 13886 -27663
rect 13946 -27663 13976 -27643
rect 13946 -27703 13996 -27663
rect 13836 -27773 13996 -27703
rect 13836 -27813 13886 -27773
rect 13856 -27833 13886 -27813
rect 13946 -27813 13996 -27773
rect 13946 -27833 13976 -27813
rect 14056 -27863 14116 -27603
rect 14046 -27873 14116 -27863
rect 13716 -27883 13796 -27873
rect 13716 -27943 13726 -27883
rect 13786 -27893 13796 -27883
rect 14036 -27883 14116 -27873
rect 14036 -27893 14046 -27883
rect 13786 -27943 14046 -27893
rect 14106 -27943 14116 -27883
rect 13716 -27953 14116 -27943
rect 14172 -27533 14572 -27523
rect 14172 -27593 14182 -27533
rect 14242 -27583 14502 -27533
rect 14242 -27593 14252 -27583
rect 14172 -27603 14252 -27593
rect 14492 -27593 14502 -27583
rect 14562 -27593 14572 -27533
rect 14492 -27603 14572 -27593
rect 14172 -27873 14232 -27603
rect 14312 -27663 14342 -27643
rect 14292 -27703 14342 -27663
rect 14402 -27663 14432 -27643
rect 14402 -27703 14452 -27663
rect 14292 -27773 14452 -27703
rect 14292 -27813 14342 -27773
rect 14312 -27833 14342 -27813
rect 14402 -27813 14452 -27773
rect 14402 -27833 14432 -27813
rect 14512 -27863 14572 -27603
rect 14502 -27873 14572 -27863
rect 14172 -27883 14252 -27873
rect 14172 -27943 14182 -27883
rect 14242 -27893 14252 -27883
rect 14492 -27883 14572 -27873
rect 14492 -27893 14502 -27883
rect 14242 -27943 14502 -27893
rect 14562 -27943 14572 -27883
rect 14172 -27953 14572 -27943
rect 14630 -27533 15030 -27523
rect 14630 -27593 14640 -27533
rect 14700 -27583 14960 -27533
rect 14700 -27593 14710 -27583
rect 14630 -27603 14710 -27593
rect 14950 -27593 14960 -27583
rect 15020 -27593 15030 -27533
rect 14950 -27603 15030 -27593
rect 14630 -27873 14690 -27603
rect 14770 -27663 14800 -27643
rect 14750 -27703 14800 -27663
rect 14860 -27663 14890 -27643
rect 14860 -27703 14910 -27663
rect 14750 -27773 14910 -27703
rect 14750 -27813 14800 -27773
rect 14770 -27833 14800 -27813
rect 14860 -27813 14910 -27773
rect 14860 -27833 14890 -27813
rect 14970 -27863 15030 -27603
rect 14960 -27873 15030 -27863
rect 14630 -27883 14710 -27873
rect 14630 -27943 14640 -27883
rect 14700 -27893 14710 -27883
rect 14950 -27883 15030 -27873
rect 14950 -27893 14960 -27883
rect 14700 -27943 14960 -27893
rect 15020 -27943 15030 -27883
rect 14630 -27953 15030 -27943
rect 15086 -27533 15486 -27523
rect 15086 -27593 15096 -27533
rect 15156 -27583 15416 -27533
rect 15156 -27593 15166 -27583
rect 15086 -27603 15166 -27593
rect 15406 -27593 15416 -27583
rect 15476 -27593 15486 -27533
rect 15406 -27603 15486 -27593
rect 15086 -27873 15146 -27603
rect 15226 -27663 15256 -27643
rect 15206 -27703 15256 -27663
rect 15316 -27663 15346 -27643
rect 15316 -27703 15366 -27663
rect 15206 -27773 15366 -27703
rect 15206 -27813 15256 -27773
rect 15226 -27833 15256 -27813
rect 15316 -27813 15366 -27773
rect 15316 -27833 15346 -27813
rect 15426 -27863 15486 -27603
rect 15416 -27873 15486 -27863
rect 15086 -27883 15166 -27873
rect 15086 -27943 15096 -27883
rect 15156 -27893 15166 -27883
rect 15406 -27883 15486 -27873
rect 15406 -27893 15416 -27883
rect 15156 -27943 15416 -27893
rect 15476 -27943 15486 -27883
rect 15086 -27953 15486 -27943
rect 0 -28025 400 -28015
rect 0 -28085 10 -28025
rect 70 -28075 330 -28025
rect 70 -28085 80 -28075
rect 0 -28095 80 -28085
rect 320 -28085 330 -28075
rect 390 -28085 400 -28025
rect 320 -28095 400 -28085
rect 0 -28365 60 -28095
rect 140 -28155 170 -28135
rect 120 -28195 170 -28155
rect 230 -28155 260 -28135
rect 230 -28195 280 -28155
rect 120 -28265 280 -28195
rect 120 -28305 170 -28265
rect 140 -28325 170 -28305
rect 230 -28305 280 -28265
rect 230 -28325 260 -28305
rect 340 -28355 400 -28095
rect 330 -28365 400 -28355
rect 0 -28375 80 -28365
rect 0 -28435 10 -28375
rect 70 -28385 80 -28375
rect 320 -28375 400 -28365
rect 320 -28385 330 -28375
rect 70 -28435 330 -28385
rect 390 -28435 400 -28375
rect 0 -28445 400 -28435
rect 456 -28025 856 -28015
rect 456 -28085 466 -28025
rect 526 -28075 786 -28025
rect 526 -28085 536 -28075
rect 456 -28095 536 -28085
rect 776 -28085 786 -28075
rect 846 -28085 856 -28025
rect 776 -28095 856 -28085
rect 456 -28365 516 -28095
rect 596 -28155 626 -28135
rect 576 -28195 626 -28155
rect 686 -28155 716 -28135
rect 686 -28195 736 -28155
rect 576 -28265 736 -28195
rect 576 -28305 626 -28265
rect 596 -28325 626 -28305
rect 686 -28305 736 -28265
rect 686 -28325 716 -28305
rect 796 -28355 856 -28095
rect 786 -28365 856 -28355
rect 456 -28375 536 -28365
rect 456 -28435 466 -28375
rect 526 -28385 536 -28375
rect 776 -28375 856 -28365
rect 776 -28385 786 -28375
rect 526 -28435 786 -28385
rect 846 -28435 856 -28375
rect 456 -28445 856 -28435
rect 912 -28025 1312 -28015
rect 912 -28085 922 -28025
rect 982 -28075 1242 -28025
rect 982 -28085 992 -28075
rect 912 -28095 992 -28085
rect 1232 -28085 1242 -28075
rect 1302 -28085 1312 -28025
rect 1232 -28095 1312 -28085
rect 912 -28365 972 -28095
rect 1052 -28155 1082 -28135
rect 1032 -28195 1082 -28155
rect 1142 -28155 1172 -28135
rect 1142 -28195 1192 -28155
rect 1032 -28265 1192 -28195
rect 1032 -28305 1082 -28265
rect 1052 -28325 1082 -28305
rect 1142 -28305 1192 -28265
rect 1142 -28325 1172 -28305
rect 1252 -28355 1312 -28095
rect 1242 -28365 1312 -28355
rect 912 -28375 992 -28365
rect 912 -28435 922 -28375
rect 982 -28385 992 -28375
rect 1232 -28375 1312 -28365
rect 1232 -28385 1242 -28375
rect 982 -28435 1242 -28385
rect 1302 -28435 1312 -28375
rect 912 -28445 1312 -28435
rect 1370 -28025 1770 -28015
rect 1370 -28085 1380 -28025
rect 1440 -28075 1700 -28025
rect 1440 -28085 1450 -28075
rect 1370 -28095 1450 -28085
rect 1690 -28085 1700 -28075
rect 1760 -28085 1770 -28025
rect 1690 -28095 1770 -28085
rect 1370 -28365 1430 -28095
rect 1510 -28155 1540 -28135
rect 1490 -28195 1540 -28155
rect 1600 -28155 1630 -28135
rect 1600 -28195 1650 -28155
rect 1490 -28265 1650 -28195
rect 1490 -28305 1540 -28265
rect 1510 -28325 1540 -28305
rect 1600 -28305 1650 -28265
rect 1600 -28325 1630 -28305
rect 1710 -28355 1770 -28095
rect 1700 -28365 1770 -28355
rect 1370 -28375 1450 -28365
rect 1370 -28435 1380 -28375
rect 1440 -28385 1450 -28375
rect 1690 -28375 1770 -28365
rect 1690 -28385 1700 -28375
rect 1440 -28435 1700 -28385
rect 1760 -28435 1770 -28375
rect 1370 -28445 1770 -28435
rect 1826 -28025 2226 -28015
rect 1826 -28085 1836 -28025
rect 1896 -28075 2156 -28025
rect 1896 -28085 1906 -28075
rect 1826 -28095 1906 -28085
rect 2146 -28085 2156 -28075
rect 2216 -28085 2226 -28025
rect 2146 -28095 2226 -28085
rect 1826 -28365 1886 -28095
rect 1966 -28155 1996 -28135
rect 1946 -28195 1996 -28155
rect 2056 -28155 2086 -28135
rect 2056 -28195 2106 -28155
rect 1946 -28265 2106 -28195
rect 1946 -28305 1996 -28265
rect 1966 -28325 1996 -28305
rect 2056 -28305 2106 -28265
rect 2056 -28325 2086 -28305
rect 2166 -28355 2226 -28095
rect 2156 -28365 2226 -28355
rect 1826 -28375 1906 -28365
rect 1826 -28435 1836 -28375
rect 1896 -28385 1906 -28375
rect 2146 -28375 2226 -28365
rect 2146 -28385 2156 -28375
rect 1896 -28435 2156 -28385
rect 2216 -28435 2226 -28375
rect 1826 -28445 2226 -28435
rect 2282 -28025 2682 -28015
rect 2282 -28085 2292 -28025
rect 2352 -28075 2612 -28025
rect 2352 -28085 2362 -28075
rect 2282 -28095 2362 -28085
rect 2602 -28085 2612 -28075
rect 2672 -28085 2682 -28025
rect 2602 -28095 2682 -28085
rect 2282 -28365 2342 -28095
rect 2422 -28155 2452 -28135
rect 2402 -28195 2452 -28155
rect 2512 -28155 2542 -28135
rect 2512 -28195 2562 -28155
rect 2402 -28265 2562 -28195
rect 2402 -28305 2452 -28265
rect 2422 -28325 2452 -28305
rect 2512 -28305 2562 -28265
rect 2512 -28325 2542 -28305
rect 2622 -28355 2682 -28095
rect 2612 -28365 2682 -28355
rect 2282 -28375 2362 -28365
rect 2282 -28435 2292 -28375
rect 2352 -28385 2362 -28375
rect 2602 -28375 2682 -28365
rect 2602 -28385 2612 -28375
rect 2352 -28435 2612 -28385
rect 2672 -28435 2682 -28375
rect 2282 -28445 2682 -28435
rect 2740 -28025 3140 -28015
rect 2740 -28085 2750 -28025
rect 2810 -28075 3070 -28025
rect 2810 -28085 2820 -28075
rect 2740 -28095 2820 -28085
rect 3060 -28085 3070 -28075
rect 3130 -28085 3140 -28025
rect 3060 -28095 3140 -28085
rect 2740 -28365 2800 -28095
rect 2880 -28155 2910 -28135
rect 2860 -28195 2910 -28155
rect 2970 -28155 3000 -28135
rect 2970 -28195 3020 -28155
rect 2860 -28265 3020 -28195
rect 2860 -28305 2910 -28265
rect 2880 -28325 2910 -28305
rect 2970 -28305 3020 -28265
rect 2970 -28325 3000 -28305
rect 3080 -28355 3140 -28095
rect 3070 -28365 3140 -28355
rect 2740 -28375 2820 -28365
rect 2740 -28435 2750 -28375
rect 2810 -28385 2820 -28375
rect 3060 -28375 3140 -28365
rect 3060 -28385 3070 -28375
rect 2810 -28435 3070 -28385
rect 3130 -28435 3140 -28375
rect 2740 -28445 3140 -28435
rect 3196 -28025 3596 -28015
rect 3196 -28085 3206 -28025
rect 3266 -28075 3526 -28025
rect 3266 -28085 3276 -28075
rect 3196 -28095 3276 -28085
rect 3516 -28085 3526 -28075
rect 3586 -28085 3596 -28025
rect 3516 -28095 3596 -28085
rect 3196 -28365 3256 -28095
rect 3336 -28155 3366 -28135
rect 3316 -28195 3366 -28155
rect 3426 -28155 3456 -28135
rect 3426 -28195 3476 -28155
rect 3316 -28265 3476 -28195
rect 3316 -28305 3366 -28265
rect 3336 -28325 3366 -28305
rect 3426 -28305 3476 -28265
rect 3426 -28325 3456 -28305
rect 3536 -28355 3596 -28095
rect 3526 -28365 3596 -28355
rect 3196 -28375 3276 -28365
rect 3196 -28435 3206 -28375
rect 3266 -28385 3276 -28375
rect 3516 -28375 3596 -28365
rect 3516 -28385 3526 -28375
rect 3266 -28435 3526 -28385
rect 3586 -28435 3596 -28375
rect 3196 -28445 3596 -28435
rect 3652 -28025 4052 -28015
rect 3652 -28085 3662 -28025
rect 3722 -28075 3982 -28025
rect 3722 -28085 3732 -28075
rect 3652 -28095 3732 -28085
rect 3972 -28085 3982 -28075
rect 4042 -28085 4052 -28025
rect 3972 -28095 4052 -28085
rect 3652 -28365 3712 -28095
rect 3792 -28155 3822 -28135
rect 3772 -28195 3822 -28155
rect 3882 -28155 3912 -28135
rect 3882 -28195 3932 -28155
rect 3772 -28265 3932 -28195
rect 3772 -28305 3822 -28265
rect 3792 -28325 3822 -28305
rect 3882 -28305 3932 -28265
rect 3882 -28325 3912 -28305
rect 3992 -28355 4052 -28095
rect 3982 -28365 4052 -28355
rect 3652 -28375 3732 -28365
rect 3652 -28435 3662 -28375
rect 3722 -28385 3732 -28375
rect 3972 -28375 4052 -28365
rect 3972 -28385 3982 -28375
rect 3722 -28435 3982 -28385
rect 4042 -28435 4052 -28375
rect 3652 -28445 4052 -28435
rect 4110 -28025 4510 -28015
rect 4110 -28085 4120 -28025
rect 4180 -28075 4440 -28025
rect 4180 -28085 4190 -28075
rect 4110 -28095 4190 -28085
rect 4430 -28085 4440 -28075
rect 4500 -28085 4510 -28025
rect 4430 -28095 4510 -28085
rect 4110 -28365 4170 -28095
rect 4250 -28155 4280 -28135
rect 4230 -28195 4280 -28155
rect 4340 -28155 4370 -28135
rect 4340 -28195 4390 -28155
rect 4230 -28265 4390 -28195
rect 4230 -28305 4280 -28265
rect 4250 -28325 4280 -28305
rect 4340 -28305 4390 -28265
rect 4340 -28325 4370 -28305
rect 4450 -28355 4510 -28095
rect 4440 -28365 4510 -28355
rect 4110 -28375 4190 -28365
rect 4110 -28435 4120 -28375
rect 4180 -28385 4190 -28375
rect 4430 -28375 4510 -28365
rect 4430 -28385 4440 -28375
rect 4180 -28435 4440 -28385
rect 4500 -28435 4510 -28375
rect 4110 -28445 4510 -28435
rect 4566 -28025 4966 -28015
rect 4566 -28085 4576 -28025
rect 4636 -28075 4896 -28025
rect 4636 -28085 4646 -28075
rect 4566 -28095 4646 -28085
rect 4886 -28085 4896 -28075
rect 4956 -28085 4966 -28025
rect 4886 -28095 4966 -28085
rect 4566 -28365 4626 -28095
rect 4706 -28155 4736 -28135
rect 4686 -28195 4736 -28155
rect 4796 -28155 4826 -28135
rect 4796 -28195 4846 -28155
rect 4686 -28265 4846 -28195
rect 4686 -28305 4736 -28265
rect 4706 -28325 4736 -28305
rect 4796 -28305 4846 -28265
rect 4796 -28325 4826 -28305
rect 4906 -28355 4966 -28095
rect 4896 -28365 4966 -28355
rect 4566 -28375 4646 -28365
rect 4566 -28435 4576 -28375
rect 4636 -28385 4646 -28375
rect 4886 -28375 4966 -28365
rect 4886 -28385 4896 -28375
rect 4636 -28435 4896 -28385
rect 4956 -28435 4966 -28375
rect 4566 -28445 4966 -28435
rect 5022 -28025 5422 -28015
rect 5022 -28085 5032 -28025
rect 5092 -28075 5352 -28025
rect 5092 -28085 5102 -28075
rect 5022 -28095 5102 -28085
rect 5342 -28085 5352 -28075
rect 5412 -28085 5422 -28025
rect 5342 -28095 5422 -28085
rect 5022 -28365 5082 -28095
rect 5162 -28155 5192 -28135
rect 5142 -28195 5192 -28155
rect 5252 -28155 5282 -28135
rect 5252 -28195 5302 -28155
rect 5142 -28265 5302 -28195
rect 5142 -28305 5192 -28265
rect 5162 -28325 5192 -28305
rect 5252 -28305 5302 -28265
rect 5252 -28325 5282 -28305
rect 5362 -28355 5422 -28095
rect 5352 -28365 5422 -28355
rect 5022 -28375 5102 -28365
rect 5022 -28435 5032 -28375
rect 5092 -28385 5102 -28375
rect 5342 -28375 5422 -28365
rect 5342 -28385 5352 -28375
rect 5092 -28435 5352 -28385
rect 5412 -28435 5422 -28375
rect 5022 -28445 5422 -28435
rect 5480 -28025 5880 -28015
rect 5480 -28085 5490 -28025
rect 5550 -28075 5810 -28025
rect 5550 -28085 5560 -28075
rect 5480 -28095 5560 -28085
rect 5800 -28085 5810 -28075
rect 5870 -28085 5880 -28025
rect 5800 -28095 5880 -28085
rect 5480 -28365 5540 -28095
rect 5620 -28155 5650 -28135
rect 5600 -28195 5650 -28155
rect 5710 -28155 5740 -28135
rect 5710 -28195 5760 -28155
rect 5600 -28265 5760 -28195
rect 5600 -28305 5650 -28265
rect 5620 -28325 5650 -28305
rect 5710 -28305 5760 -28265
rect 5710 -28325 5740 -28305
rect 5820 -28355 5880 -28095
rect 5810 -28365 5880 -28355
rect 5480 -28375 5560 -28365
rect 5480 -28435 5490 -28375
rect 5550 -28385 5560 -28375
rect 5800 -28375 5880 -28365
rect 5800 -28385 5810 -28375
rect 5550 -28435 5810 -28385
rect 5870 -28435 5880 -28375
rect 5480 -28445 5880 -28435
rect 5936 -28025 6336 -28015
rect 5936 -28085 5946 -28025
rect 6006 -28075 6266 -28025
rect 6006 -28085 6016 -28075
rect 5936 -28095 6016 -28085
rect 6256 -28085 6266 -28075
rect 6326 -28085 6336 -28025
rect 6256 -28095 6336 -28085
rect 5936 -28365 5996 -28095
rect 6076 -28155 6106 -28135
rect 6056 -28195 6106 -28155
rect 6166 -28155 6196 -28135
rect 6166 -28195 6216 -28155
rect 6056 -28265 6216 -28195
rect 6056 -28305 6106 -28265
rect 6076 -28325 6106 -28305
rect 6166 -28305 6216 -28265
rect 6166 -28325 6196 -28305
rect 6276 -28355 6336 -28095
rect 6266 -28365 6336 -28355
rect 5936 -28375 6016 -28365
rect 5936 -28435 5946 -28375
rect 6006 -28385 6016 -28375
rect 6256 -28375 6336 -28365
rect 6256 -28385 6266 -28375
rect 6006 -28435 6266 -28385
rect 6326 -28435 6336 -28375
rect 5936 -28445 6336 -28435
rect 6392 -28025 6792 -28015
rect 6392 -28085 6402 -28025
rect 6462 -28075 6722 -28025
rect 6462 -28085 6472 -28075
rect 6392 -28095 6472 -28085
rect 6712 -28085 6722 -28075
rect 6782 -28085 6792 -28025
rect 6712 -28095 6792 -28085
rect 6392 -28365 6452 -28095
rect 6532 -28155 6562 -28135
rect 6512 -28195 6562 -28155
rect 6622 -28155 6652 -28135
rect 6622 -28195 6672 -28155
rect 6512 -28265 6672 -28195
rect 6512 -28305 6562 -28265
rect 6532 -28325 6562 -28305
rect 6622 -28305 6672 -28265
rect 6622 -28325 6652 -28305
rect 6732 -28355 6792 -28095
rect 6722 -28365 6792 -28355
rect 6392 -28375 6472 -28365
rect 6392 -28435 6402 -28375
rect 6462 -28385 6472 -28375
rect 6712 -28375 6792 -28365
rect 6712 -28385 6722 -28375
rect 6462 -28435 6722 -28385
rect 6782 -28435 6792 -28375
rect 6392 -28445 6792 -28435
rect 6850 -28025 7250 -28015
rect 6850 -28085 6860 -28025
rect 6920 -28075 7180 -28025
rect 6920 -28085 6930 -28075
rect 6850 -28095 6930 -28085
rect 7170 -28085 7180 -28075
rect 7240 -28085 7250 -28025
rect 7170 -28095 7250 -28085
rect 6850 -28365 6910 -28095
rect 6990 -28155 7020 -28135
rect 6970 -28195 7020 -28155
rect 7080 -28155 7110 -28135
rect 7080 -28195 7130 -28155
rect 6970 -28265 7130 -28195
rect 6970 -28305 7020 -28265
rect 6990 -28325 7020 -28305
rect 7080 -28305 7130 -28265
rect 7080 -28325 7110 -28305
rect 7190 -28355 7250 -28095
rect 7180 -28365 7250 -28355
rect 6850 -28375 6930 -28365
rect 6850 -28435 6860 -28375
rect 6920 -28385 6930 -28375
rect 7170 -28375 7250 -28365
rect 7170 -28385 7180 -28375
rect 6920 -28435 7180 -28385
rect 7240 -28435 7250 -28375
rect 6850 -28445 7250 -28435
rect 7306 -28025 7706 -28015
rect 7306 -28085 7316 -28025
rect 7376 -28075 7636 -28025
rect 7376 -28085 7386 -28075
rect 7306 -28095 7386 -28085
rect 7626 -28085 7636 -28075
rect 7696 -28085 7706 -28025
rect 7626 -28095 7706 -28085
rect 7306 -28365 7366 -28095
rect 7446 -28155 7476 -28135
rect 7426 -28195 7476 -28155
rect 7536 -28155 7566 -28135
rect 7536 -28195 7586 -28155
rect 7426 -28265 7586 -28195
rect 7426 -28305 7476 -28265
rect 7446 -28325 7476 -28305
rect 7536 -28305 7586 -28265
rect 7536 -28325 7566 -28305
rect 7646 -28355 7706 -28095
rect 7636 -28365 7706 -28355
rect 7306 -28375 7386 -28365
rect 7306 -28435 7316 -28375
rect 7376 -28385 7386 -28375
rect 7626 -28375 7706 -28365
rect 7626 -28385 7636 -28375
rect 7376 -28435 7636 -28385
rect 7696 -28435 7706 -28375
rect 7306 -28445 7706 -28435
rect 7762 -28025 8162 -28015
rect 7762 -28085 7772 -28025
rect 7832 -28075 8092 -28025
rect 7832 -28085 7842 -28075
rect 7762 -28095 7842 -28085
rect 8082 -28085 8092 -28075
rect 8152 -28085 8162 -28025
rect 8082 -28095 8162 -28085
rect 7762 -28365 7822 -28095
rect 7902 -28155 7932 -28135
rect 7882 -28195 7932 -28155
rect 7992 -28155 8022 -28135
rect 7992 -28195 8042 -28155
rect 7882 -28265 8042 -28195
rect 7882 -28305 7932 -28265
rect 7902 -28325 7932 -28305
rect 7992 -28305 8042 -28265
rect 7992 -28325 8022 -28305
rect 8102 -28355 8162 -28095
rect 8092 -28365 8162 -28355
rect 7762 -28375 7842 -28365
rect 7762 -28435 7772 -28375
rect 7832 -28385 7842 -28375
rect 8082 -28375 8162 -28365
rect 8082 -28385 8092 -28375
rect 7832 -28435 8092 -28385
rect 8152 -28435 8162 -28375
rect 7762 -28445 8162 -28435
rect 8236 -28025 8636 -28015
rect 8236 -28085 8246 -28025
rect 8306 -28075 8566 -28025
rect 8306 -28085 8316 -28075
rect 8236 -28095 8316 -28085
rect 8556 -28085 8566 -28075
rect 8626 -28085 8636 -28025
rect 8556 -28095 8636 -28085
rect 8236 -28365 8296 -28095
rect 8376 -28155 8406 -28135
rect 8356 -28195 8406 -28155
rect 8466 -28155 8496 -28135
rect 8466 -28195 8516 -28155
rect 8356 -28265 8516 -28195
rect 8356 -28305 8406 -28265
rect 8376 -28325 8406 -28305
rect 8466 -28305 8516 -28265
rect 8466 -28325 8496 -28305
rect 8576 -28355 8636 -28095
rect 8566 -28365 8636 -28355
rect 8236 -28375 8316 -28365
rect 8236 -28435 8246 -28375
rect 8306 -28385 8316 -28375
rect 8556 -28375 8636 -28365
rect 8556 -28385 8566 -28375
rect 8306 -28435 8566 -28385
rect 8626 -28435 8636 -28375
rect 8236 -28445 8636 -28435
rect 8692 -28025 9092 -28015
rect 8692 -28085 8702 -28025
rect 8762 -28075 9022 -28025
rect 8762 -28085 8772 -28075
rect 8692 -28095 8772 -28085
rect 9012 -28085 9022 -28075
rect 9082 -28085 9092 -28025
rect 9012 -28095 9092 -28085
rect 8692 -28365 8752 -28095
rect 8832 -28155 8862 -28135
rect 8812 -28195 8862 -28155
rect 8922 -28155 8952 -28135
rect 8922 -28195 8972 -28155
rect 8812 -28265 8972 -28195
rect 8812 -28305 8862 -28265
rect 8832 -28325 8862 -28305
rect 8922 -28305 8972 -28265
rect 8922 -28325 8952 -28305
rect 9032 -28355 9092 -28095
rect 9022 -28365 9092 -28355
rect 8692 -28375 8772 -28365
rect 8692 -28435 8702 -28375
rect 8762 -28385 8772 -28375
rect 9012 -28375 9092 -28365
rect 9012 -28385 9022 -28375
rect 8762 -28435 9022 -28385
rect 9082 -28435 9092 -28375
rect 8692 -28445 9092 -28435
rect 9150 -28025 9550 -28015
rect 9150 -28085 9160 -28025
rect 9220 -28075 9480 -28025
rect 9220 -28085 9230 -28075
rect 9150 -28095 9230 -28085
rect 9470 -28085 9480 -28075
rect 9540 -28085 9550 -28025
rect 9470 -28095 9550 -28085
rect 9150 -28365 9210 -28095
rect 9290 -28155 9320 -28135
rect 9270 -28195 9320 -28155
rect 9380 -28155 9410 -28135
rect 9380 -28195 9430 -28155
rect 9270 -28265 9430 -28195
rect 9270 -28305 9320 -28265
rect 9290 -28325 9320 -28305
rect 9380 -28305 9430 -28265
rect 9380 -28325 9410 -28305
rect 9490 -28355 9550 -28095
rect 9480 -28365 9550 -28355
rect 9150 -28375 9230 -28365
rect 9150 -28435 9160 -28375
rect 9220 -28385 9230 -28375
rect 9470 -28375 9550 -28365
rect 9470 -28385 9480 -28375
rect 9220 -28435 9480 -28385
rect 9540 -28435 9550 -28375
rect 9150 -28445 9550 -28435
rect 9606 -28025 10006 -28015
rect 9606 -28085 9616 -28025
rect 9676 -28075 9936 -28025
rect 9676 -28085 9686 -28075
rect 9606 -28095 9686 -28085
rect 9926 -28085 9936 -28075
rect 9996 -28085 10006 -28025
rect 9926 -28095 10006 -28085
rect 9606 -28365 9666 -28095
rect 9746 -28155 9776 -28135
rect 9726 -28195 9776 -28155
rect 9836 -28155 9866 -28135
rect 9836 -28195 9886 -28155
rect 9726 -28265 9886 -28195
rect 9726 -28305 9776 -28265
rect 9746 -28325 9776 -28305
rect 9836 -28305 9886 -28265
rect 9836 -28325 9866 -28305
rect 9946 -28355 10006 -28095
rect 9936 -28365 10006 -28355
rect 9606 -28375 9686 -28365
rect 9606 -28435 9616 -28375
rect 9676 -28385 9686 -28375
rect 9926 -28375 10006 -28365
rect 9926 -28385 9936 -28375
rect 9676 -28435 9936 -28385
rect 9996 -28435 10006 -28375
rect 9606 -28445 10006 -28435
rect 10062 -28025 10462 -28015
rect 10062 -28085 10072 -28025
rect 10132 -28075 10392 -28025
rect 10132 -28085 10142 -28075
rect 10062 -28095 10142 -28085
rect 10382 -28085 10392 -28075
rect 10452 -28085 10462 -28025
rect 10382 -28095 10462 -28085
rect 10062 -28365 10122 -28095
rect 10202 -28155 10232 -28135
rect 10182 -28195 10232 -28155
rect 10292 -28155 10322 -28135
rect 10292 -28195 10342 -28155
rect 10182 -28265 10342 -28195
rect 10182 -28305 10232 -28265
rect 10202 -28325 10232 -28305
rect 10292 -28305 10342 -28265
rect 10292 -28325 10322 -28305
rect 10402 -28355 10462 -28095
rect 10392 -28365 10462 -28355
rect 10062 -28375 10142 -28365
rect 10062 -28435 10072 -28375
rect 10132 -28385 10142 -28375
rect 10382 -28375 10462 -28365
rect 10382 -28385 10392 -28375
rect 10132 -28435 10392 -28385
rect 10452 -28435 10462 -28375
rect 10062 -28445 10462 -28435
rect 10520 -28025 10920 -28015
rect 10520 -28085 10530 -28025
rect 10590 -28075 10850 -28025
rect 10590 -28085 10600 -28075
rect 10520 -28095 10600 -28085
rect 10840 -28085 10850 -28075
rect 10910 -28085 10920 -28025
rect 10840 -28095 10920 -28085
rect 10520 -28365 10580 -28095
rect 10660 -28155 10690 -28135
rect 10640 -28195 10690 -28155
rect 10750 -28155 10780 -28135
rect 10750 -28195 10800 -28155
rect 10640 -28265 10800 -28195
rect 10640 -28305 10690 -28265
rect 10660 -28325 10690 -28305
rect 10750 -28305 10800 -28265
rect 10750 -28325 10780 -28305
rect 10860 -28355 10920 -28095
rect 10850 -28365 10920 -28355
rect 10520 -28375 10600 -28365
rect 10520 -28435 10530 -28375
rect 10590 -28385 10600 -28375
rect 10840 -28375 10920 -28365
rect 10840 -28385 10850 -28375
rect 10590 -28435 10850 -28385
rect 10910 -28435 10920 -28375
rect 10520 -28445 10920 -28435
rect 10976 -28025 11376 -28015
rect 10976 -28085 10986 -28025
rect 11046 -28075 11306 -28025
rect 11046 -28085 11056 -28075
rect 10976 -28095 11056 -28085
rect 11296 -28085 11306 -28075
rect 11366 -28085 11376 -28025
rect 11296 -28095 11376 -28085
rect 10976 -28365 11036 -28095
rect 11116 -28155 11146 -28135
rect 11096 -28195 11146 -28155
rect 11206 -28155 11236 -28135
rect 11206 -28195 11256 -28155
rect 11096 -28265 11256 -28195
rect 11096 -28305 11146 -28265
rect 11116 -28325 11146 -28305
rect 11206 -28305 11256 -28265
rect 11206 -28325 11236 -28305
rect 11316 -28355 11376 -28095
rect 11306 -28365 11376 -28355
rect 10976 -28375 11056 -28365
rect 10976 -28435 10986 -28375
rect 11046 -28385 11056 -28375
rect 11296 -28375 11376 -28365
rect 11296 -28385 11306 -28375
rect 11046 -28435 11306 -28385
rect 11366 -28435 11376 -28375
rect 10976 -28445 11376 -28435
rect 11432 -28025 11832 -28015
rect 11432 -28085 11442 -28025
rect 11502 -28075 11762 -28025
rect 11502 -28085 11512 -28075
rect 11432 -28095 11512 -28085
rect 11752 -28085 11762 -28075
rect 11822 -28085 11832 -28025
rect 11752 -28095 11832 -28085
rect 11432 -28365 11492 -28095
rect 11572 -28155 11602 -28135
rect 11552 -28195 11602 -28155
rect 11662 -28155 11692 -28135
rect 11662 -28195 11712 -28155
rect 11552 -28265 11712 -28195
rect 11552 -28305 11602 -28265
rect 11572 -28325 11602 -28305
rect 11662 -28305 11712 -28265
rect 11662 -28325 11692 -28305
rect 11772 -28355 11832 -28095
rect 11762 -28365 11832 -28355
rect 11432 -28375 11512 -28365
rect 11432 -28435 11442 -28375
rect 11502 -28385 11512 -28375
rect 11752 -28375 11832 -28365
rect 11752 -28385 11762 -28375
rect 11502 -28435 11762 -28385
rect 11822 -28435 11832 -28375
rect 11432 -28445 11832 -28435
rect 11890 -28025 12290 -28015
rect 11890 -28085 11900 -28025
rect 11960 -28075 12220 -28025
rect 11960 -28085 11970 -28075
rect 11890 -28095 11970 -28085
rect 12210 -28085 12220 -28075
rect 12280 -28085 12290 -28025
rect 12210 -28095 12290 -28085
rect 11890 -28365 11950 -28095
rect 12030 -28155 12060 -28135
rect 12010 -28195 12060 -28155
rect 12120 -28155 12150 -28135
rect 12120 -28195 12170 -28155
rect 12010 -28265 12170 -28195
rect 12010 -28305 12060 -28265
rect 12030 -28325 12060 -28305
rect 12120 -28305 12170 -28265
rect 12120 -28325 12150 -28305
rect 12230 -28355 12290 -28095
rect 12220 -28365 12290 -28355
rect 11890 -28375 11970 -28365
rect 11890 -28435 11900 -28375
rect 11960 -28385 11970 -28375
rect 12210 -28375 12290 -28365
rect 12210 -28385 12220 -28375
rect 11960 -28435 12220 -28385
rect 12280 -28435 12290 -28375
rect 11890 -28445 12290 -28435
rect 12346 -28025 12746 -28015
rect 12346 -28085 12356 -28025
rect 12416 -28075 12676 -28025
rect 12416 -28085 12426 -28075
rect 12346 -28095 12426 -28085
rect 12666 -28085 12676 -28075
rect 12736 -28085 12746 -28025
rect 12666 -28095 12746 -28085
rect 12346 -28365 12406 -28095
rect 12486 -28155 12516 -28135
rect 12466 -28195 12516 -28155
rect 12576 -28155 12606 -28135
rect 12576 -28195 12626 -28155
rect 12466 -28265 12626 -28195
rect 12466 -28305 12516 -28265
rect 12486 -28325 12516 -28305
rect 12576 -28305 12626 -28265
rect 12576 -28325 12606 -28305
rect 12686 -28355 12746 -28095
rect 12676 -28365 12746 -28355
rect 12346 -28375 12426 -28365
rect 12346 -28435 12356 -28375
rect 12416 -28385 12426 -28375
rect 12666 -28375 12746 -28365
rect 12666 -28385 12676 -28375
rect 12416 -28435 12676 -28385
rect 12736 -28435 12746 -28375
rect 12346 -28445 12746 -28435
rect 12802 -28025 13202 -28015
rect 12802 -28085 12812 -28025
rect 12872 -28075 13132 -28025
rect 12872 -28085 12882 -28075
rect 12802 -28095 12882 -28085
rect 13122 -28085 13132 -28075
rect 13192 -28085 13202 -28025
rect 13122 -28095 13202 -28085
rect 12802 -28365 12862 -28095
rect 12942 -28155 12972 -28135
rect 12922 -28195 12972 -28155
rect 13032 -28155 13062 -28135
rect 13032 -28195 13082 -28155
rect 12922 -28265 13082 -28195
rect 12922 -28305 12972 -28265
rect 12942 -28325 12972 -28305
rect 13032 -28305 13082 -28265
rect 13032 -28325 13062 -28305
rect 13142 -28355 13202 -28095
rect 13132 -28365 13202 -28355
rect 12802 -28375 12882 -28365
rect 12802 -28435 12812 -28375
rect 12872 -28385 12882 -28375
rect 13122 -28375 13202 -28365
rect 13122 -28385 13132 -28375
rect 12872 -28435 13132 -28385
rect 13192 -28435 13202 -28375
rect 12802 -28445 13202 -28435
rect 13260 -28025 13660 -28015
rect 13260 -28085 13270 -28025
rect 13330 -28075 13590 -28025
rect 13330 -28085 13340 -28075
rect 13260 -28095 13340 -28085
rect 13580 -28085 13590 -28075
rect 13650 -28085 13660 -28025
rect 13580 -28095 13660 -28085
rect 13260 -28365 13320 -28095
rect 13400 -28155 13430 -28135
rect 13380 -28195 13430 -28155
rect 13490 -28155 13520 -28135
rect 13490 -28195 13540 -28155
rect 13380 -28265 13540 -28195
rect 13380 -28305 13430 -28265
rect 13400 -28325 13430 -28305
rect 13490 -28305 13540 -28265
rect 13490 -28325 13520 -28305
rect 13600 -28355 13660 -28095
rect 13590 -28365 13660 -28355
rect 13260 -28375 13340 -28365
rect 13260 -28435 13270 -28375
rect 13330 -28385 13340 -28375
rect 13580 -28375 13660 -28365
rect 13580 -28385 13590 -28375
rect 13330 -28435 13590 -28385
rect 13650 -28435 13660 -28375
rect 13260 -28445 13660 -28435
rect 13716 -28025 14116 -28015
rect 13716 -28085 13726 -28025
rect 13786 -28075 14046 -28025
rect 13786 -28085 13796 -28075
rect 13716 -28095 13796 -28085
rect 14036 -28085 14046 -28075
rect 14106 -28085 14116 -28025
rect 14036 -28095 14116 -28085
rect 13716 -28365 13776 -28095
rect 13856 -28155 13886 -28135
rect 13836 -28195 13886 -28155
rect 13946 -28155 13976 -28135
rect 13946 -28195 13996 -28155
rect 13836 -28265 13996 -28195
rect 13836 -28305 13886 -28265
rect 13856 -28325 13886 -28305
rect 13946 -28305 13996 -28265
rect 13946 -28325 13976 -28305
rect 14056 -28355 14116 -28095
rect 14046 -28365 14116 -28355
rect 13716 -28375 13796 -28365
rect 13716 -28435 13726 -28375
rect 13786 -28385 13796 -28375
rect 14036 -28375 14116 -28365
rect 14036 -28385 14046 -28375
rect 13786 -28435 14046 -28385
rect 14106 -28435 14116 -28375
rect 13716 -28445 14116 -28435
rect 14172 -28025 14572 -28015
rect 14172 -28085 14182 -28025
rect 14242 -28075 14502 -28025
rect 14242 -28085 14252 -28075
rect 14172 -28095 14252 -28085
rect 14492 -28085 14502 -28075
rect 14562 -28085 14572 -28025
rect 14492 -28095 14572 -28085
rect 14172 -28365 14232 -28095
rect 14312 -28155 14342 -28135
rect 14292 -28195 14342 -28155
rect 14402 -28155 14432 -28135
rect 14402 -28195 14452 -28155
rect 14292 -28265 14452 -28195
rect 14292 -28305 14342 -28265
rect 14312 -28325 14342 -28305
rect 14402 -28305 14452 -28265
rect 14402 -28325 14432 -28305
rect 14512 -28355 14572 -28095
rect 14502 -28365 14572 -28355
rect 14172 -28375 14252 -28365
rect 14172 -28435 14182 -28375
rect 14242 -28385 14252 -28375
rect 14492 -28375 14572 -28365
rect 14492 -28385 14502 -28375
rect 14242 -28435 14502 -28385
rect 14562 -28435 14572 -28375
rect 14172 -28445 14572 -28435
rect 14630 -28025 15030 -28015
rect 14630 -28085 14640 -28025
rect 14700 -28075 14960 -28025
rect 14700 -28085 14710 -28075
rect 14630 -28095 14710 -28085
rect 14950 -28085 14960 -28075
rect 15020 -28085 15030 -28025
rect 14950 -28095 15030 -28085
rect 14630 -28365 14690 -28095
rect 14770 -28155 14800 -28135
rect 14750 -28195 14800 -28155
rect 14860 -28155 14890 -28135
rect 14860 -28195 14910 -28155
rect 14750 -28265 14910 -28195
rect 14750 -28305 14800 -28265
rect 14770 -28325 14800 -28305
rect 14860 -28305 14910 -28265
rect 14860 -28325 14890 -28305
rect 14970 -28355 15030 -28095
rect 14960 -28365 15030 -28355
rect 14630 -28375 14710 -28365
rect 14630 -28435 14640 -28375
rect 14700 -28385 14710 -28375
rect 14950 -28375 15030 -28365
rect 14950 -28385 14960 -28375
rect 14700 -28435 14960 -28385
rect 15020 -28435 15030 -28375
rect 14630 -28445 15030 -28435
rect 15086 -28025 15486 -28015
rect 15086 -28085 15096 -28025
rect 15156 -28075 15416 -28025
rect 15156 -28085 15166 -28075
rect 15086 -28095 15166 -28085
rect 15406 -28085 15416 -28075
rect 15476 -28085 15486 -28025
rect 15406 -28095 15486 -28085
rect 15086 -28365 15146 -28095
rect 15226 -28155 15256 -28135
rect 15206 -28195 15256 -28155
rect 15316 -28155 15346 -28135
rect 15316 -28195 15366 -28155
rect 15206 -28265 15366 -28195
rect 15206 -28305 15256 -28265
rect 15226 -28325 15256 -28305
rect 15316 -28305 15366 -28265
rect 15316 -28325 15346 -28305
rect 15426 -28355 15486 -28095
rect 15416 -28365 15486 -28355
rect 15086 -28375 15166 -28365
rect 15086 -28435 15096 -28375
rect 15156 -28385 15166 -28375
rect 15406 -28375 15486 -28365
rect 15406 -28385 15416 -28375
rect 15156 -28435 15416 -28385
rect 15476 -28435 15486 -28375
rect 15086 -28445 15486 -28435
rect 0 -28527 400 -28517
rect 0 -28587 10 -28527
rect 70 -28577 330 -28527
rect 70 -28587 80 -28577
rect 0 -28597 80 -28587
rect 320 -28587 330 -28577
rect 390 -28587 400 -28527
rect 320 -28597 400 -28587
rect 0 -28867 60 -28597
rect 140 -28657 170 -28637
rect 120 -28697 170 -28657
rect 230 -28657 260 -28637
rect 230 -28697 280 -28657
rect 120 -28767 280 -28697
rect 120 -28807 170 -28767
rect 140 -28827 170 -28807
rect 230 -28807 280 -28767
rect 230 -28827 260 -28807
rect 340 -28857 400 -28597
rect 330 -28867 400 -28857
rect 0 -28877 80 -28867
rect 0 -28937 10 -28877
rect 70 -28887 80 -28877
rect 320 -28877 400 -28867
rect 320 -28887 330 -28877
rect 70 -28937 330 -28887
rect 390 -28937 400 -28877
rect 0 -28947 400 -28937
rect 456 -28527 856 -28517
rect 456 -28587 466 -28527
rect 526 -28577 786 -28527
rect 526 -28587 536 -28577
rect 456 -28597 536 -28587
rect 776 -28587 786 -28577
rect 846 -28587 856 -28527
rect 776 -28597 856 -28587
rect 456 -28867 516 -28597
rect 596 -28657 626 -28637
rect 576 -28697 626 -28657
rect 686 -28657 716 -28637
rect 686 -28697 736 -28657
rect 576 -28767 736 -28697
rect 576 -28807 626 -28767
rect 596 -28827 626 -28807
rect 686 -28807 736 -28767
rect 686 -28827 716 -28807
rect 796 -28857 856 -28597
rect 786 -28867 856 -28857
rect 456 -28877 536 -28867
rect 456 -28937 466 -28877
rect 526 -28887 536 -28877
rect 776 -28877 856 -28867
rect 776 -28887 786 -28877
rect 526 -28937 786 -28887
rect 846 -28937 856 -28877
rect 456 -28947 856 -28937
rect 912 -28527 1312 -28517
rect 912 -28587 922 -28527
rect 982 -28577 1242 -28527
rect 982 -28587 992 -28577
rect 912 -28597 992 -28587
rect 1232 -28587 1242 -28577
rect 1302 -28587 1312 -28527
rect 1232 -28597 1312 -28587
rect 912 -28867 972 -28597
rect 1052 -28657 1082 -28637
rect 1032 -28697 1082 -28657
rect 1142 -28657 1172 -28637
rect 1142 -28697 1192 -28657
rect 1032 -28767 1192 -28697
rect 1032 -28807 1082 -28767
rect 1052 -28827 1082 -28807
rect 1142 -28807 1192 -28767
rect 1142 -28827 1172 -28807
rect 1252 -28857 1312 -28597
rect 1242 -28867 1312 -28857
rect 912 -28877 992 -28867
rect 912 -28937 922 -28877
rect 982 -28887 992 -28877
rect 1232 -28877 1312 -28867
rect 1232 -28887 1242 -28877
rect 982 -28937 1242 -28887
rect 1302 -28937 1312 -28877
rect 912 -28947 1312 -28937
rect 1370 -28527 1770 -28517
rect 1370 -28587 1380 -28527
rect 1440 -28577 1700 -28527
rect 1440 -28587 1450 -28577
rect 1370 -28597 1450 -28587
rect 1690 -28587 1700 -28577
rect 1760 -28587 1770 -28527
rect 1690 -28597 1770 -28587
rect 1370 -28867 1430 -28597
rect 1510 -28657 1540 -28637
rect 1490 -28697 1540 -28657
rect 1600 -28657 1630 -28637
rect 1600 -28697 1650 -28657
rect 1490 -28767 1650 -28697
rect 1490 -28807 1540 -28767
rect 1510 -28827 1540 -28807
rect 1600 -28807 1650 -28767
rect 1600 -28827 1630 -28807
rect 1710 -28857 1770 -28597
rect 1700 -28867 1770 -28857
rect 1370 -28877 1450 -28867
rect 1370 -28937 1380 -28877
rect 1440 -28887 1450 -28877
rect 1690 -28877 1770 -28867
rect 1690 -28887 1700 -28877
rect 1440 -28937 1700 -28887
rect 1760 -28937 1770 -28877
rect 1370 -28947 1770 -28937
rect 1826 -28527 2226 -28517
rect 1826 -28587 1836 -28527
rect 1896 -28577 2156 -28527
rect 1896 -28587 1906 -28577
rect 1826 -28597 1906 -28587
rect 2146 -28587 2156 -28577
rect 2216 -28587 2226 -28527
rect 2146 -28597 2226 -28587
rect 1826 -28867 1886 -28597
rect 1966 -28657 1996 -28637
rect 1946 -28697 1996 -28657
rect 2056 -28657 2086 -28637
rect 2056 -28697 2106 -28657
rect 1946 -28767 2106 -28697
rect 1946 -28807 1996 -28767
rect 1966 -28827 1996 -28807
rect 2056 -28807 2106 -28767
rect 2056 -28827 2086 -28807
rect 2166 -28857 2226 -28597
rect 2156 -28867 2226 -28857
rect 1826 -28877 1906 -28867
rect 1826 -28937 1836 -28877
rect 1896 -28887 1906 -28877
rect 2146 -28877 2226 -28867
rect 2146 -28887 2156 -28877
rect 1896 -28937 2156 -28887
rect 2216 -28937 2226 -28877
rect 1826 -28947 2226 -28937
rect 2282 -28527 2682 -28517
rect 2282 -28587 2292 -28527
rect 2352 -28577 2612 -28527
rect 2352 -28587 2362 -28577
rect 2282 -28597 2362 -28587
rect 2602 -28587 2612 -28577
rect 2672 -28587 2682 -28527
rect 2602 -28597 2682 -28587
rect 2282 -28867 2342 -28597
rect 2422 -28657 2452 -28637
rect 2402 -28697 2452 -28657
rect 2512 -28657 2542 -28637
rect 2512 -28697 2562 -28657
rect 2402 -28767 2562 -28697
rect 2402 -28807 2452 -28767
rect 2422 -28827 2452 -28807
rect 2512 -28807 2562 -28767
rect 2512 -28827 2542 -28807
rect 2622 -28857 2682 -28597
rect 2612 -28867 2682 -28857
rect 2282 -28877 2362 -28867
rect 2282 -28937 2292 -28877
rect 2352 -28887 2362 -28877
rect 2602 -28877 2682 -28867
rect 2602 -28887 2612 -28877
rect 2352 -28937 2612 -28887
rect 2672 -28937 2682 -28877
rect 2282 -28947 2682 -28937
rect 2740 -28527 3140 -28517
rect 2740 -28587 2750 -28527
rect 2810 -28577 3070 -28527
rect 2810 -28587 2820 -28577
rect 2740 -28597 2820 -28587
rect 3060 -28587 3070 -28577
rect 3130 -28587 3140 -28527
rect 3060 -28597 3140 -28587
rect 2740 -28867 2800 -28597
rect 2880 -28657 2910 -28637
rect 2860 -28697 2910 -28657
rect 2970 -28657 3000 -28637
rect 2970 -28697 3020 -28657
rect 2860 -28767 3020 -28697
rect 2860 -28807 2910 -28767
rect 2880 -28827 2910 -28807
rect 2970 -28807 3020 -28767
rect 2970 -28827 3000 -28807
rect 3080 -28857 3140 -28597
rect 3070 -28867 3140 -28857
rect 2740 -28877 2820 -28867
rect 2740 -28937 2750 -28877
rect 2810 -28887 2820 -28877
rect 3060 -28877 3140 -28867
rect 3060 -28887 3070 -28877
rect 2810 -28937 3070 -28887
rect 3130 -28937 3140 -28877
rect 2740 -28947 3140 -28937
rect 3196 -28527 3596 -28517
rect 3196 -28587 3206 -28527
rect 3266 -28577 3526 -28527
rect 3266 -28587 3276 -28577
rect 3196 -28597 3276 -28587
rect 3516 -28587 3526 -28577
rect 3586 -28587 3596 -28527
rect 3516 -28597 3596 -28587
rect 3196 -28867 3256 -28597
rect 3336 -28657 3366 -28637
rect 3316 -28697 3366 -28657
rect 3426 -28657 3456 -28637
rect 3426 -28697 3476 -28657
rect 3316 -28767 3476 -28697
rect 3316 -28807 3366 -28767
rect 3336 -28827 3366 -28807
rect 3426 -28807 3476 -28767
rect 3426 -28827 3456 -28807
rect 3536 -28857 3596 -28597
rect 3526 -28867 3596 -28857
rect 3196 -28877 3276 -28867
rect 3196 -28937 3206 -28877
rect 3266 -28887 3276 -28877
rect 3516 -28877 3596 -28867
rect 3516 -28887 3526 -28877
rect 3266 -28937 3526 -28887
rect 3586 -28937 3596 -28877
rect 3196 -28947 3596 -28937
rect 3652 -28527 4052 -28517
rect 3652 -28587 3662 -28527
rect 3722 -28577 3982 -28527
rect 3722 -28587 3732 -28577
rect 3652 -28597 3732 -28587
rect 3972 -28587 3982 -28577
rect 4042 -28587 4052 -28527
rect 3972 -28597 4052 -28587
rect 3652 -28867 3712 -28597
rect 3792 -28657 3822 -28637
rect 3772 -28697 3822 -28657
rect 3882 -28657 3912 -28637
rect 3882 -28697 3932 -28657
rect 3772 -28767 3932 -28697
rect 3772 -28807 3822 -28767
rect 3792 -28827 3822 -28807
rect 3882 -28807 3932 -28767
rect 3882 -28827 3912 -28807
rect 3992 -28857 4052 -28597
rect 3982 -28867 4052 -28857
rect 3652 -28877 3732 -28867
rect 3652 -28937 3662 -28877
rect 3722 -28887 3732 -28877
rect 3972 -28877 4052 -28867
rect 3972 -28887 3982 -28877
rect 3722 -28937 3982 -28887
rect 4042 -28937 4052 -28877
rect 3652 -28947 4052 -28937
rect 4110 -28527 4510 -28517
rect 4110 -28587 4120 -28527
rect 4180 -28577 4440 -28527
rect 4180 -28587 4190 -28577
rect 4110 -28597 4190 -28587
rect 4430 -28587 4440 -28577
rect 4500 -28587 4510 -28527
rect 4430 -28597 4510 -28587
rect 4110 -28867 4170 -28597
rect 4250 -28657 4280 -28637
rect 4230 -28697 4280 -28657
rect 4340 -28657 4370 -28637
rect 4340 -28697 4390 -28657
rect 4230 -28767 4390 -28697
rect 4230 -28807 4280 -28767
rect 4250 -28827 4280 -28807
rect 4340 -28807 4390 -28767
rect 4340 -28827 4370 -28807
rect 4450 -28857 4510 -28597
rect 4440 -28867 4510 -28857
rect 4110 -28877 4190 -28867
rect 4110 -28937 4120 -28877
rect 4180 -28887 4190 -28877
rect 4430 -28877 4510 -28867
rect 4430 -28887 4440 -28877
rect 4180 -28937 4440 -28887
rect 4500 -28937 4510 -28877
rect 4110 -28947 4510 -28937
rect 4566 -28527 4966 -28517
rect 4566 -28587 4576 -28527
rect 4636 -28577 4896 -28527
rect 4636 -28587 4646 -28577
rect 4566 -28597 4646 -28587
rect 4886 -28587 4896 -28577
rect 4956 -28587 4966 -28527
rect 4886 -28597 4966 -28587
rect 4566 -28867 4626 -28597
rect 4706 -28657 4736 -28637
rect 4686 -28697 4736 -28657
rect 4796 -28657 4826 -28637
rect 4796 -28697 4846 -28657
rect 4686 -28767 4846 -28697
rect 4686 -28807 4736 -28767
rect 4706 -28827 4736 -28807
rect 4796 -28807 4846 -28767
rect 4796 -28827 4826 -28807
rect 4906 -28857 4966 -28597
rect 4896 -28867 4966 -28857
rect 4566 -28877 4646 -28867
rect 4566 -28937 4576 -28877
rect 4636 -28887 4646 -28877
rect 4886 -28877 4966 -28867
rect 4886 -28887 4896 -28877
rect 4636 -28937 4896 -28887
rect 4956 -28937 4966 -28877
rect 4566 -28947 4966 -28937
rect 5022 -28527 5422 -28517
rect 5022 -28587 5032 -28527
rect 5092 -28577 5352 -28527
rect 5092 -28587 5102 -28577
rect 5022 -28597 5102 -28587
rect 5342 -28587 5352 -28577
rect 5412 -28587 5422 -28527
rect 5342 -28597 5422 -28587
rect 5022 -28867 5082 -28597
rect 5162 -28657 5192 -28637
rect 5142 -28697 5192 -28657
rect 5252 -28657 5282 -28637
rect 5252 -28697 5302 -28657
rect 5142 -28767 5302 -28697
rect 5142 -28807 5192 -28767
rect 5162 -28827 5192 -28807
rect 5252 -28807 5302 -28767
rect 5252 -28827 5282 -28807
rect 5362 -28857 5422 -28597
rect 5352 -28867 5422 -28857
rect 5022 -28877 5102 -28867
rect 5022 -28937 5032 -28877
rect 5092 -28887 5102 -28877
rect 5342 -28877 5422 -28867
rect 5342 -28887 5352 -28877
rect 5092 -28937 5352 -28887
rect 5412 -28937 5422 -28877
rect 5022 -28947 5422 -28937
rect 5480 -28527 5880 -28517
rect 5480 -28587 5490 -28527
rect 5550 -28577 5810 -28527
rect 5550 -28587 5560 -28577
rect 5480 -28597 5560 -28587
rect 5800 -28587 5810 -28577
rect 5870 -28587 5880 -28527
rect 5800 -28597 5880 -28587
rect 5480 -28867 5540 -28597
rect 5620 -28657 5650 -28637
rect 5600 -28697 5650 -28657
rect 5710 -28657 5740 -28637
rect 5710 -28697 5760 -28657
rect 5600 -28767 5760 -28697
rect 5600 -28807 5650 -28767
rect 5620 -28827 5650 -28807
rect 5710 -28807 5760 -28767
rect 5710 -28827 5740 -28807
rect 5820 -28857 5880 -28597
rect 5810 -28867 5880 -28857
rect 5480 -28877 5560 -28867
rect 5480 -28937 5490 -28877
rect 5550 -28887 5560 -28877
rect 5800 -28877 5880 -28867
rect 5800 -28887 5810 -28877
rect 5550 -28937 5810 -28887
rect 5870 -28937 5880 -28877
rect 5480 -28947 5880 -28937
rect 5936 -28527 6336 -28517
rect 5936 -28587 5946 -28527
rect 6006 -28577 6266 -28527
rect 6006 -28587 6016 -28577
rect 5936 -28597 6016 -28587
rect 6256 -28587 6266 -28577
rect 6326 -28587 6336 -28527
rect 6256 -28597 6336 -28587
rect 5936 -28867 5996 -28597
rect 6076 -28657 6106 -28637
rect 6056 -28697 6106 -28657
rect 6166 -28657 6196 -28637
rect 6166 -28697 6216 -28657
rect 6056 -28767 6216 -28697
rect 6056 -28807 6106 -28767
rect 6076 -28827 6106 -28807
rect 6166 -28807 6216 -28767
rect 6166 -28827 6196 -28807
rect 6276 -28857 6336 -28597
rect 6266 -28867 6336 -28857
rect 5936 -28877 6016 -28867
rect 5936 -28937 5946 -28877
rect 6006 -28887 6016 -28877
rect 6256 -28877 6336 -28867
rect 6256 -28887 6266 -28877
rect 6006 -28937 6266 -28887
rect 6326 -28937 6336 -28877
rect 5936 -28947 6336 -28937
rect 6392 -28527 6792 -28517
rect 6392 -28587 6402 -28527
rect 6462 -28577 6722 -28527
rect 6462 -28587 6472 -28577
rect 6392 -28597 6472 -28587
rect 6712 -28587 6722 -28577
rect 6782 -28587 6792 -28527
rect 6712 -28597 6792 -28587
rect 6392 -28867 6452 -28597
rect 6532 -28657 6562 -28637
rect 6512 -28697 6562 -28657
rect 6622 -28657 6652 -28637
rect 6622 -28697 6672 -28657
rect 6512 -28767 6672 -28697
rect 6512 -28807 6562 -28767
rect 6532 -28827 6562 -28807
rect 6622 -28807 6672 -28767
rect 6622 -28827 6652 -28807
rect 6732 -28857 6792 -28597
rect 6722 -28867 6792 -28857
rect 6392 -28877 6472 -28867
rect 6392 -28937 6402 -28877
rect 6462 -28887 6472 -28877
rect 6712 -28877 6792 -28867
rect 6712 -28887 6722 -28877
rect 6462 -28937 6722 -28887
rect 6782 -28937 6792 -28877
rect 6392 -28947 6792 -28937
rect 6850 -28527 7250 -28517
rect 6850 -28587 6860 -28527
rect 6920 -28577 7180 -28527
rect 6920 -28587 6930 -28577
rect 6850 -28597 6930 -28587
rect 7170 -28587 7180 -28577
rect 7240 -28587 7250 -28527
rect 7170 -28597 7250 -28587
rect 6850 -28867 6910 -28597
rect 6990 -28657 7020 -28637
rect 6970 -28697 7020 -28657
rect 7080 -28657 7110 -28637
rect 7080 -28697 7130 -28657
rect 6970 -28767 7130 -28697
rect 6970 -28807 7020 -28767
rect 6990 -28827 7020 -28807
rect 7080 -28807 7130 -28767
rect 7080 -28827 7110 -28807
rect 7190 -28857 7250 -28597
rect 7180 -28867 7250 -28857
rect 6850 -28877 6930 -28867
rect 6850 -28937 6860 -28877
rect 6920 -28887 6930 -28877
rect 7170 -28877 7250 -28867
rect 7170 -28887 7180 -28877
rect 6920 -28937 7180 -28887
rect 7240 -28937 7250 -28877
rect 6850 -28947 7250 -28937
rect 7306 -28527 7706 -28517
rect 7306 -28587 7316 -28527
rect 7376 -28577 7636 -28527
rect 7376 -28587 7386 -28577
rect 7306 -28597 7386 -28587
rect 7626 -28587 7636 -28577
rect 7696 -28587 7706 -28527
rect 7626 -28597 7706 -28587
rect 7306 -28867 7366 -28597
rect 7446 -28657 7476 -28637
rect 7426 -28697 7476 -28657
rect 7536 -28657 7566 -28637
rect 7536 -28697 7586 -28657
rect 7426 -28767 7586 -28697
rect 7426 -28807 7476 -28767
rect 7446 -28827 7476 -28807
rect 7536 -28807 7586 -28767
rect 7536 -28827 7566 -28807
rect 7646 -28857 7706 -28597
rect 7636 -28867 7706 -28857
rect 7306 -28877 7386 -28867
rect 7306 -28937 7316 -28877
rect 7376 -28887 7386 -28877
rect 7626 -28877 7706 -28867
rect 7626 -28887 7636 -28877
rect 7376 -28937 7636 -28887
rect 7696 -28937 7706 -28877
rect 7306 -28947 7706 -28937
rect 7762 -28527 8162 -28517
rect 7762 -28587 7772 -28527
rect 7832 -28577 8092 -28527
rect 7832 -28587 7842 -28577
rect 7762 -28597 7842 -28587
rect 8082 -28587 8092 -28577
rect 8152 -28587 8162 -28527
rect 8082 -28597 8162 -28587
rect 7762 -28867 7822 -28597
rect 7902 -28657 7932 -28637
rect 7882 -28697 7932 -28657
rect 7992 -28657 8022 -28637
rect 7992 -28697 8042 -28657
rect 7882 -28767 8042 -28697
rect 7882 -28807 7932 -28767
rect 7902 -28827 7932 -28807
rect 7992 -28807 8042 -28767
rect 7992 -28827 8022 -28807
rect 8102 -28857 8162 -28597
rect 8092 -28867 8162 -28857
rect 7762 -28877 7842 -28867
rect 7762 -28937 7772 -28877
rect 7832 -28887 7842 -28877
rect 8082 -28877 8162 -28867
rect 8082 -28887 8092 -28877
rect 7832 -28937 8092 -28887
rect 8152 -28937 8162 -28877
rect 7762 -28947 8162 -28937
rect 8236 -28527 8636 -28517
rect 8236 -28587 8246 -28527
rect 8306 -28577 8566 -28527
rect 8306 -28587 8316 -28577
rect 8236 -28597 8316 -28587
rect 8556 -28587 8566 -28577
rect 8626 -28587 8636 -28527
rect 8556 -28597 8636 -28587
rect 8236 -28867 8296 -28597
rect 8376 -28657 8406 -28637
rect 8356 -28697 8406 -28657
rect 8466 -28657 8496 -28637
rect 8466 -28697 8516 -28657
rect 8356 -28767 8516 -28697
rect 8356 -28807 8406 -28767
rect 8376 -28827 8406 -28807
rect 8466 -28807 8516 -28767
rect 8466 -28827 8496 -28807
rect 8576 -28857 8636 -28597
rect 8566 -28867 8636 -28857
rect 8236 -28877 8316 -28867
rect 8236 -28937 8246 -28877
rect 8306 -28887 8316 -28877
rect 8556 -28877 8636 -28867
rect 8556 -28887 8566 -28877
rect 8306 -28937 8566 -28887
rect 8626 -28937 8636 -28877
rect 8236 -28947 8636 -28937
rect 8692 -28527 9092 -28517
rect 8692 -28587 8702 -28527
rect 8762 -28577 9022 -28527
rect 8762 -28587 8772 -28577
rect 8692 -28597 8772 -28587
rect 9012 -28587 9022 -28577
rect 9082 -28587 9092 -28527
rect 9012 -28597 9092 -28587
rect 8692 -28867 8752 -28597
rect 8832 -28657 8862 -28637
rect 8812 -28697 8862 -28657
rect 8922 -28657 8952 -28637
rect 8922 -28697 8972 -28657
rect 8812 -28767 8972 -28697
rect 8812 -28807 8862 -28767
rect 8832 -28827 8862 -28807
rect 8922 -28807 8972 -28767
rect 8922 -28827 8952 -28807
rect 9032 -28857 9092 -28597
rect 9022 -28867 9092 -28857
rect 8692 -28877 8772 -28867
rect 8692 -28937 8702 -28877
rect 8762 -28887 8772 -28877
rect 9012 -28877 9092 -28867
rect 9012 -28887 9022 -28877
rect 8762 -28937 9022 -28887
rect 9082 -28937 9092 -28877
rect 8692 -28947 9092 -28937
rect 9150 -28527 9550 -28517
rect 9150 -28587 9160 -28527
rect 9220 -28577 9480 -28527
rect 9220 -28587 9230 -28577
rect 9150 -28597 9230 -28587
rect 9470 -28587 9480 -28577
rect 9540 -28587 9550 -28527
rect 9470 -28597 9550 -28587
rect 9150 -28867 9210 -28597
rect 9290 -28657 9320 -28637
rect 9270 -28697 9320 -28657
rect 9380 -28657 9410 -28637
rect 9380 -28697 9430 -28657
rect 9270 -28767 9430 -28697
rect 9270 -28807 9320 -28767
rect 9290 -28827 9320 -28807
rect 9380 -28807 9430 -28767
rect 9380 -28827 9410 -28807
rect 9490 -28857 9550 -28597
rect 9480 -28867 9550 -28857
rect 9150 -28877 9230 -28867
rect 9150 -28937 9160 -28877
rect 9220 -28887 9230 -28877
rect 9470 -28877 9550 -28867
rect 9470 -28887 9480 -28877
rect 9220 -28937 9480 -28887
rect 9540 -28937 9550 -28877
rect 9150 -28947 9550 -28937
rect 9606 -28527 10006 -28517
rect 9606 -28587 9616 -28527
rect 9676 -28577 9936 -28527
rect 9676 -28587 9686 -28577
rect 9606 -28597 9686 -28587
rect 9926 -28587 9936 -28577
rect 9996 -28587 10006 -28527
rect 9926 -28597 10006 -28587
rect 9606 -28867 9666 -28597
rect 9746 -28657 9776 -28637
rect 9726 -28697 9776 -28657
rect 9836 -28657 9866 -28637
rect 9836 -28697 9886 -28657
rect 9726 -28767 9886 -28697
rect 9726 -28807 9776 -28767
rect 9746 -28827 9776 -28807
rect 9836 -28807 9886 -28767
rect 9836 -28827 9866 -28807
rect 9946 -28857 10006 -28597
rect 9936 -28867 10006 -28857
rect 9606 -28877 9686 -28867
rect 9606 -28937 9616 -28877
rect 9676 -28887 9686 -28877
rect 9926 -28877 10006 -28867
rect 9926 -28887 9936 -28877
rect 9676 -28937 9936 -28887
rect 9996 -28937 10006 -28877
rect 9606 -28947 10006 -28937
rect 10062 -28527 10462 -28517
rect 10062 -28587 10072 -28527
rect 10132 -28577 10392 -28527
rect 10132 -28587 10142 -28577
rect 10062 -28597 10142 -28587
rect 10382 -28587 10392 -28577
rect 10452 -28587 10462 -28527
rect 10382 -28597 10462 -28587
rect 10062 -28867 10122 -28597
rect 10202 -28657 10232 -28637
rect 10182 -28697 10232 -28657
rect 10292 -28657 10322 -28637
rect 10292 -28697 10342 -28657
rect 10182 -28767 10342 -28697
rect 10182 -28807 10232 -28767
rect 10202 -28827 10232 -28807
rect 10292 -28807 10342 -28767
rect 10292 -28827 10322 -28807
rect 10402 -28857 10462 -28597
rect 10392 -28867 10462 -28857
rect 10062 -28877 10142 -28867
rect 10062 -28937 10072 -28877
rect 10132 -28887 10142 -28877
rect 10382 -28877 10462 -28867
rect 10382 -28887 10392 -28877
rect 10132 -28937 10392 -28887
rect 10452 -28937 10462 -28877
rect 10062 -28947 10462 -28937
rect 10520 -28527 10920 -28517
rect 10520 -28587 10530 -28527
rect 10590 -28577 10850 -28527
rect 10590 -28587 10600 -28577
rect 10520 -28597 10600 -28587
rect 10840 -28587 10850 -28577
rect 10910 -28587 10920 -28527
rect 10840 -28597 10920 -28587
rect 10520 -28867 10580 -28597
rect 10660 -28657 10690 -28637
rect 10640 -28697 10690 -28657
rect 10750 -28657 10780 -28637
rect 10750 -28697 10800 -28657
rect 10640 -28767 10800 -28697
rect 10640 -28807 10690 -28767
rect 10660 -28827 10690 -28807
rect 10750 -28807 10800 -28767
rect 10750 -28827 10780 -28807
rect 10860 -28857 10920 -28597
rect 10850 -28867 10920 -28857
rect 10520 -28877 10600 -28867
rect 10520 -28937 10530 -28877
rect 10590 -28887 10600 -28877
rect 10840 -28877 10920 -28867
rect 10840 -28887 10850 -28877
rect 10590 -28937 10850 -28887
rect 10910 -28937 10920 -28877
rect 10520 -28947 10920 -28937
rect 10976 -28527 11376 -28517
rect 10976 -28587 10986 -28527
rect 11046 -28577 11306 -28527
rect 11046 -28587 11056 -28577
rect 10976 -28597 11056 -28587
rect 11296 -28587 11306 -28577
rect 11366 -28587 11376 -28527
rect 11296 -28597 11376 -28587
rect 10976 -28867 11036 -28597
rect 11116 -28657 11146 -28637
rect 11096 -28697 11146 -28657
rect 11206 -28657 11236 -28637
rect 11206 -28697 11256 -28657
rect 11096 -28767 11256 -28697
rect 11096 -28807 11146 -28767
rect 11116 -28827 11146 -28807
rect 11206 -28807 11256 -28767
rect 11206 -28827 11236 -28807
rect 11316 -28857 11376 -28597
rect 11306 -28867 11376 -28857
rect 10976 -28877 11056 -28867
rect 10976 -28937 10986 -28877
rect 11046 -28887 11056 -28877
rect 11296 -28877 11376 -28867
rect 11296 -28887 11306 -28877
rect 11046 -28937 11306 -28887
rect 11366 -28937 11376 -28877
rect 10976 -28947 11376 -28937
rect 11432 -28527 11832 -28517
rect 11432 -28587 11442 -28527
rect 11502 -28577 11762 -28527
rect 11502 -28587 11512 -28577
rect 11432 -28597 11512 -28587
rect 11752 -28587 11762 -28577
rect 11822 -28587 11832 -28527
rect 11752 -28597 11832 -28587
rect 11432 -28867 11492 -28597
rect 11572 -28657 11602 -28637
rect 11552 -28697 11602 -28657
rect 11662 -28657 11692 -28637
rect 11662 -28697 11712 -28657
rect 11552 -28767 11712 -28697
rect 11552 -28807 11602 -28767
rect 11572 -28827 11602 -28807
rect 11662 -28807 11712 -28767
rect 11662 -28827 11692 -28807
rect 11772 -28857 11832 -28597
rect 11762 -28867 11832 -28857
rect 11432 -28877 11512 -28867
rect 11432 -28937 11442 -28877
rect 11502 -28887 11512 -28877
rect 11752 -28877 11832 -28867
rect 11752 -28887 11762 -28877
rect 11502 -28937 11762 -28887
rect 11822 -28937 11832 -28877
rect 11432 -28947 11832 -28937
rect 11890 -28527 12290 -28517
rect 11890 -28587 11900 -28527
rect 11960 -28577 12220 -28527
rect 11960 -28587 11970 -28577
rect 11890 -28597 11970 -28587
rect 12210 -28587 12220 -28577
rect 12280 -28587 12290 -28527
rect 12210 -28597 12290 -28587
rect 11890 -28867 11950 -28597
rect 12030 -28657 12060 -28637
rect 12010 -28697 12060 -28657
rect 12120 -28657 12150 -28637
rect 12120 -28697 12170 -28657
rect 12010 -28767 12170 -28697
rect 12010 -28807 12060 -28767
rect 12030 -28827 12060 -28807
rect 12120 -28807 12170 -28767
rect 12120 -28827 12150 -28807
rect 12230 -28857 12290 -28597
rect 12220 -28867 12290 -28857
rect 11890 -28877 11970 -28867
rect 11890 -28937 11900 -28877
rect 11960 -28887 11970 -28877
rect 12210 -28877 12290 -28867
rect 12210 -28887 12220 -28877
rect 11960 -28937 12220 -28887
rect 12280 -28937 12290 -28877
rect 11890 -28947 12290 -28937
rect 12346 -28527 12746 -28517
rect 12346 -28587 12356 -28527
rect 12416 -28577 12676 -28527
rect 12416 -28587 12426 -28577
rect 12346 -28597 12426 -28587
rect 12666 -28587 12676 -28577
rect 12736 -28587 12746 -28527
rect 12666 -28597 12746 -28587
rect 12346 -28867 12406 -28597
rect 12486 -28657 12516 -28637
rect 12466 -28697 12516 -28657
rect 12576 -28657 12606 -28637
rect 12576 -28697 12626 -28657
rect 12466 -28767 12626 -28697
rect 12466 -28807 12516 -28767
rect 12486 -28827 12516 -28807
rect 12576 -28807 12626 -28767
rect 12576 -28827 12606 -28807
rect 12686 -28857 12746 -28597
rect 12676 -28867 12746 -28857
rect 12346 -28877 12426 -28867
rect 12346 -28937 12356 -28877
rect 12416 -28887 12426 -28877
rect 12666 -28877 12746 -28867
rect 12666 -28887 12676 -28877
rect 12416 -28937 12676 -28887
rect 12736 -28937 12746 -28877
rect 12346 -28947 12746 -28937
rect 12802 -28527 13202 -28517
rect 12802 -28587 12812 -28527
rect 12872 -28577 13132 -28527
rect 12872 -28587 12882 -28577
rect 12802 -28597 12882 -28587
rect 13122 -28587 13132 -28577
rect 13192 -28587 13202 -28527
rect 13122 -28597 13202 -28587
rect 12802 -28867 12862 -28597
rect 12942 -28657 12972 -28637
rect 12922 -28697 12972 -28657
rect 13032 -28657 13062 -28637
rect 13032 -28697 13082 -28657
rect 12922 -28767 13082 -28697
rect 12922 -28807 12972 -28767
rect 12942 -28827 12972 -28807
rect 13032 -28807 13082 -28767
rect 13032 -28827 13062 -28807
rect 13142 -28857 13202 -28597
rect 13132 -28867 13202 -28857
rect 12802 -28877 12882 -28867
rect 12802 -28937 12812 -28877
rect 12872 -28887 12882 -28877
rect 13122 -28877 13202 -28867
rect 13122 -28887 13132 -28877
rect 12872 -28937 13132 -28887
rect 13192 -28937 13202 -28877
rect 12802 -28947 13202 -28937
rect 13260 -28527 13660 -28517
rect 13260 -28587 13270 -28527
rect 13330 -28577 13590 -28527
rect 13330 -28587 13340 -28577
rect 13260 -28597 13340 -28587
rect 13580 -28587 13590 -28577
rect 13650 -28587 13660 -28527
rect 13580 -28597 13660 -28587
rect 13260 -28867 13320 -28597
rect 13400 -28657 13430 -28637
rect 13380 -28697 13430 -28657
rect 13490 -28657 13520 -28637
rect 13490 -28697 13540 -28657
rect 13380 -28767 13540 -28697
rect 13380 -28807 13430 -28767
rect 13400 -28827 13430 -28807
rect 13490 -28807 13540 -28767
rect 13490 -28827 13520 -28807
rect 13600 -28857 13660 -28597
rect 13590 -28867 13660 -28857
rect 13260 -28877 13340 -28867
rect 13260 -28937 13270 -28877
rect 13330 -28887 13340 -28877
rect 13580 -28877 13660 -28867
rect 13580 -28887 13590 -28877
rect 13330 -28937 13590 -28887
rect 13650 -28937 13660 -28877
rect 13260 -28947 13660 -28937
rect 13716 -28527 14116 -28517
rect 13716 -28587 13726 -28527
rect 13786 -28577 14046 -28527
rect 13786 -28587 13796 -28577
rect 13716 -28597 13796 -28587
rect 14036 -28587 14046 -28577
rect 14106 -28587 14116 -28527
rect 14036 -28597 14116 -28587
rect 13716 -28867 13776 -28597
rect 13856 -28657 13886 -28637
rect 13836 -28697 13886 -28657
rect 13946 -28657 13976 -28637
rect 13946 -28697 13996 -28657
rect 13836 -28767 13996 -28697
rect 13836 -28807 13886 -28767
rect 13856 -28827 13886 -28807
rect 13946 -28807 13996 -28767
rect 13946 -28827 13976 -28807
rect 14056 -28857 14116 -28597
rect 14046 -28867 14116 -28857
rect 13716 -28877 13796 -28867
rect 13716 -28937 13726 -28877
rect 13786 -28887 13796 -28877
rect 14036 -28877 14116 -28867
rect 14036 -28887 14046 -28877
rect 13786 -28937 14046 -28887
rect 14106 -28937 14116 -28877
rect 13716 -28947 14116 -28937
rect 14172 -28527 14572 -28517
rect 14172 -28587 14182 -28527
rect 14242 -28577 14502 -28527
rect 14242 -28587 14252 -28577
rect 14172 -28597 14252 -28587
rect 14492 -28587 14502 -28577
rect 14562 -28587 14572 -28527
rect 14492 -28597 14572 -28587
rect 14172 -28867 14232 -28597
rect 14312 -28657 14342 -28637
rect 14292 -28697 14342 -28657
rect 14402 -28657 14432 -28637
rect 14402 -28697 14452 -28657
rect 14292 -28767 14452 -28697
rect 14292 -28807 14342 -28767
rect 14312 -28827 14342 -28807
rect 14402 -28807 14452 -28767
rect 14402 -28827 14432 -28807
rect 14512 -28857 14572 -28597
rect 14502 -28867 14572 -28857
rect 14172 -28877 14252 -28867
rect 14172 -28937 14182 -28877
rect 14242 -28887 14252 -28877
rect 14492 -28877 14572 -28867
rect 14492 -28887 14502 -28877
rect 14242 -28937 14502 -28887
rect 14562 -28937 14572 -28877
rect 14172 -28947 14572 -28937
rect 14630 -28527 15030 -28517
rect 14630 -28587 14640 -28527
rect 14700 -28577 14960 -28527
rect 14700 -28587 14710 -28577
rect 14630 -28597 14710 -28587
rect 14950 -28587 14960 -28577
rect 15020 -28587 15030 -28527
rect 14950 -28597 15030 -28587
rect 14630 -28867 14690 -28597
rect 14770 -28657 14800 -28637
rect 14750 -28697 14800 -28657
rect 14860 -28657 14890 -28637
rect 14860 -28697 14910 -28657
rect 14750 -28767 14910 -28697
rect 14750 -28807 14800 -28767
rect 14770 -28827 14800 -28807
rect 14860 -28807 14910 -28767
rect 14860 -28827 14890 -28807
rect 14970 -28857 15030 -28597
rect 14960 -28867 15030 -28857
rect 14630 -28877 14710 -28867
rect 14630 -28937 14640 -28877
rect 14700 -28887 14710 -28877
rect 14950 -28877 15030 -28867
rect 14950 -28887 14960 -28877
rect 14700 -28937 14960 -28887
rect 15020 -28937 15030 -28877
rect 14630 -28947 15030 -28937
rect 15086 -28527 15486 -28517
rect 15086 -28587 15096 -28527
rect 15156 -28577 15416 -28527
rect 15156 -28587 15166 -28577
rect 15086 -28597 15166 -28587
rect 15406 -28587 15416 -28577
rect 15476 -28587 15486 -28527
rect 15406 -28597 15486 -28587
rect 15086 -28867 15146 -28597
rect 15226 -28657 15256 -28637
rect 15206 -28697 15256 -28657
rect 15316 -28657 15346 -28637
rect 15316 -28697 15366 -28657
rect 15206 -28767 15366 -28697
rect 15206 -28807 15256 -28767
rect 15226 -28827 15256 -28807
rect 15316 -28807 15366 -28767
rect 15316 -28827 15346 -28807
rect 15426 -28857 15486 -28597
rect 15416 -28867 15486 -28857
rect 15086 -28877 15166 -28867
rect 15086 -28937 15096 -28877
rect 15156 -28887 15166 -28877
rect 15406 -28877 15486 -28867
rect 15406 -28887 15416 -28877
rect 15156 -28937 15416 -28887
rect 15476 -28937 15486 -28877
rect 15086 -28947 15486 -28937
rect 0 -29021 400 -29011
rect 0 -29081 10 -29021
rect 70 -29071 330 -29021
rect 70 -29081 80 -29071
rect 0 -29091 80 -29081
rect 320 -29081 330 -29071
rect 390 -29081 400 -29021
rect 320 -29091 400 -29081
rect 0 -29361 60 -29091
rect 140 -29151 170 -29131
rect 120 -29191 170 -29151
rect 230 -29151 260 -29131
rect 230 -29191 280 -29151
rect 120 -29261 280 -29191
rect 120 -29301 170 -29261
rect 140 -29321 170 -29301
rect 230 -29301 280 -29261
rect 230 -29321 260 -29301
rect 340 -29351 400 -29091
rect 330 -29361 400 -29351
rect 0 -29371 80 -29361
rect 0 -29431 10 -29371
rect 70 -29381 80 -29371
rect 320 -29371 400 -29361
rect 320 -29381 330 -29371
rect 70 -29431 330 -29381
rect 390 -29431 400 -29371
rect 0 -29441 400 -29431
rect 456 -29021 856 -29011
rect 456 -29081 466 -29021
rect 526 -29071 786 -29021
rect 526 -29081 536 -29071
rect 456 -29091 536 -29081
rect 776 -29081 786 -29071
rect 846 -29081 856 -29021
rect 776 -29091 856 -29081
rect 456 -29361 516 -29091
rect 596 -29151 626 -29131
rect 576 -29191 626 -29151
rect 686 -29151 716 -29131
rect 686 -29191 736 -29151
rect 576 -29261 736 -29191
rect 576 -29301 626 -29261
rect 596 -29321 626 -29301
rect 686 -29301 736 -29261
rect 686 -29321 716 -29301
rect 796 -29351 856 -29091
rect 786 -29361 856 -29351
rect 456 -29371 536 -29361
rect 456 -29431 466 -29371
rect 526 -29381 536 -29371
rect 776 -29371 856 -29361
rect 776 -29381 786 -29371
rect 526 -29431 786 -29381
rect 846 -29431 856 -29371
rect 456 -29441 856 -29431
rect 912 -29021 1312 -29011
rect 912 -29081 922 -29021
rect 982 -29071 1242 -29021
rect 982 -29081 992 -29071
rect 912 -29091 992 -29081
rect 1232 -29081 1242 -29071
rect 1302 -29081 1312 -29021
rect 1232 -29091 1312 -29081
rect 912 -29361 972 -29091
rect 1052 -29151 1082 -29131
rect 1032 -29191 1082 -29151
rect 1142 -29151 1172 -29131
rect 1142 -29191 1192 -29151
rect 1032 -29261 1192 -29191
rect 1032 -29301 1082 -29261
rect 1052 -29321 1082 -29301
rect 1142 -29301 1192 -29261
rect 1142 -29321 1172 -29301
rect 1252 -29351 1312 -29091
rect 1242 -29361 1312 -29351
rect 912 -29371 992 -29361
rect 912 -29431 922 -29371
rect 982 -29381 992 -29371
rect 1232 -29371 1312 -29361
rect 1232 -29381 1242 -29371
rect 982 -29431 1242 -29381
rect 1302 -29431 1312 -29371
rect 912 -29441 1312 -29431
rect 1370 -29021 1770 -29011
rect 1370 -29081 1380 -29021
rect 1440 -29071 1700 -29021
rect 1440 -29081 1450 -29071
rect 1370 -29091 1450 -29081
rect 1690 -29081 1700 -29071
rect 1760 -29081 1770 -29021
rect 1690 -29091 1770 -29081
rect 1370 -29361 1430 -29091
rect 1510 -29151 1540 -29131
rect 1490 -29191 1540 -29151
rect 1600 -29151 1630 -29131
rect 1600 -29191 1650 -29151
rect 1490 -29261 1650 -29191
rect 1490 -29301 1540 -29261
rect 1510 -29321 1540 -29301
rect 1600 -29301 1650 -29261
rect 1600 -29321 1630 -29301
rect 1710 -29351 1770 -29091
rect 1700 -29361 1770 -29351
rect 1370 -29371 1450 -29361
rect 1370 -29431 1380 -29371
rect 1440 -29381 1450 -29371
rect 1690 -29371 1770 -29361
rect 1690 -29381 1700 -29371
rect 1440 -29431 1700 -29381
rect 1760 -29431 1770 -29371
rect 1370 -29441 1770 -29431
rect 1826 -29021 2226 -29011
rect 1826 -29081 1836 -29021
rect 1896 -29071 2156 -29021
rect 1896 -29081 1906 -29071
rect 1826 -29091 1906 -29081
rect 2146 -29081 2156 -29071
rect 2216 -29081 2226 -29021
rect 2146 -29091 2226 -29081
rect 1826 -29361 1886 -29091
rect 1966 -29151 1996 -29131
rect 1946 -29191 1996 -29151
rect 2056 -29151 2086 -29131
rect 2056 -29191 2106 -29151
rect 1946 -29261 2106 -29191
rect 1946 -29301 1996 -29261
rect 1966 -29321 1996 -29301
rect 2056 -29301 2106 -29261
rect 2056 -29321 2086 -29301
rect 2166 -29351 2226 -29091
rect 2156 -29361 2226 -29351
rect 1826 -29371 1906 -29361
rect 1826 -29431 1836 -29371
rect 1896 -29381 1906 -29371
rect 2146 -29371 2226 -29361
rect 2146 -29381 2156 -29371
rect 1896 -29431 2156 -29381
rect 2216 -29431 2226 -29371
rect 1826 -29441 2226 -29431
rect 2282 -29021 2682 -29011
rect 2282 -29081 2292 -29021
rect 2352 -29071 2612 -29021
rect 2352 -29081 2362 -29071
rect 2282 -29091 2362 -29081
rect 2602 -29081 2612 -29071
rect 2672 -29081 2682 -29021
rect 2602 -29091 2682 -29081
rect 2282 -29361 2342 -29091
rect 2422 -29151 2452 -29131
rect 2402 -29191 2452 -29151
rect 2512 -29151 2542 -29131
rect 2512 -29191 2562 -29151
rect 2402 -29261 2562 -29191
rect 2402 -29301 2452 -29261
rect 2422 -29321 2452 -29301
rect 2512 -29301 2562 -29261
rect 2512 -29321 2542 -29301
rect 2622 -29351 2682 -29091
rect 2612 -29361 2682 -29351
rect 2282 -29371 2362 -29361
rect 2282 -29431 2292 -29371
rect 2352 -29381 2362 -29371
rect 2602 -29371 2682 -29361
rect 2602 -29381 2612 -29371
rect 2352 -29431 2612 -29381
rect 2672 -29431 2682 -29371
rect 2282 -29441 2682 -29431
rect 2740 -29021 3140 -29011
rect 2740 -29081 2750 -29021
rect 2810 -29071 3070 -29021
rect 2810 -29081 2820 -29071
rect 2740 -29091 2820 -29081
rect 3060 -29081 3070 -29071
rect 3130 -29081 3140 -29021
rect 3060 -29091 3140 -29081
rect 2740 -29361 2800 -29091
rect 2880 -29151 2910 -29131
rect 2860 -29191 2910 -29151
rect 2970 -29151 3000 -29131
rect 2970 -29191 3020 -29151
rect 2860 -29261 3020 -29191
rect 2860 -29301 2910 -29261
rect 2880 -29321 2910 -29301
rect 2970 -29301 3020 -29261
rect 2970 -29321 3000 -29301
rect 3080 -29351 3140 -29091
rect 3070 -29361 3140 -29351
rect 2740 -29371 2820 -29361
rect 2740 -29431 2750 -29371
rect 2810 -29381 2820 -29371
rect 3060 -29371 3140 -29361
rect 3060 -29381 3070 -29371
rect 2810 -29431 3070 -29381
rect 3130 -29431 3140 -29371
rect 2740 -29441 3140 -29431
rect 3196 -29021 3596 -29011
rect 3196 -29081 3206 -29021
rect 3266 -29071 3526 -29021
rect 3266 -29081 3276 -29071
rect 3196 -29091 3276 -29081
rect 3516 -29081 3526 -29071
rect 3586 -29081 3596 -29021
rect 3516 -29091 3596 -29081
rect 3196 -29361 3256 -29091
rect 3336 -29151 3366 -29131
rect 3316 -29191 3366 -29151
rect 3426 -29151 3456 -29131
rect 3426 -29191 3476 -29151
rect 3316 -29261 3476 -29191
rect 3316 -29301 3366 -29261
rect 3336 -29321 3366 -29301
rect 3426 -29301 3476 -29261
rect 3426 -29321 3456 -29301
rect 3536 -29351 3596 -29091
rect 3526 -29361 3596 -29351
rect 3196 -29371 3276 -29361
rect 3196 -29431 3206 -29371
rect 3266 -29381 3276 -29371
rect 3516 -29371 3596 -29361
rect 3516 -29381 3526 -29371
rect 3266 -29431 3526 -29381
rect 3586 -29431 3596 -29371
rect 3196 -29441 3596 -29431
rect 3652 -29021 4052 -29011
rect 3652 -29081 3662 -29021
rect 3722 -29071 3982 -29021
rect 3722 -29081 3732 -29071
rect 3652 -29091 3732 -29081
rect 3972 -29081 3982 -29071
rect 4042 -29081 4052 -29021
rect 3972 -29091 4052 -29081
rect 3652 -29361 3712 -29091
rect 3792 -29151 3822 -29131
rect 3772 -29191 3822 -29151
rect 3882 -29151 3912 -29131
rect 3882 -29191 3932 -29151
rect 3772 -29261 3932 -29191
rect 3772 -29301 3822 -29261
rect 3792 -29321 3822 -29301
rect 3882 -29301 3932 -29261
rect 3882 -29321 3912 -29301
rect 3992 -29351 4052 -29091
rect 3982 -29361 4052 -29351
rect 3652 -29371 3732 -29361
rect 3652 -29431 3662 -29371
rect 3722 -29381 3732 -29371
rect 3972 -29371 4052 -29361
rect 3972 -29381 3982 -29371
rect 3722 -29431 3982 -29381
rect 4042 -29431 4052 -29371
rect 3652 -29441 4052 -29431
rect 4110 -29021 4510 -29011
rect 4110 -29081 4120 -29021
rect 4180 -29071 4440 -29021
rect 4180 -29081 4190 -29071
rect 4110 -29091 4190 -29081
rect 4430 -29081 4440 -29071
rect 4500 -29081 4510 -29021
rect 4430 -29091 4510 -29081
rect 4110 -29361 4170 -29091
rect 4250 -29151 4280 -29131
rect 4230 -29191 4280 -29151
rect 4340 -29151 4370 -29131
rect 4340 -29191 4390 -29151
rect 4230 -29261 4390 -29191
rect 4230 -29301 4280 -29261
rect 4250 -29321 4280 -29301
rect 4340 -29301 4390 -29261
rect 4340 -29321 4370 -29301
rect 4450 -29351 4510 -29091
rect 4440 -29361 4510 -29351
rect 4110 -29371 4190 -29361
rect 4110 -29431 4120 -29371
rect 4180 -29381 4190 -29371
rect 4430 -29371 4510 -29361
rect 4430 -29381 4440 -29371
rect 4180 -29431 4440 -29381
rect 4500 -29431 4510 -29371
rect 4110 -29441 4510 -29431
rect 4566 -29021 4966 -29011
rect 4566 -29081 4576 -29021
rect 4636 -29071 4896 -29021
rect 4636 -29081 4646 -29071
rect 4566 -29091 4646 -29081
rect 4886 -29081 4896 -29071
rect 4956 -29081 4966 -29021
rect 4886 -29091 4966 -29081
rect 4566 -29361 4626 -29091
rect 4706 -29151 4736 -29131
rect 4686 -29191 4736 -29151
rect 4796 -29151 4826 -29131
rect 4796 -29191 4846 -29151
rect 4686 -29261 4846 -29191
rect 4686 -29301 4736 -29261
rect 4706 -29321 4736 -29301
rect 4796 -29301 4846 -29261
rect 4796 -29321 4826 -29301
rect 4906 -29351 4966 -29091
rect 4896 -29361 4966 -29351
rect 4566 -29371 4646 -29361
rect 4566 -29431 4576 -29371
rect 4636 -29381 4646 -29371
rect 4886 -29371 4966 -29361
rect 4886 -29381 4896 -29371
rect 4636 -29431 4896 -29381
rect 4956 -29431 4966 -29371
rect 4566 -29441 4966 -29431
rect 5022 -29021 5422 -29011
rect 5022 -29081 5032 -29021
rect 5092 -29071 5352 -29021
rect 5092 -29081 5102 -29071
rect 5022 -29091 5102 -29081
rect 5342 -29081 5352 -29071
rect 5412 -29081 5422 -29021
rect 5342 -29091 5422 -29081
rect 5022 -29361 5082 -29091
rect 5162 -29151 5192 -29131
rect 5142 -29191 5192 -29151
rect 5252 -29151 5282 -29131
rect 5252 -29191 5302 -29151
rect 5142 -29261 5302 -29191
rect 5142 -29301 5192 -29261
rect 5162 -29321 5192 -29301
rect 5252 -29301 5302 -29261
rect 5252 -29321 5282 -29301
rect 5362 -29351 5422 -29091
rect 5352 -29361 5422 -29351
rect 5022 -29371 5102 -29361
rect 5022 -29431 5032 -29371
rect 5092 -29381 5102 -29371
rect 5342 -29371 5422 -29361
rect 5342 -29381 5352 -29371
rect 5092 -29431 5352 -29381
rect 5412 -29431 5422 -29371
rect 5022 -29441 5422 -29431
rect 5480 -29021 5880 -29011
rect 5480 -29081 5490 -29021
rect 5550 -29071 5810 -29021
rect 5550 -29081 5560 -29071
rect 5480 -29091 5560 -29081
rect 5800 -29081 5810 -29071
rect 5870 -29081 5880 -29021
rect 5800 -29091 5880 -29081
rect 5480 -29361 5540 -29091
rect 5620 -29151 5650 -29131
rect 5600 -29191 5650 -29151
rect 5710 -29151 5740 -29131
rect 5710 -29191 5760 -29151
rect 5600 -29261 5760 -29191
rect 5600 -29301 5650 -29261
rect 5620 -29321 5650 -29301
rect 5710 -29301 5760 -29261
rect 5710 -29321 5740 -29301
rect 5820 -29351 5880 -29091
rect 5810 -29361 5880 -29351
rect 5480 -29371 5560 -29361
rect 5480 -29431 5490 -29371
rect 5550 -29381 5560 -29371
rect 5800 -29371 5880 -29361
rect 5800 -29381 5810 -29371
rect 5550 -29431 5810 -29381
rect 5870 -29431 5880 -29371
rect 5480 -29441 5880 -29431
rect 5936 -29021 6336 -29011
rect 5936 -29081 5946 -29021
rect 6006 -29071 6266 -29021
rect 6006 -29081 6016 -29071
rect 5936 -29091 6016 -29081
rect 6256 -29081 6266 -29071
rect 6326 -29081 6336 -29021
rect 6256 -29091 6336 -29081
rect 5936 -29361 5996 -29091
rect 6076 -29151 6106 -29131
rect 6056 -29191 6106 -29151
rect 6166 -29151 6196 -29131
rect 6166 -29191 6216 -29151
rect 6056 -29261 6216 -29191
rect 6056 -29301 6106 -29261
rect 6076 -29321 6106 -29301
rect 6166 -29301 6216 -29261
rect 6166 -29321 6196 -29301
rect 6276 -29351 6336 -29091
rect 6266 -29361 6336 -29351
rect 5936 -29371 6016 -29361
rect 5936 -29431 5946 -29371
rect 6006 -29381 6016 -29371
rect 6256 -29371 6336 -29361
rect 6256 -29381 6266 -29371
rect 6006 -29431 6266 -29381
rect 6326 -29431 6336 -29371
rect 5936 -29441 6336 -29431
rect 6392 -29021 6792 -29011
rect 6392 -29081 6402 -29021
rect 6462 -29071 6722 -29021
rect 6462 -29081 6472 -29071
rect 6392 -29091 6472 -29081
rect 6712 -29081 6722 -29071
rect 6782 -29081 6792 -29021
rect 6712 -29091 6792 -29081
rect 6392 -29361 6452 -29091
rect 6532 -29151 6562 -29131
rect 6512 -29191 6562 -29151
rect 6622 -29151 6652 -29131
rect 6622 -29191 6672 -29151
rect 6512 -29261 6672 -29191
rect 6512 -29301 6562 -29261
rect 6532 -29321 6562 -29301
rect 6622 -29301 6672 -29261
rect 6622 -29321 6652 -29301
rect 6732 -29351 6792 -29091
rect 6722 -29361 6792 -29351
rect 6392 -29371 6472 -29361
rect 6392 -29431 6402 -29371
rect 6462 -29381 6472 -29371
rect 6712 -29371 6792 -29361
rect 6712 -29381 6722 -29371
rect 6462 -29431 6722 -29381
rect 6782 -29431 6792 -29371
rect 6392 -29441 6792 -29431
rect 6850 -29021 7250 -29011
rect 6850 -29081 6860 -29021
rect 6920 -29071 7180 -29021
rect 6920 -29081 6930 -29071
rect 6850 -29091 6930 -29081
rect 7170 -29081 7180 -29071
rect 7240 -29081 7250 -29021
rect 7170 -29091 7250 -29081
rect 6850 -29361 6910 -29091
rect 6990 -29151 7020 -29131
rect 6970 -29191 7020 -29151
rect 7080 -29151 7110 -29131
rect 7080 -29191 7130 -29151
rect 6970 -29261 7130 -29191
rect 6970 -29301 7020 -29261
rect 6990 -29321 7020 -29301
rect 7080 -29301 7130 -29261
rect 7080 -29321 7110 -29301
rect 7190 -29351 7250 -29091
rect 7180 -29361 7250 -29351
rect 6850 -29371 6930 -29361
rect 6850 -29431 6860 -29371
rect 6920 -29381 6930 -29371
rect 7170 -29371 7250 -29361
rect 7170 -29381 7180 -29371
rect 6920 -29431 7180 -29381
rect 7240 -29431 7250 -29371
rect 6850 -29441 7250 -29431
rect 7306 -29021 7706 -29011
rect 7306 -29081 7316 -29021
rect 7376 -29071 7636 -29021
rect 7376 -29081 7386 -29071
rect 7306 -29091 7386 -29081
rect 7626 -29081 7636 -29071
rect 7696 -29081 7706 -29021
rect 7626 -29091 7706 -29081
rect 7306 -29361 7366 -29091
rect 7446 -29151 7476 -29131
rect 7426 -29191 7476 -29151
rect 7536 -29151 7566 -29131
rect 7536 -29191 7586 -29151
rect 7426 -29261 7586 -29191
rect 7426 -29301 7476 -29261
rect 7446 -29321 7476 -29301
rect 7536 -29301 7586 -29261
rect 7536 -29321 7566 -29301
rect 7646 -29351 7706 -29091
rect 7636 -29361 7706 -29351
rect 7306 -29371 7386 -29361
rect 7306 -29431 7316 -29371
rect 7376 -29381 7386 -29371
rect 7626 -29371 7706 -29361
rect 7626 -29381 7636 -29371
rect 7376 -29431 7636 -29381
rect 7696 -29431 7706 -29371
rect 7306 -29441 7706 -29431
rect 7762 -29021 8162 -29011
rect 7762 -29081 7772 -29021
rect 7832 -29071 8092 -29021
rect 7832 -29081 7842 -29071
rect 7762 -29091 7842 -29081
rect 8082 -29081 8092 -29071
rect 8152 -29081 8162 -29021
rect 8082 -29091 8162 -29081
rect 7762 -29361 7822 -29091
rect 7902 -29151 7932 -29131
rect 7882 -29191 7932 -29151
rect 7992 -29151 8022 -29131
rect 7992 -29191 8042 -29151
rect 7882 -29261 8042 -29191
rect 7882 -29301 7932 -29261
rect 7902 -29321 7932 -29301
rect 7992 -29301 8042 -29261
rect 7992 -29321 8022 -29301
rect 8102 -29351 8162 -29091
rect 8092 -29361 8162 -29351
rect 7762 -29371 7842 -29361
rect 7762 -29431 7772 -29371
rect 7832 -29381 7842 -29371
rect 8082 -29371 8162 -29361
rect 8082 -29381 8092 -29371
rect 7832 -29431 8092 -29381
rect 8152 -29431 8162 -29371
rect 7762 -29441 8162 -29431
rect 8236 -29021 8636 -29011
rect 8236 -29081 8246 -29021
rect 8306 -29071 8566 -29021
rect 8306 -29081 8316 -29071
rect 8236 -29091 8316 -29081
rect 8556 -29081 8566 -29071
rect 8626 -29081 8636 -29021
rect 8556 -29091 8636 -29081
rect 8236 -29361 8296 -29091
rect 8376 -29151 8406 -29131
rect 8356 -29191 8406 -29151
rect 8466 -29151 8496 -29131
rect 8466 -29191 8516 -29151
rect 8356 -29261 8516 -29191
rect 8356 -29301 8406 -29261
rect 8376 -29321 8406 -29301
rect 8466 -29301 8516 -29261
rect 8466 -29321 8496 -29301
rect 8576 -29351 8636 -29091
rect 8566 -29361 8636 -29351
rect 8236 -29371 8316 -29361
rect 8236 -29431 8246 -29371
rect 8306 -29381 8316 -29371
rect 8556 -29371 8636 -29361
rect 8556 -29381 8566 -29371
rect 8306 -29431 8566 -29381
rect 8626 -29431 8636 -29371
rect 8236 -29441 8636 -29431
rect 8692 -29021 9092 -29011
rect 8692 -29081 8702 -29021
rect 8762 -29071 9022 -29021
rect 8762 -29081 8772 -29071
rect 8692 -29091 8772 -29081
rect 9012 -29081 9022 -29071
rect 9082 -29081 9092 -29021
rect 9012 -29091 9092 -29081
rect 8692 -29361 8752 -29091
rect 8832 -29151 8862 -29131
rect 8812 -29191 8862 -29151
rect 8922 -29151 8952 -29131
rect 8922 -29191 8972 -29151
rect 8812 -29261 8972 -29191
rect 8812 -29301 8862 -29261
rect 8832 -29321 8862 -29301
rect 8922 -29301 8972 -29261
rect 8922 -29321 8952 -29301
rect 9032 -29351 9092 -29091
rect 9022 -29361 9092 -29351
rect 8692 -29371 8772 -29361
rect 8692 -29431 8702 -29371
rect 8762 -29381 8772 -29371
rect 9012 -29371 9092 -29361
rect 9012 -29381 9022 -29371
rect 8762 -29431 9022 -29381
rect 9082 -29431 9092 -29371
rect 8692 -29441 9092 -29431
rect 9150 -29021 9550 -29011
rect 9150 -29081 9160 -29021
rect 9220 -29071 9480 -29021
rect 9220 -29081 9230 -29071
rect 9150 -29091 9230 -29081
rect 9470 -29081 9480 -29071
rect 9540 -29081 9550 -29021
rect 9470 -29091 9550 -29081
rect 9150 -29361 9210 -29091
rect 9290 -29151 9320 -29131
rect 9270 -29191 9320 -29151
rect 9380 -29151 9410 -29131
rect 9380 -29191 9430 -29151
rect 9270 -29261 9430 -29191
rect 9270 -29301 9320 -29261
rect 9290 -29321 9320 -29301
rect 9380 -29301 9430 -29261
rect 9380 -29321 9410 -29301
rect 9490 -29351 9550 -29091
rect 9480 -29361 9550 -29351
rect 9150 -29371 9230 -29361
rect 9150 -29431 9160 -29371
rect 9220 -29381 9230 -29371
rect 9470 -29371 9550 -29361
rect 9470 -29381 9480 -29371
rect 9220 -29431 9480 -29381
rect 9540 -29431 9550 -29371
rect 9150 -29441 9550 -29431
rect 9606 -29021 10006 -29011
rect 9606 -29081 9616 -29021
rect 9676 -29071 9936 -29021
rect 9676 -29081 9686 -29071
rect 9606 -29091 9686 -29081
rect 9926 -29081 9936 -29071
rect 9996 -29081 10006 -29021
rect 9926 -29091 10006 -29081
rect 9606 -29361 9666 -29091
rect 9746 -29151 9776 -29131
rect 9726 -29191 9776 -29151
rect 9836 -29151 9866 -29131
rect 9836 -29191 9886 -29151
rect 9726 -29261 9886 -29191
rect 9726 -29301 9776 -29261
rect 9746 -29321 9776 -29301
rect 9836 -29301 9886 -29261
rect 9836 -29321 9866 -29301
rect 9946 -29351 10006 -29091
rect 9936 -29361 10006 -29351
rect 9606 -29371 9686 -29361
rect 9606 -29431 9616 -29371
rect 9676 -29381 9686 -29371
rect 9926 -29371 10006 -29361
rect 9926 -29381 9936 -29371
rect 9676 -29431 9936 -29381
rect 9996 -29431 10006 -29371
rect 9606 -29441 10006 -29431
rect 10062 -29021 10462 -29011
rect 10062 -29081 10072 -29021
rect 10132 -29071 10392 -29021
rect 10132 -29081 10142 -29071
rect 10062 -29091 10142 -29081
rect 10382 -29081 10392 -29071
rect 10452 -29081 10462 -29021
rect 10382 -29091 10462 -29081
rect 10062 -29361 10122 -29091
rect 10202 -29151 10232 -29131
rect 10182 -29191 10232 -29151
rect 10292 -29151 10322 -29131
rect 10292 -29191 10342 -29151
rect 10182 -29261 10342 -29191
rect 10182 -29301 10232 -29261
rect 10202 -29321 10232 -29301
rect 10292 -29301 10342 -29261
rect 10292 -29321 10322 -29301
rect 10402 -29351 10462 -29091
rect 10392 -29361 10462 -29351
rect 10062 -29371 10142 -29361
rect 10062 -29431 10072 -29371
rect 10132 -29381 10142 -29371
rect 10382 -29371 10462 -29361
rect 10382 -29381 10392 -29371
rect 10132 -29431 10392 -29381
rect 10452 -29431 10462 -29371
rect 10062 -29441 10462 -29431
rect 10520 -29021 10920 -29011
rect 10520 -29081 10530 -29021
rect 10590 -29071 10850 -29021
rect 10590 -29081 10600 -29071
rect 10520 -29091 10600 -29081
rect 10840 -29081 10850 -29071
rect 10910 -29081 10920 -29021
rect 10840 -29091 10920 -29081
rect 10520 -29361 10580 -29091
rect 10660 -29151 10690 -29131
rect 10640 -29191 10690 -29151
rect 10750 -29151 10780 -29131
rect 10750 -29191 10800 -29151
rect 10640 -29261 10800 -29191
rect 10640 -29301 10690 -29261
rect 10660 -29321 10690 -29301
rect 10750 -29301 10800 -29261
rect 10750 -29321 10780 -29301
rect 10860 -29351 10920 -29091
rect 10850 -29361 10920 -29351
rect 10520 -29371 10600 -29361
rect 10520 -29431 10530 -29371
rect 10590 -29381 10600 -29371
rect 10840 -29371 10920 -29361
rect 10840 -29381 10850 -29371
rect 10590 -29431 10850 -29381
rect 10910 -29431 10920 -29371
rect 10520 -29441 10920 -29431
rect 10976 -29021 11376 -29011
rect 10976 -29081 10986 -29021
rect 11046 -29071 11306 -29021
rect 11046 -29081 11056 -29071
rect 10976 -29091 11056 -29081
rect 11296 -29081 11306 -29071
rect 11366 -29081 11376 -29021
rect 11296 -29091 11376 -29081
rect 10976 -29361 11036 -29091
rect 11116 -29151 11146 -29131
rect 11096 -29191 11146 -29151
rect 11206 -29151 11236 -29131
rect 11206 -29191 11256 -29151
rect 11096 -29261 11256 -29191
rect 11096 -29301 11146 -29261
rect 11116 -29321 11146 -29301
rect 11206 -29301 11256 -29261
rect 11206 -29321 11236 -29301
rect 11316 -29351 11376 -29091
rect 11306 -29361 11376 -29351
rect 10976 -29371 11056 -29361
rect 10976 -29431 10986 -29371
rect 11046 -29381 11056 -29371
rect 11296 -29371 11376 -29361
rect 11296 -29381 11306 -29371
rect 11046 -29431 11306 -29381
rect 11366 -29431 11376 -29371
rect 10976 -29441 11376 -29431
rect 11432 -29021 11832 -29011
rect 11432 -29081 11442 -29021
rect 11502 -29071 11762 -29021
rect 11502 -29081 11512 -29071
rect 11432 -29091 11512 -29081
rect 11752 -29081 11762 -29071
rect 11822 -29081 11832 -29021
rect 11752 -29091 11832 -29081
rect 11432 -29361 11492 -29091
rect 11572 -29151 11602 -29131
rect 11552 -29191 11602 -29151
rect 11662 -29151 11692 -29131
rect 11662 -29191 11712 -29151
rect 11552 -29261 11712 -29191
rect 11552 -29301 11602 -29261
rect 11572 -29321 11602 -29301
rect 11662 -29301 11712 -29261
rect 11662 -29321 11692 -29301
rect 11772 -29351 11832 -29091
rect 11762 -29361 11832 -29351
rect 11432 -29371 11512 -29361
rect 11432 -29431 11442 -29371
rect 11502 -29381 11512 -29371
rect 11752 -29371 11832 -29361
rect 11752 -29381 11762 -29371
rect 11502 -29431 11762 -29381
rect 11822 -29431 11832 -29371
rect 11432 -29441 11832 -29431
rect 11890 -29021 12290 -29011
rect 11890 -29081 11900 -29021
rect 11960 -29071 12220 -29021
rect 11960 -29081 11970 -29071
rect 11890 -29091 11970 -29081
rect 12210 -29081 12220 -29071
rect 12280 -29081 12290 -29021
rect 12210 -29091 12290 -29081
rect 11890 -29361 11950 -29091
rect 12030 -29151 12060 -29131
rect 12010 -29191 12060 -29151
rect 12120 -29151 12150 -29131
rect 12120 -29191 12170 -29151
rect 12010 -29261 12170 -29191
rect 12010 -29301 12060 -29261
rect 12030 -29321 12060 -29301
rect 12120 -29301 12170 -29261
rect 12120 -29321 12150 -29301
rect 12230 -29351 12290 -29091
rect 12220 -29361 12290 -29351
rect 11890 -29371 11970 -29361
rect 11890 -29431 11900 -29371
rect 11960 -29381 11970 -29371
rect 12210 -29371 12290 -29361
rect 12210 -29381 12220 -29371
rect 11960 -29431 12220 -29381
rect 12280 -29431 12290 -29371
rect 11890 -29441 12290 -29431
rect 12346 -29021 12746 -29011
rect 12346 -29081 12356 -29021
rect 12416 -29071 12676 -29021
rect 12416 -29081 12426 -29071
rect 12346 -29091 12426 -29081
rect 12666 -29081 12676 -29071
rect 12736 -29081 12746 -29021
rect 12666 -29091 12746 -29081
rect 12346 -29361 12406 -29091
rect 12486 -29151 12516 -29131
rect 12466 -29191 12516 -29151
rect 12576 -29151 12606 -29131
rect 12576 -29191 12626 -29151
rect 12466 -29261 12626 -29191
rect 12466 -29301 12516 -29261
rect 12486 -29321 12516 -29301
rect 12576 -29301 12626 -29261
rect 12576 -29321 12606 -29301
rect 12686 -29351 12746 -29091
rect 12676 -29361 12746 -29351
rect 12346 -29371 12426 -29361
rect 12346 -29431 12356 -29371
rect 12416 -29381 12426 -29371
rect 12666 -29371 12746 -29361
rect 12666 -29381 12676 -29371
rect 12416 -29431 12676 -29381
rect 12736 -29431 12746 -29371
rect 12346 -29441 12746 -29431
rect 12802 -29021 13202 -29011
rect 12802 -29081 12812 -29021
rect 12872 -29071 13132 -29021
rect 12872 -29081 12882 -29071
rect 12802 -29091 12882 -29081
rect 13122 -29081 13132 -29071
rect 13192 -29081 13202 -29021
rect 13122 -29091 13202 -29081
rect 12802 -29361 12862 -29091
rect 12942 -29151 12972 -29131
rect 12922 -29191 12972 -29151
rect 13032 -29151 13062 -29131
rect 13032 -29191 13082 -29151
rect 12922 -29261 13082 -29191
rect 12922 -29301 12972 -29261
rect 12942 -29321 12972 -29301
rect 13032 -29301 13082 -29261
rect 13032 -29321 13062 -29301
rect 13142 -29351 13202 -29091
rect 13132 -29361 13202 -29351
rect 12802 -29371 12882 -29361
rect 12802 -29431 12812 -29371
rect 12872 -29381 12882 -29371
rect 13122 -29371 13202 -29361
rect 13122 -29381 13132 -29371
rect 12872 -29431 13132 -29381
rect 13192 -29431 13202 -29371
rect 12802 -29441 13202 -29431
rect 13260 -29021 13660 -29011
rect 13260 -29081 13270 -29021
rect 13330 -29071 13590 -29021
rect 13330 -29081 13340 -29071
rect 13260 -29091 13340 -29081
rect 13580 -29081 13590 -29071
rect 13650 -29081 13660 -29021
rect 13580 -29091 13660 -29081
rect 13260 -29361 13320 -29091
rect 13400 -29151 13430 -29131
rect 13380 -29191 13430 -29151
rect 13490 -29151 13520 -29131
rect 13490 -29191 13540 -29151
rect 13380 -29261 13540 -29191
rect 13380 -29301 13430 -29261
rect 13400 -29321 13430 -29301
rect 13490 -29301 13540 -29261
rect 13490 -29321 13520 -29301
rect 13600 -29351 13660 -29091
rect 13590 -29361 13660 -29351
rect 13260 -29371 13340 -29361
rect 13260 -29431 13270 -29371
rect 13330 -29381 13340 -29371
rect 13580 -29371 13660 -29361
rect 13580 -29381 13590 -29371
rect 13330 -29431 13590 -29381
rect 13650 -29431 13660 -29371
rect 13260 -29441 13660 -29431
rect 13716 -29021 14116 -29011
rect 13716 -29081 13726 -29021
rect 13786 -29071 14046 -29021
rect 13786 -29081 13796 -29071
rect 13716 -29091 13796 -29081
rect 14036 -29081 14046 -29071
rect 14106 -29081 14116 -29021
rect 14036 -29091 14116 -29081
rect 13716 -29361 13776 -29091
rect 13856 -29151 13886 -29131
rect 13836 -29191 13886 -29151
rect 13946 -29151 13976 -29131
rect 13946 -29191 13996 -29151
rect 13836 -29261 13996 -29191
rect 13836 -29301 13886 -29261
rect 13856 -29321 13886 -29301
rect 13946 -29301 13996 -29261
rect 13946 -29321 13976 -29301
rect 14056 -29351 14116 -29091
rect 14046 -29361 14116 -29351
rect 13716 -29371 13796 -29361
rect 13716 -29431 13726 -29371
rect 13786 -29381 13796 -29371
rect 14036 -29371 14116 -29361
rect 14036 -29381 14046 -29371
rect 13786 -29431 14046 -29381
rect 14106 -29431 14116 -29371
rect 13716 -29441 14116 -29431
rect 14172 -29021 14572 -29011
rect 14172 -29081 14182 -29021
rect 14242 -29071 14502 -29021
rect 14242 -29081 14252 -29071
rect 14172 -29091 14252 -29081
rect 14492 -29081 14502 -29071
rect 14562 -29081 14572 -29021
rect 14492 -29091 14572 -29081
rect 14172 -29361 14232 -29091
rect 14312 -29151 14342 -29131
rect 14292 -29191 14342 -29151
rect 14402 -29151 14432 -29131
rect 14402 -29191 14452 -29151
rect 14292 -29261 14452 -29191
rect 14292 -29301 14342 -29261
rect 14312 -29321 14342 -29301
rect 14402 -29301 14452 -29261
rect 14402 -29321 14432 -29301
rect 14512 -29351 14572 -29091
rect 14502 -29361 14572 -29351
rect 14172 -29371 14252 -29361
rect 14172 -29431 14182 -29371
rect 14242 -29381 14252 -29371
rect 14492 -29371 14572 -29361
rect 14492 -29381 14502 -29371
rect 14242 -29431 14502 -29381
rect 14562 -29431 14572 -29371
rect 14172 -29441 14572 -29431
rect 14630 -29021 15030 -29011
rect 14630 -29081 14640 -29021
rect 14700 -29071 14960 -29021
rect 14700 -29081 14710 -29071
rect 14630 -29091 14710 -29081
rect 14950 -29081 14960 -29071
rect 15020 -29081 15030 -29021
rect 14950 -29091 15030 -29081
rect 14630 -29361 14690 -29091
rect 14770 -29151 14800 -29131
rect 14750 -29191 14800 -29151
rect 14860 -29151 14890 -29131
rect 14860 -29191 14910 -29151
rect 14750 -29261 14910 -29191
rect 14750 -29301 14800 -29261
rect 14770 -29321 14800 -29301
rect 14860 -29301 14910 -29261
rect 14860 -29321 14890 -29301
rect 14970 -29351 15030 -29091
rect 14960 -29361 15030 -29351
rect 14630 -29371 14710 -29361
rect 14630 -29431 14640 -29371
rect 14700 -29381 14710 -29371
rect 14950 -29371 15030 -29361
rect 14950 -29381 14960 -29371
rect 14700 -29431 14960 -29381
rect 15020 -29431 15030 -29371
rect 14630 -29441 15030 -29431
rect 15086 -29021 15486 -29011
rect 15086 -29081 15096 -29021
rect 15156 -29071 15416 -29021
rect 15156 -29081 15166 -29071
rect 15086 -29091 15166 -29081
rect 15406 -29081 15416 -29071
rect 15476 -29081 15486 -29021
rect 15406 -29091 15486 -29081
rect 15086 -29361 15146 -29091
rect 15226 -29151 15256 -29131
rect 15206 -29191 15256 -29151
rect 15316 -29151 15346 -29131
rect 15316 -29191 15366 -29151
rect 15206 -29261 15366 -29191
rect 15206 -29301 15256 -29261
rect 15226 -29321 15256 -29301
rect 15316 -29301 15366 -29261
rect 15316 -29321 15346 -29301
rect 15426 -29351 15486 -29091
rect 15416 -29361 15486 -29351
rect 15086 -29371 15166 -29361
rect 15086 -29431 15096 -29371
rect 15156 -29381 15166 -29371
rect 15406 -29371 15486 -29361
rect 15406 -29381 15416 -29371
rect 15156 -29431 15416 -29381
rect 15476 -29431 15486 -29371
rect 15086 -29441 15486 -29431
rect 0 -29513 400 -29503
rect 0 -29573 10 -29513
rect 70 -29563 330 -29513
rect 70 -29573 80 -29563
rect 0 -29583 80 -29573
rect 320 -29573 330 -29563
rect 390 -29573 400 -29513
rect 320 -29583 400 -29573
rect 0 -29853 60 -29583
rect 140 -29643 170 -29623
rect 120 -29683 170 -29643
rect 230 -29643 260 -29623
rect 230 -29683 280 -29643
rect 120 -29753 280 -29683
rect 120 -29793 170 -29753
rect 140 -29813 170 -29793
rect 230 -29793 280 -29753
rect 230 -29813 260 -29793
rect 340 -29843 400 -29583
rect 330 -29853 400 -29843
rect 0 -29863 80 -29853
rect 0 -29923 10 -29863
rect 70 -29873 80 -29863
rect 320 -29863 400 -29853
rect 320 -29873 330 -29863
rect 70 -29923 330 -29873
rect 390 -29923 400 -29863
rect 0 -29933 400 -29923
rect 456 -29513 856 -29503
rect 456 -29573 466 -29513
rect 526 -29563 786 -29513
rect 526 -29573 536 -29563
rect 456 -29583 536 -29573
rect 776 -29573 786 -29563
rect 846 -29573 856 -29513
rect 776 -29583 856 -29573
rect 456 -29853 516 -29583
rect 596 -29643 626 -29623
rect 576 -29683 626 -29643
rect 686 -29643 716 -29623
rect 686 -29683 736 -29643
rect 576 -29753 736 -29683
rect 576 -29793 626 -29753
rect 596 -29813 626 -29793
rect 686 -29793 736 -29753
rect 686 -29813 716 -29793
rect 796 -29843 856 -29583
rect 786 -29853 856 -29843
rect 456 -29863 536 -29853
rect 456 -29923 466 -29863
rect 526 -29873 536 -29863
rect 776 -29863 856 -29853
rect 776 -29873 786 -29863
rect 526 -29923 786 -29873
rect 846 -29923 856 -29863
rect 456 -29933 856 -29923
rect 912 -29513 1312 -29503
rect 912 -29573 922 -29513
rect 982 -29563 1242 -29513
rect 982 -29573 992 -29563
rect 912 -29583 992 -29573
rect 1232 -29573 1242 -29563
rect 1302 -29573 1312 -29513
rect 1232 -29583 1312 -29573
rect 912 -29853 972 -29583
rect 1052 -29643 1082 -29623
rect 1032 -29683 1082 -29643
rect 1142 -29643 1172 -29623
rect 1142 -29683 1192 -29643
rect 1032 -29753 1192 -29683
rect 1032 -29793 1082 -29753
rect 1052 -29813 1082 -29793
rect 1142 -29793 1192 -29753
rect 1142 -29813 1172 -29793
rect 1252 -29843 1312 -29583
rect 1242 -29853 1312 -29843
rect 912 -29863 992 -29853
rect 912 -29923 922 -29863
rect 982 -29873 992 -29863
rect 1232 -29863 1312 -29853
rect 1232 -29873 1242 -29863
rect 982 -29923 1242 -29873
rect 1302 -29923 1312 -29863
rect 912 -29933 1312 -29923
rect 1370 -29513 1770 -29503
rect 1370 -29573 1380 -29513
rect 1440 -29563 1700 -29513
rect 1440 -29573 1450 -29563
rect 1370 -29583 1450 -29573
rect 1690 -29573 1700 -29563
rect 1760 -29573 1770 -29513
rect 1690 -29583 1770 -29573
rect 1370 -29853 1430 -29583
rect 1510 -29643 1540 -29623
rect 1490 -29683 1540 -29643
rect 1600 -29643 1630 -29623
rect 1600 -29683 1650 -29643
rect 1490 -29753 1650 -29683
rect 1490 -29793 1540 -29753
rect 1510 -29813 1540 -29793
rect 1600 -29793 1650 -29753
rect 1600 -29813 1630 -29793
rect 1710 -29843 1770 -29583
rect 1700 -29853 1770 -29843
rect 1370 -29863 1450 -29853
rect 1370 -29923 1380 -29863
rect 1440 -29873 1450 -29863
rect 1690 -29863 1770 -29853
rect 1690 -29873 1700 -29863
rect 1440 -29923 1700 -29873
rect 1760 -29923 1770 -29863
rect 1370 -29933 1770 -29923
rect 1826 -29513 2226 -29503
rect 1826 -29573 1836 -29513
rect 1896 -29563 2156 -29513
rect 1896 -29573 1906 -29563
rect 1826 -29583 1906 -29573
rect 2146 -29573 2156 -29563
rect 2216 -29573 2226 -29513
rect 2146 -29583 2226 -29573
rect 1826 -29853 1886 -29583
rect 1966 -29643 1996 -29623
rect 1946 -29683 1996 -29643
rect 2056 -29643 2086 -29623
rect 2056 -29683 2106 -29643
rect 1946 -29753 2106 -29683
rect 1946 -29793 1996 -29753
rect 1966 -29813 1996 -29793
rect 2056 -29793 2106 -29753
rect 2056 -29813 2086 -29793
rect 2166 -29843 2226 -29583
rect 2156 -29853 2226 -29843
rect 1826 -29863 1906 -29853
rect 1826 -29923 1836 -29863
rect 1896 -29873 1906 -29863
rect 2146 -29863 2226 -29853
rect 2146 -29873 2156 -29863
rect 1896 -29923 2156 -29873
rect 2216 -29923 2226 -29863
rect 1826 -29933 2226 -29923
rect 2282 -29513 2682 -29503
rect 2282 -29573 2292 -29513
rect 2352 -29563 2612 -29513
rect 2352 -29573 2362 -29563
rect 2282 -29583 2362 -29573
rect 2602 -29573 2612 -29563
rect 2672 -29573 2682 -29513
rect 2602 -29583 2682 -29573
rect 2282 -29853 2342 -29583
rect 2422 -29643 2452 -29623
rect 2402 -29683 2452 -29643
rect 2512 -29643 2542 -29623
rect 2512 -29683 2562 -29643
rect 2402 -29753 2562 -29683
rect 2402 -29793 2452 -29753
rect 2422 -29813 2452 -29793
rect 2512 -29793 2562 -29753
rect 2512 -29813 2542 -29793
rect 2622 -29843 2682 -29583
rect 2612 -29853 2682 -29843
rect 2282 -29863 2362 -29853
rect 2282 -29923 2292 -29863
rect 2352 -29873 2362 -29863
rect 2602 -29863 2682 -29853
rect 2602 -29873 2612 -29863
rect 2352 -29923 2612 -29873
rect 2672 -29923 2682 -29863
rect 2282 -29933 2682 -29923
rect 2740 -29513 3140 -29503
rect 2740 -29573 2750 -29513
rect 2810 -29563 3070 -29513
rect 2810 -29573 2820 -29563
rect 2740 -29583 2820 -29573
rect 3060 -29573 3070 -29563
rect 3130 -29573 3140 -29513
rect 3060 -29583 3140 -29573
rect 2740 -29853 2800 -29583
rect 2880 -29643 2910 -29623
rect 2860 -29683 2910 -29643
rect 2970 -29643 3000 -29623
rect 2970 -29683 3020 -29643
rect 2860 -29753 3020 -29683
rect 2860 -29793 2910 -29753
rect 2880 -29813 2910 -29793
rect 2970 -29793 3020 -29753
rect 2970 -29813 3000 -29793
rect 3080 -29843 3140 -29583
rect 3070 -29853 3140 -29843
rect 2740 -29863 2820 -29853
rect 2740 -29923 2750 -29863
rect 2810 -29873 2820 -29863
rect 3060 -29863 3140 -29853
rect 3060 -29873 3070 -29863
rect 2810 -29923 3070 -29873
rect 3130 -29923 3140 -29863
rect 2740 -29933 3140 -29923
rect 3196 -29513 3596 -29503
rect 3196 -29573 3206 -29513
rect 3266 -29563 3526 -29513
rect 3266 -29573 3276 -29563
rect 3196 -29583 3276 -29573
rect 3516 -29573 3526 -29563
rect 3586 -29573 3596 -29513
rect 3516 -29583 3596 -29573
rect 3196 -29853 3256 -29583
rect 3336 -29643 3366 -29623
rect 3316 -29683 3366 -29643
rect 3426 -29643 3456 -29623
rect 3426 -29683 3476 -29643
rect 3316 -29753 3476 -29683
rect 3316 -29793 3366 -29753
rect 3336 -29813 3366 -29793
rect 3426 -29793 3476 -29753
rect 3426 -29813 3456 -29793
rect 3536 -29843 3596 -29583
rect 3526 -29853 3596 -29843
rect 3196 -29863 3276 -29853
rect 3196 -29923 3206 -29863
rect 3266 -29873 3276 -29863
rect 3516 -29863 3596 -29853
rect 3516 -29873 3526 -29863
rect 3266 -29923 3526 -29873
rect 3586 -29923 3596 -29863
rect 3196 -29933 3596 -29923
rect 3652 -29513 4052 -29503
rect 3652 -29573 3662 -29513
rect 3722 -29563 3982 -29513
rect 3722 -29573 3732 -29563
rect 3652 -29583 3732 -29573
rect 3972 -29573 3982 -29563
rect 4042 -29573 4052 -29513
rect 3972 -29583 4052 -29573
rect 3652 -29853 3712 -29583
rect 3792 -29643 3822 -29623
rect 3772 -29683 3822 -29643
rect 3882 -29643 3912 -29623
rect 3882 -29683 3932 -29643
rect 3772 -29753 3932 -29683
rect 3772 -29793 3822 -29753
rect 3792 -29813 3822 -29793
rect 3882 -29793 3932 -29753
rect 3882 -29813 3912 -29793
rect 3992 -29843 4052 -29583
rect 3982 -29853 4052 -29843
rect 3652 -29863 3732 -29853
rect 3652 -29923 3662 -29863
rect 3722 -29873 3732 -29863
rect 3972 -29863 4052 -29853
rect 3972 -29873 3982 -29863
rect 3722 -29923 3982 -29873
rect 4042 -29923 4052 -29863
rect 3652 -29933 4052 -29923
rect 4110 -29513 4510 -29503
rect 4110 -29573 4120 -29513
rect 4180 -29563 4440 -29513
rect 4180 -29573 4190 -29563
rect 4110 -29583 4190 -29573
rect 4430 -29573 4440 -29563
rect 4500 -29573 4510 -29513
rect 4430 -29583 4510 -29573
rect 4110 -29853 4170 -29583
rect 4250 -29643 4280 -29623
rect 4230 -29683 4280 -29643
rect 4340 -29643 4370 -29623
rect 4340 -29683 4390 -29643
rect 4230 -29753 4390 -29683
rect 4230 -29793 4280 -29753
rect 4250 -29813 4280 -29793
rect 4340 -29793 4390 -29753
rect 4340 -29813 4370 -29793
rect 4450 -29843 4510 -29583
rect 4440 -29853 4510 -29843
rect 4110 -29863 4190 -29853
rect 4110 -29923 4120 -29863
rect 4180 -29873 4190 -29863
rect 4430 -29863 4510 -29853
rect 4430 -29873 4440 -29863
rect 4180 -29923 4440 -29873
rect 4500 -29923 4510 -29863
rect 4110 -29933 4510 -29923
rect 4566 -29513 4966 -29503
rect 4566 -29573 4576 -29513
rect 4636 -29563 4896 -29513
rect 4636 -29573 4646 -29563
rect 4566 -29583 4646 -29573
rect 4886 -29573 4896 -29563
rect 4956 -29573 4966 -29513
rect 4886 -29583 4966 -29573
rect 4566 -29853 4626 -29583
rect 4706 -29643 4736 -29623
rect 4686 -29683 4736 -29643
rect 4796 -29643 4826 -29623
rect 4796 -29683 4846 -29643
rect 4686 -29753 4846 -29683
rect 4686 -29793 4736 -29753
rect 4706 -29813 4736 -29793
rect 4796 -29793 4846 -29753
rect 4796 -29813 4826 -29793
rect 4906 -29843 4966 -29583
rect 4896 -29853 4966 -29843
rect 4566 -29863 4646 -29853
rect 4566 -29923 4576 -29863
rect 4636 -29873 4646 -29863
rect 4886 -29863 4966 -29853
rect 4886 -29873 4896 -29863
rect 4636 -29923 4896 -29873
rect 4956 -29923 4966 -29863
rect 4566 -29933 4966 -29923
rect 5022 -29513 5422 -29503
rect 5022 -29573 5032 -29513
rect 5092 -29563 5352 -29513
rect 5092 -29573 5102 -29563
rect 5022 -29583 5102 -29573
rect 5342 -29573 5352 -29563
rect 5412 -29573 5422 -29513
rect 5342 -29583 5422 -29573
rect 5022 -29853 5082 -29583
rect 5162 -29643 5192 -29623
rect 5142 -29683 5192 -29643
rect 5252 -29643 5282 -29623
rect 5252 -29683 5302 -29643
rect 5142 -29753 5302 -29683
rect 5142 -29793 5192 -29753
rect 5162 -29813 5192 -29793
rect 5252 -29793 5302 -29753
rect 5252 -29813 5282 -29793
rect 5362 -29843 5422 -29583
rect 5352 -29853 5422 -29843
rect 5022 -29863 5102 -29853
rect 5022 -29923 5032 -29863
rect 5092 -29873 5102 -29863
rect 5342 -29863 5422 -29853
rect 5342 -29873 5352 -29863
rect 5092 -29923 5352 -29873
rect 5412 -29923 5422 -29863
rect 5022 -29933 5422 -29923
rect 5480 -29513 5880 -29503
rect 5480 -29573 5490 -29513
rect 5550 -29563 5810 -29513
rect 5550 -29573 5560 -29563
rect 5480 -29583 5560 -29573
rect 5800 -29573 5810 -29563
rect 5870 -29573 5880 -29513
rect 5800 -29583 5880 -29573
rect 5480 -29853 5540 -29583
rect 5620 -29643 5650 -29623
rect 5600 -29683 5650 -29643
rect 5710 -29643 5740 -29623
rect 5710 -29683 5760 -29643
rect 5600 -29753 5760 -29683
rect 5600 -29793 5650 -29753
rect 5620 -29813 5650 -29793
rect 5710 -29793 5760 -29753
rect 5710 -29813 5740 -29793
rect 5820 -29843 5880 -29583
rect 5810 -29853 5880 -29843
rect 5480 -29863 5560 -29853
rect 5480 -29923 5490 -29863
rect 5550 -29873 5560 -29863
rect 5800 -29863 5880 -29853
rect 5800 -29873 5810 -29863
rect 5550 -29923 5810 -29873
rect 5870 -29923 5880 -29863
rect 5480 -29933 5880 -29923
rect 5936 -29513 6336 -29503
rect 5936 -29573 5946 -29513
rect 6006 -29563 6266 -29513
rect 6006 -29573 6016 -29563
rect 5936 -29583 6016 -29573
rect 6256 -29573 6266 -29563
rect 6326 -29573 6336 -29513
rect 6256 -29583 6336 -29573
rect 5936 -29853 5996 -29583
rect 6076 -29643 6106 -29623
rect 6056 -29683 6106 -29643
rect 6166 -29643 6196 -29623
rect 6166 -29683 6216 -29643
rect 6056 -29753 6216 -29683
rect 6056 -29793 6106 -29753
rect 6076 -29813 6106 -29793
rect 6166 -29793 6216 -29753
rect 6166 -29813 6196 -29793
rect 6276 -29843 6336 -29583
rect 6266 -29853 6336 -29843
rect 5936 -29863 6016 -29853
rect 5936 -29923 5946 -29863
rect 6006 -29873 6016 -29863
rect 6256 -29863 6336 -29853
rect 6256 -29873 6266 -29863
rect 6006 -29923 6266 -29873
rect 6326 -29923 6336 -29863
rect 5936 -29933 6336 -29923
rect 6392 -29513 6792 -29503
rect 6392 -29573 6402 -29513
rect 6462 -29563 6722 -29513
rect 6462 -29573 6472 -29563
rect 6392 -29583 6472 -29573
rect 6712 -29573 6722 -29563
rect 6782 -29573 6792 -29513
rect 6712 -29583 6792 -29573
rect 6392 -29853 6452 -29583
rect 6532 -29643 6562 -29623
rect 6512 -29683 6562 -29643
rect 6622 -29643 6652 -29623
rect 6622 -29683 6672 -29643
rect 6512 -29753 6672 -29683
rect 6512 -29793 6562 -29753
rect 6532 -29813 6562 -29793
rect 6622 -29793 6672 -29753
rect 6622 -29813 6652 -29793
rect 6732 -29843 6792 -29583
rect 6722 -29853 6792 -29843
rect 6392 -29863 6472 -29853
rect 6392 -29923 6402 -29863
rect 6462 -29873 6472 -29863
rect 6712 -29863 6792 -29853
rect 6712 -29873 6722 -29863
rect 6462 -29923 6722 -29873
rect 6782 -29923 6792 -29863
rect 6392 -29933 6792 -29923
rect 6850 -29513 7250 -29503
rect 6850 -29573 6860 -29513
rect 6920 -29563 7180 -29513
rect 6920 -29573 6930 -29563
rect 6850 -29583 6930 -29573
rect 7170 -29573 7180 -29563
rect 7240 -29573 7250 -29513
rect 7170 -29583 7250 -29573
rect 6850 -29853 6910 -29583
rect 6990 -29643 7020 -29623
rect 6970 -29683 7020 -29643
rect 7080 -29643 7110 -29623
rect 7080 -29683 7130 -29643
rect 6970 -29753 7130 -29683
rect 6970 -29793 7020 -29753
rect 6990 -29813 7020 -29793
rect 7080 -29793 7130 -29753
rect 7080 -29813 7110 -29793
rect 7190 -29843 7250 -29583
rect 7180 -29853 7250 -29843
rect 6850 -29863 6930 -29853
rect 6850 -29923 6860 -29863
rect 6920 -29873 6930 -29863
rect 7170 -29863 7250 -29853
rect 7170 -29873 7180 -29863
rect 6920 -29923 7180 -29873
rect 7240 -29923 7250 -29863
rect 6850 -29933 7250 -29923
rect 7306 -29513 7706 -29503
rect 7306 -29573 7316 -29513
rect 7376 -29563 7636 -29513
rect 7376 -29573 7386 -29563
rect 7306 -29583 7386 -29573
rect 7626 -29573 7636 -29563
rect 7696 -29573 7706 -29513
rect 7626 -29583 7706 -29573
rect 7306 -29853 7366 -29583
rect 7446 -29643 7476 -29623
rect 7426 -29683 7476 -29643
rect 7536 -29643 7566 -29623
rect 7536 -29683 7586 -29643
rect 7426 -29753 7586 -29683
rect 7426 -29793 7476 -29753
rect 7446 -29813 7476 -29793
rect 7536 -29793 7586 -29753
rect 7536 -29813 7566 -29793
rect 7646 -29843 7706 -29583
rect 7636 -29853 7706 -29843
rect 7306 -29863 7386 -29853
rect 7306 -29923 7316 -29863
rect 7376 -29873 7386 -29863
rect 7626 -29863 7706 -29853
rect 7626 -29873 7636 -29863
rect 7376 -29923 7636 -29873
rect 7696 -29923 7706 -29863
rect 7306 -29933 7706 -29923
rect 7762 -29513 8162 -29503
rect 7762 -29573 7772 -29513
rect 7832 -29563 8092 -29513
rect 7832 -29573 7842 -29563
rect 7762 -29583 7842 -29573
rect 8082 -29573 8092 -29563
rect 8152 -29573 8162 -29513
rect 8082 -29583 8162 -29573
rect 7762 -29853 7822 -29583
rect 7902 -29643 7932 -29623
rect 7882 -29683 7932 -29643
rect 7992 -29643 8022 -29623
rect 7992 -29683 8042 -29643
rect 7882 -29753 8042 -29683
rect 7882 -29793 7932 -29753
rect 7902 -29813 7932 -29793
rect 7992 -29793 8042 -29753
rect 7992 -29813 8022 -29793
rect 8102 -29843 8162 -29583
rect 8092 -29853 8162 -29843
rect 7762 -29863 7842 -29853
rect 7762 -29923 7772 -29863
rect 7832 -29873 7842 -29863
rect 8082 -29863 8162 -29853
rect 8082 -29873 8092 -29863
rect 7832 -29923 8092 -29873
rect 8152 -29923 8162 -29863
rect 7762 -29933 8162 -29923
rect 8236 -29513 8636 -29503
rect 8236 -29573 8246 -29513
rect 8306 -29563 8566 -29513
rect 8306 -29573 8316 -29563
rect 8236 -29583 8316 -29573
rect 8556 -29573 8566 -29563
rect 8626 -29573 8636 -29513
rect 8556 -29583 8636 -29573
rect 8236 -29853 8296 -29583
rect 8376 -29643 8406 -29623
rect 8356 -29683 8406 -29643
rect 8466 -29643 8496 -29623
rect 8466 -29683 8516 -29643
rect 8356 -29753 8516 -29683
rect 8356 -29793 8406 -29753
rect 8376 -29813 8406 -29793
rect 8466 -29793 8516 -29753
rect 8466 -29813 8496 -29793
rect 8576 -29843 8636 -29583
rect 8566 -29853 8636 -29843
rect 8236 -29863 8316 -29853
rect 8236 -29923 8246 -29863
rect 8306 -29873 8316 -29863
rect 8556 -29863 8636 -29853
rect 8556 -29873 8566 -29863
rect 8306 -29923 8566 -29873
rect 8626 -29923 8636 -29863
rect 8236 -29933 8636 -29923
rect 8692 -29513 9092 -29503
rect 8692 -29573 8702 -29513
rect 8762 -29563 9022 -29513
rect 8762 -29573 8772 -29563
rect 8692 -29583 8772 -29573
rect 9012 -29573 9022 -29563
rect 9082 -29573 9092 -29513
rect 9012 -29583 9092 -29573
rect 8692 -29853 8752 -29583
rect 8832 -29643 8862 -29623
rect 8812 -29683 8862 -29643
rect 8922 -29643 8952 -29623
rect 8922 -29683 8972 -29643
rect 8812 -29753 8972 -29683
rect 8812 -29793 8862 -29753
rect 8832 -29813 8862 -29793
rect 8922 -29793 8972 -29753
rect 8922 -29813 8952 -29793
rect 9032 -29843 9092 -29583
rect 9022 -29853 9092 -29843
rect 8692 -29863 8772 -29853
rect 8692 -29923 8702 -29863
rect 8762 -29873 8772 -29863
rect 9012 -29863 9092 -29853
rect 9012 -29873 9022 -29863
rect 8762 -29923 9022 -29873
rect 9082 -29923 9092 -29863
rect 8692 -29933 9092 -29923
rect 9150 -29513 9550 -29503
rect 9150 -29573 9160 -29513
rect 9220 -29563 9480 -29513
rect 9220 -29573 9230 -29563
rect 9150 -29583 9230 -29573
rect 9470 -29573 9480 -29563
rect 9540 -29573 9550 -29513
rect 9470 -29583 9550 -29573
rect 9150 -29853 9210 -29583
rect 9290 -29643 9320 -29623
rect 9270 -29683 9320 -29643
rect 9380 -29643 9410 -29623
rect 9380 -29683 9430 -29643
rect 9270 -29753 9430 -29683
rect 9270 -29793 9320 -29753
rect 9290 -29813 9320 -29793
rect 9380 -29793 9430 -29753
rect 9380 -29813 9410 -29793
rect 9490 -29843 9550 -29583
rect 9480 -29853 9550 -29843
rect 9150 -29863 9230 -29853
rect 9150 -29923 9160 -29863
rect 9220 -29873 9230 -29863
rect 9470 -29863 9550 -29853
rect 9470 -29873 9480 -29863
rect 9220 -29923 9480 -29873
rect 9540 -29923 9550 -29863
rect 9150 -29933 9550 -29923
rect 9606 -29513 10006 -29503
rect 9606 -29573 9616 -29513
rect 9676 -29563 9936 -29513
rect 9676 -29573 9686 -29563
rect 9606 -29583 9686 -29573
rect 9926 -29573 9936 -29563
rect 9996 -29573 10006 -29513
rect 9926 -29583 10006 -29573
rect 9606 -29853 9666 -29583
rect 9746 -29643 9776 -29623
rect 9726 -29683 9776 -29643
rect 9836 -29643 9866 -29623
rect 9836 -29683 9886 -29643
rect 9726 -29753 9886 -29683
rect 9726 -29793 9776 -29753
rect 9746 -29813 9776 -29793
rect 9836 -29793 9886 -29753
rect 9836 -29813 9866 -29793
rect 9946 -29843 10006 -29583
rect 9936 -29853 10006 -29843
rect 9606 -29863 9686 -29853
rect 9606 -29923 9616 -29863
rect 9676 -29873 9686 -29863
rect 9926 -29863 10006 -29853
rect 9926 -29873 9936 -29863
rect 9676 -29923 9936 -29873
rect 9996 -29923 10006 -29863
rect 9606 -29933 10006 -29923
rect 10062 -29513 10462 -29503
rect 10062 -29573 10072 -29513
rect 10132 -29563 10392 -29513
rect 10132 -29573 10142 -29563
rect 10062 -29583 10142 -29573
rect 10382 -29573 10392 -29563
rect 10452 -29573 10462 -29513
rect 10382 -29583 10462 -29573
rect 10062 -29853 10122 -29583
rect 10202 -29643 10232 -29623
rect 10182 -29683 10232 -29643
rect 10292 -29643 10322 -29623
rect 10292 -29683 10342 -29643
rect 10182 -29753 10342 -29683
rect 10182 -29793 10232 -29753
rect 10202 -29813 10232 -29793
rect 10292 -29793 10342 -29753
rect 10292 -29813 10322 -29793
rect 10402 -29843 10462 -29583
rect 10392 -29853 10462 -29843
rect 10062 -29863 10142 -29853
rect 10062 -29923 10072 -29863
rect 10132 -29873 10142 -29863
rect 10382 -29863 10462 -29853
rect 10382 -29873 10392 -29863
rect 10132 -29923 10392 -29873
rect 10452 -29923 10462 -29863
rect 10062 -29933 10462 -29923
rect 10520 -29513 10920 -29503
rect 10520 -29573 10530 -29513
rect 10590 -29563 10850 -29513
rect 10590 -29573 10600 -29563
rect 10520 -29583 10600 -29573
rect 10840 -29573 10850 -29563
rect 10910 -29573 10920 -29513
rect 10840 -29583 10920 -29573
rect 10520 -29853 10580 -29583
rect 10660 -29643 10690 -29623
rect 10640 -29683 10690 -29643
rect 10750 -29643 10780 -29623
rect 10750 -29683 10800 -29643
rect 10640 -29753 10800 -29683
rect 10640 -29793 10690 -29753
rect 10660 -29813 10690 -29793
rect 10750 -29793 10800 -29753
rect 10750 -29813 10780 -29793
rect 10860 -29843 10920 -29583
rect 10850 -29853 10920 -29843
rect 10520 -29863 10600 -29853
rect 10520 -29923 10530 -29863
rect 10590 -29873 10600 -29863
rect 10840 -29863 10920 -29853
rect 10840 -29873 10850 -29863
rect 10590 -29923 10850 -29873
rect 10910 -29923 10920 -29863
rect 10520 -29933 10920 -29923
rect 10976 -29513 11376 -29503
rect 10976 -29573 10986 -29513
rect 11046 -29563 11306 -29513
rect 11046 -29573 11056 -29563
rect 10976 -29583 11056 -29573
rect 11296 -29573 11306 -29563
rect 11366 -29573 11376 -29513
rect 11296 -29583 11376 -29573
rect 10976 -29853 11036 -29583
rect 11116 -29643 11146 -29623
rect 11096 -29683 11146 -29643
rect 11206 -29643 11236 -29623
rect 11206 -29683 11256 -29643
rect 11096 -29753 11256 -29683
rect 11096 -29793 11146 -29753
rect 11116 -29813 11146 -29793
rect 11206 -29793 11256 -29753
rect 11206 -29813 11236 -29793
rect 11316 -29843 11376 -29583
rect 11306 -29853 11376 -29843
rect 10976 -29863 11056 -29853
rect 10976 -29923 10986 -29863
rect 11046 -29873 11056 -29863
rect 11296 -29863 11376 -29853
rect 11296 -29873 11306 -29863
rect 11046 -29923 11306 -29873
rect 11366 -29923 11376 -29863
rect 10976 -29933 11376 -29923
rect 11432 -29513 11832 -29503
rect 11432 -29573 11442 -29513
rect 11502 -29563 11762 -29513
rect 11502 -29573 11512 -29563
rect 11432 -29583 11512 -29573
rect 11752 -29573 11762 -29563
rect 11822 -29573 11832 -29513
rect 11752 -29583 11832 -29573
rect 11432 -29853 11492 -29583
rect 11572 -29643 11602 -29623
rect 11552 -29683 11602 -29643
rect 11662 -29643 11692 -29623
rect 11662 -29683 11712 -29643
rect 11552 -29753 11712 -29683
rect 11552 -29793 11602 -29753
rect 11572 -29813 11602 -29793
rect 11662 -29793 11712 -29753
rect 11662 -29813 11692 -29793
rect 11772 -29843 11832 -29583
rect 11762 -29853 11832 -29843
rect 11432 -29863 11512 -29853
rect 11432 -29923 11442 -29863
rect 11502 -29873 11512 -29863
rect 11752 -29863 11832 -29853
rect 11752 -29873 11762 -29863
rect 11502 -29923 11762 -29873
rect 11822 -29923 11832 -29863
rect 11432 -29933 11832 -29923
rect 11890 -29513 12290 -29503
rect 11890 -29573 11900 -29513
rect 11960 -29563 12220 -29513
rect 11960 -29573 11970 -29563
rect 11890 -29583 11970 -29573
rect 12210 -29573 12220 -29563
rect 12280 -29573 12290 -29513
rect 12210 -29583 12290 -29573
rect 11890 -29853 11950 -29583
rect 12030 -29643 12060 -29623
rect 12010 -29683 12060 -29643
rect 12120 -29643 12150 -29623
rect 12120 -29683 12170 -29643
rect 12010 -29753 12170 -29683
rect 12010 -29793 12060 -29753
rect 12030 -29813 12060 -29793
rect 12120 -29793 12170 -29753
rect 12120 -29813 12150 -29793
rect 12230 -29843 12290 -29583
rect 12220 -29853 12290 -29843
rect 11890 -29863 11970 -29853
rect 11890 -29923 11900 -29863
rect 11960 -29873 11970 -29863
rect 12210 -29863 12290 -29853
rect 12210 -29873 12220 -29863
rect 11960 -29923 12220 -29873
rect 12280 -29923 12290 -29863
rect 11890 -29933 12290 -29923
rect 12346 -29513 12746 -29503
rect 12346 -29573 12356 -29513
rect 12416 -29563 12676 -29513
rect 12416 -29573 12426 -29563
rect 12346 -29583 12426 -29573
rect 12666 -29573 12676 -29563
rect 12736 -29573 12746 -29513
rect 12666 -29583 12746 -29573
rect 12346 -29853 12406 -29583
rect 12486 -29643 12516 -29623
rect 12466 -29683 12516 -29643
rect 12576 -29643 12606 -29623
rect 12576 -29683 12626 -29643
rect 12466 -29753 12626 -29683
rect 12466 -29793 12516 -29753
rect 12486 -29813 12516 -29793
rect 12576 -29793 12626 -29753
rect 12576 -29813 12606 -29793
rect 12686 -29843 12746 -29583
rect 12676 -29853 12746 -29843
rect 12346 -29863 12426 -29853
rect 12346 -29923 12356 -29863
rect 12416 -29873 12426 -29863
rect 12666 -29863 12746 -29853
rect 12666 -29873 12676 -29863
rect 12416 -29923 12676 -29873
rect 12736 -29923 12746 -29863
rect 12346 -29933 12746 -29923
rect 12802 -29513 13202 -29503
rect 12802 -29573 12812 -29513
rect 12872 -29563 13132 -29513
rect 12872 -29573 12882 -29563
rect 12802 -29583 12882 -29573
rect 13122 -29573 13132 -29563
rect 13192 -29573 13202 -29513
rect 13122 -29583 13202 -29573
rect 12802 -29853 12862 -29583
rect 12942 -29643 12972 -29623
rect 12922 -29683 12972 -29643
rect 13032 -29643 13062 -29623
rect 13032 -29683 13082 -29643
rect 12922 -29753 13082 -29683
rect 12922 -29793 12972 -29753
rect 12942 -29813 12972 -29793
rect 13032 -29793 13082 -29753
rect 13032 -29813 13062 -29793
rect 13142 -29843 13202 -29583
rect 13132 -29853 13202 -29843
rect 12802 -29863 12882 -29853
rect 12802 -29923 12812 -29863
rect 12872 -29873 12882 -29863
rect 13122 -29863 13202 -29853
rect 13122 -29873 13132 -29863
rect 12872 -29923 13132 -29873
rect 13192 -29923 13202 -29863
rect 12802 -29933 13202 -29923
rect 13260 -29513 13660 -29503
rect 13260 -29573 13270 -29513
rect 13330 -29563 13590 -29513
rect 13330 -29573 13340 -29563
rect 13260 -29583 13340 -29573
rect 13580 -29573 13590 -29563
rect 13650 -29573 13660 -29513
rect 13580 -29583 13660 -29573
rect 13260 -29853 13320 -29583
rect 13400 -29643 13430 -29623
rect 13380 -29683 13430 -29643
rect 13490 -29643 13520 -29623
rect 13490 -29683 13540 -29643
rect 13380 -29753 13540 -29683
rect 13380 -29793 13430 -29753
rect 13400 -29813 13430 -29793
rect 13490 -29793 13540 -29753
rect 13490 -29813 13520 -29793
rect 13600 -29843 13660 -29583
rect 13590 -29853 13660 -29843
rect 13260 -29863 13340 -29853
rect 13260 -29923 13270 -29863
rect 13330 -29873 13340 -29863
rect 13580 -29863 13660 -29853
rect 13580 -29873 13590 -29863
rect 13330 -29923 13590 -29873
rect 13650 -29923 13660 -29863
rect 13260 -29933 13660 -29923
rect 13716 -29513 14116 -29503
rect 13716 -29573 13726 -29513
rect 13786 -29563 14046 -29513
rect 13786 -29573 13796 -29563
rect 13716 -29583 13796 -29573
rect 14036 -29573 14046 -29563
rect 14106 -29573 14116 -29513
rect 14036 -29583 14116 -29573
rect 13716 -29853 13776 -29583
rect 13856 -29643 13886 -29623
rect 13836 -29683 13886 -29643
rect 13946 -29643 13976 -29623
rect 13946 -29683 13996 -29643
rect 13836 -29753 13996 -29683
rect 13836 -29793 13886 -29753
rect 13856 -29813 13886 -29793
rect 13946 -29793 13996 -29753
rect 13946 -29813 13976 -29793
rect 14056 -29843 14116 -29583
rect 14046 -29853 14116 -29843
rect 13716 -29863 13796 -29853
rect 13716 -29923 13726 -29863
rect 13786 -29873 13796 -29863
rect 14036 -29863 14116 -29853
rect 14036 -29873 14046 -29863
rect 13786 -29923 14046 -29873
rect 14106 -29923 14116 -29863
rect 13716 -29933 14116 -29923
rect 14172 -29513 14572 -29503
rect 14172 -29573 14182 -29513
rect 14242 -29563 14502 -29513
rect 14242 -29573 14252 -29563
rect 14172 -29583 14252 -29573
rect 14492 -29573 14502 -29563
rect 14562 -29573 14572 -29513
rect 14492 -29583 14572 -29573
rect 14172 -29853 14232 -29583
rect 14312 -29643 14342 -29623
rect 14292 -29683 14342 -29643
rect 14402 -29643 14432 -29623
rect 14402 -29683 14452 -29643
rect 14292 -29753 14452 -29683
rect 14292 -29793 14342 -29753
rect 14312 -29813 14342 -29793
rect 14402 -29793 14452 -29753
rect 14402 -29813 14432 -29793
rect 14512 -29843 14572 -29583
rect 14502 -29853 14572 -29843
rect 14172 -29863 14252 -29853
rect 14172 -29923 14182 -29863
rect 14242 -29873 14252 -29863
rect 14492 -29863 14572 -29853
rect 14492 -29873 14502 -29863
rect 14242 -29923 14502 -29873
rect 14562 -29923 14572 -29863
rect 14172 -29933 14572 -29923
rect 14630 -29513 15030 -29503
rect 14630 -29573 14640 -29513
rect 14700 -29563 14960 -29513
rect 14700 -29573 14710 -29563
rect 14630 -29583 14710 -29573
rect 14950 -29573 14960 -29563
rect 15020 -29573 15030 -29513
rect 14950 -29583 15030 -29573
rect 14630 -29853 14690 -29583
rect 14770 -29643 14800 -29623
rect 14750 -29683 14800 -29643
rect 14860 -29643 14890 -29623
rect 14860 -29683 14910 -29643
rect 14750 -29753 14910 -29683
rect 14750 -29793 14800 -29753
rect 14770 -29813 14800 -29793
rect 14860 -29793 14910 -29753
rect 14860 -29813 14890 -29793
rect 14970 -29843 15030 -29583
rect 14960 -29853 15030 -29843
rect 14630 -29863 14710 -29853
rect 14630 -29923 14640 -29863
rect 14700 -29873 14710 -29863
rect 14950 -29863 15030 -29853
rect 14950 -29873 14960 -29863
rect 14700 -29923 14960 -29873
rect 15020 -29923 15030 -29863
rect 14630 -29933 15030 -29923
rect 15086 -29513 15486 -29503
rect 15086 -29573 15096 -29513
rect 15156 -29563 15416 -29513
rect 15156 -29573 15166 -29563
rect 15086 -29583 15166 -29573
rect 15406 -29573 15416 -29563
rect 15476 -29573 15486 -29513
rect 15406 -29583 15486 -29573
rect 15086 -29853 15146 -29583
rect 15226 -29643 15256 -29623
rect 15206 -29683 15256 -29643
rect 15316 -29643 15346 -29623
rect 15316 -29683 15366 -29643
rect 15206 -29753 15366 -29683
rect 15206 -29793 15256 -29753
rect 15226 -29813 15256 -29793
rect 15316 -29793 15366 -29753
rect 15316 -29813 15346 -29793
rect 15426 -29843 15486 -29583
rect 15416 -29853 15486 -29843
rect 15086 -29863 15166 -29853
rect 15086 -29923 15096 -29863
rect 15156 -29873 15166 -29863
rect 15406 -29863 15486 -29853
rect 15406 -29873 15416 -29863
rect 15156 -29923 15416 -29873
rect 15476 -29923 15486 -29863
rect 15086 -29933 15486 -29923
rect 0 -30015 400 -30005
rect 0 -30075 10 -30015
rect 70 -30065 330 -30015
rect 70 -30075 80 -30065
rect 0 -30085 80 -30075
rect 320 -30075 330 -30065
rect 390 -30075 400 -30015
rect 320 -30085 400 -30075
rect 0 -30355 60 -30085
rect 140 -30145 170 -30125
rect 120 -30185 170 -30145
rect 230 -30145 260 -30125
rect 230 -30185 280 -30145
rect 120 -30255 280 -30185
rect 120 -30295 170 -30255
rect 140 -30315 170 -30295
rect 230 -30295 280 -30255
rect 230 -30315 260 -30295
rect 340 -30345 400 -30085
rect 330 -30355 400 -30345
rect 0 -30365 80 -30355
rect 0 -30425 10 -30365
rect 70 -30375 80 -30365
rect 320 -30365 400 -30355
rect 320 -30375 330 -30365
rect 70 -30425 330 -30375
rect 390 -30425 400 -30365
rect 0 -30435 400 -30425
rect 456 -30015 856 -30005
rect 456 -30075 466 -30015
rect 526 -30065 786 -30015
rect 526 -30075 536 -30065
rect 456 -30085 536 -30075
rect 776 -30075 786 -30065
rect 846 -30075 856 -30015
rect 776 -30085 856 -30075
rect 456 -30355 516 -30085
rect 596 -30145 626 -30125
rect 576 -30185 626 -30145
rect 686 -30145 716 -30125
rect 686 -30185 736 -30145
rect 576 -30255 736 -30185
rect 576 -30295 626 -30255
rect 596 -30315 626 -30295
rect 686 -30295 736 -30255
rect 686 -30315 716 -30295
rect 796 -30345 856 -30085
rect 786 -30355 856 -30345
rect 456 -30365 536 -30355
rect 456 -30425 466 -30365
rect 526 -30375 536 -30365
rect 776 -30365 856 -30355
rect 776 -30375 786 -30365
rect 526 -30425 786 -30375
rect 846 -30425 856 -30365
rect 456 -30435 856 -30425
rect 912 -30015 1312 -30005
rect 912 -30075 922 -30015
rect 982 -30065 1242 -30015
rect 982 -30075 992 -30065
rect 912 -30085 992 -30075
rect 1232 -30075 1242 -30065
rect 1302 -30075 1312 -30015
rect 1232 -30085 1312 -30075
rect 912 -30355 972 -30085
rect 1052 -30145 1082 -30125
rect 1032 -30185 1082 -30145
rect 1142 -30145 1172 -30125
rect 1142 -30185 1192 -30145
rect 1032 -30255 1192 -30185
rect 1032 -30295 1082 -30255
rect 1052 -30315 1082 -30295
rect 1142 -30295 1192 -30255
rect 1142 -30315 1172 -30295
rect 1252 -30345 1312 -30085
rect 1242 -30355 1312 -30345
rect 912 -30365 992 -30355
rect 912 -30425 922 -30365
rect 982 -30375 992 -30365
rect 1232 -30365 1312 -30355
rect 1232 -30375 1242 -30365
rect 982 -30425 1242 -30375
rect 1302 -30425 1312 -30365
rect 912 -30435 1312 -30425
rect 1370 -30015 1770 -30005
rect 1370 -30075 1380 -30015
rect 1440 -30065 1700 -30015
rect 1440 -30075 1450 -30065
rect 1370 -30085 1450 -30075
rect 1690 -30075 1700 -30065
rect 1760 -30075 1770 -30015
rect 1690 -30085 1770 -30075
rect 1370 -30355 1430 -30085
rect 1510 -30145 1540 -30125
rect 1490 -30185 1540 -30145
rect 1600 -30145 1630 -30125
rect 1600 -30185 1650 -30145
rect 1490 -30255 1650 -30185
rect 1490 -30295 1540 -30255
rect 1510 -30315 1540 -30295
rect 1600 -30295 1650 -30255
rect 1600 -30315 1630 -30295
rect 1710 -30345 1770 -30085
rect 1700 -30355 1770 -30345
rect 1370 -30365 1450 -30355
rect 1370 -30425 1380 -30365
rect 1440 -30375 1450 -30365
rect 1690 -30365 1770 -30355
rect 1690 -30375 1700 -30365
rect 1440 -30425 1700 -30375
rect 1760 -30425 1770 -30365
rect 1370 -30435 1770 -30425
rect 1826 -30015 2226 -30005
rect 1826 -30075 1836 -30015
rect 1896 -30065 2156 -30015
rect 1896 -30075 1906 -30065
rect 1826 -30085 1906 -30075
rect 2146 -30075 2156 -30065
rect 2216 -30075 2226 -30015
rect 2146 -30085 2226 -30075
rect 1826 -30355 1886 -30085
rect 1966 -30145 1996 -30125
rect 1946 -30185 1996 -30145
rect 2056 -30145 2086 -30125
rect 2056 -30185 2106 -30145
rect 1946 -30255 2106 -30185
rect 1946 -30295 1996 -30255
rect 1966 -30315 1996 -30295
rect 2056 -30295 2106 -30255
rect 2056 -30315 2086 -30295
rect 2166 -30345 2226 -30085
rect 2156 -30355 2226 -30345
rect 1826 -30365 1906 -30355
rect 1826 -30425 1836 -30365
rect 1896 -30375 1906 -30365
rect 2146 -30365 2226 -30355
rect 2146 -30375 2156 -30365
rect 1896 -30425 2156 -30375
rect 2216 -30425 2226 -30365
rect 1826 -30435 2226 -30425
rect 2282 -30015 2682 -30005
rect 2282 -30075 2292 -30015
rect 2352 -30065 2612 -30015
rect 2352 -30075 2362 -30065
rect 2282 -30085 2362 -30075
rect 2602 -30075 2612 -30065
rect 2672 -30075 2682 -30015
rect 2602 -30085 2682 -30075
rect 2282 -30355 2342 -30085
rect 2422 -30145 2452 -30125
rect 2402 -30185 2452 -30145
rect 2512 -30145 2542 -30125
rect 2512 -30185 2562 -30145
rect 2402 -30255 2562 -30185
rect 2402 -30295 2452 -30255
rect 2422 -30315 2452 -30295
rect 2512 -30295 2562 -30255
rect 2512 -30315 2542 -30295
rect 2622 -30345 2682 -30085
rect 2612 -30355 2682 -30345
rect 2282 -30365 2362 -30355
rect 2282 -30425 2292 -30365
rect 2352 -30375 2362 -30365
rect 2602 -30365 2682 -30355
rect 2602 -30375 2612 -30365
rect 2352 -30425 2612 -30375
rect 2672 -30425 2682 -30365
rect 2282 -30435 2682 -30425
rect 2740 -30015 3140 -30005
rect 2740 -30075 2750 -30015
rect 2810 -30065 3070 -30015
rect 2810 -30075 2820 -30065
rect 2740 -30085 2820 -30075
rect 3060 -30075 3070 -30065
rect 3130 -30075 3140 -30015
rect 3060 -30085 3140 -30075
rect 2740 -30355 2800 -30085
rect 2880 -30145 2910 -30125
rect 2860 -30185 2910 -30145
rect 2970 -30145 3000 -30125
rect 2970 -30185 3020 -30145
rect 2860 -30255 3020 -30185
rect 2860 -30295 2910 -30255
rect 2880 -30315 2910 -30295
rect 2970 -30295 3020 -30255
rect 2970 -30315 3000 -30295
rect 3080 -30345 3140 -30085
rect 3070 -30355 3140 -30345
rect 2740 -30365 2820 -30355
rect 2740 -30425 2750 -30365
rect 2810 -30375 2820 -30365
rect 3060 -30365 3140 -30355
rect 3060 -30375 3070 -30365
rect 2810 -30425 3070 -30375
rect 3130 -30425 3140 -30365
rect 2740 -30435 3140 -30425
rect 3196 -30015 3596 -30005
rect 3196 -30075 3206 -30015
rect 3266 -30065 3526 -30015
rect 3266 -30075 3276 -30065
rect 3196 -30085 3276 -30075
rect 3516 -30075 3526 -30065
rect 3586 -30075 3596 -30015
rect 3516 -30085 3596 -30075
rect 3196 -30355 3256 -30085
rect 3336 -30145 3366 -30125
rect 3316 -30185 3366 -30145
rect 3426 -30145 3456 -30125
rect 3426 -30185 3476 -30145
rect 3316 -30255 3476 -30185
rect 3316 -30295 3366 -30255
rect 3336 -30315 3366 -30295
rect 3426 -30295 3476 -30255
rect 3426 -30315 3456 -30295
rect 3536 -30345 3596 -30085
rect 3526 -30355 3596 -30345
rect 3196 -30365 3276 -30355
rect 3196 -30425 3206 -30365
rect 3266 -30375 3276 -30365
rect 3516 -30365 3596 -30355
rect 3516 -30375 3526 -30365
rect 3266 -30425 3526 -30375
rect 3586 -30425 3596 -30365
rect 3196 -30435 3596 -30425
rect 3652 -30015 4052 -30005
rect 3652 -30075 3662 -30015
rect 3722 -30065 3982 -30015
rect 3722 -30075 3732 -30065
rect 3652 -30085 3732 -30075
rect 3972 -30075 3982 -30065
rect 4042 -30075 4052 -30015
rect 3972 -30085 4052 -30075
rect 3652 -30355 3712 -30085
rect 3792 -30145 3822 -30125
rect 3772 -30185 3822 -30145
rect 3882 -30145 3912 -30125
rect 3882 -30185 3932 -30145
rect 3772 -30255 3932 -30185
rect 3772 -30295 3822 -30255
rect 3792 -30315 3822 -30295
rect 3882 -30295 3932 -30255
rect 3882 -30315 3912 -30295
rect 3992 -30345 4052 -30085
rect 3982 -30355 4052 -30345
rect 3652 -30365 3732 -30355
rect 3652 -30425 3662 -30365
rect 3722 -30375 3732 -30365
rect 3972 -30365 4052 -30355
rect 3972 -30375 3982 -30365
rect 3722 -30425 3982 -30375
rect 4042 -30425 4052 -30365
rect 3652 -30435 4052 -30425
rect 4110 -30015 4510 -30005
rect 4110 -30075 4120 -30015
rect 4180 -30065 4440 -30015
rect 4180 -30075 4190 -30065
rect 4110 -30085 4190 -30075
rect 4430 -30075 4440 -30065
rect 4500 -30075 4510 -30015
rect 4430 -30085 4510 -30075
rect 4110 -30355 4170 -30085
rect 4250 -30145 4280 -30125
rect 4230 -30185 4280 -30145
rect 4340 -30145 4370 -30125
rect 4340 -30185 4390 -30145
rect 4230 -30255 4390 -30185
rect 4230 -30295 4280 -30255
rect 4250 -30315 4280 -30295
rect 4340 -30295 4390 -30255
rect 4340 -30315 4370 -30295
rect 4450 -30345 4510 -30085
rect 4440 -30355 4510 -30345
rect 4110 -30365 4190 -30355
rect 4110 -30425 4120 -30365
rect 4180 -30375 4190 -30365
rect 4430 -30365 4510 -30355
rect 4430 -30375 4440 -30365
rect 4180 -30425 4440 -30375
rect 4500 -30425 4510 -30365
rect 4110 -30435 4510 -30425
rect 4566 -30015 4966 -30005
rect 4566 -30075 4576 -30015
rect 4636 -30065 4896 -30015
rect 4636 -30075 4646 -30065
rect 4566 -30085 4646 -30075
rect 4886 -30075 4896 -30065
rect 4956 -30075 4966 -30015
rect 4886 -30085 4966 -30075
rect 4566 -30355 4626 -30085
rect 4706 -30145 4736 -30125
rect 4686 -30185 4736 -30145
rect 4796 -30145 4826 -30125
rect 4796 -30185 4846 -30145
rect 4686 -30255 4846 -30185
rect 4686 -30295 4736 -30255
rect 4706 -30315 4736 -30295
rect 4796 -30295 4846 -30255
rect 4796 -30315 4826 -30295
rect 4906 -30345 4966 -30085
rect 4896 -30355 4966 -30345
rect 4566 -30365 4646 -30355
rect 4566 -30425 4576 -30365
rect 4636 -30375 4646 -30365
rect 4886 -30365 4966 -30355
rect 4886 -30375 4896 -30365
rect 4636 -30425 4896 -30375
rect 4956 -30425 4966 -30365
rect 4566 -30435 4966 -30425
rect 5022 -30015 5422 -30005
rect 5022 -30075 5032 -30015
rect 5092 -30065 5352 -30015
rect 5092 -30075 5102 -30065
rect 5022 -30085 5102 -30075
rect 5342 -30075 5352 -30065
rect 5412 -30075 5422 -30015
rect 5342 -30085 5422 -30075
rect 5022 -30355 5082 -30085
rect 5162 -30145 5192 -30125
rect 5142 -30185 5192 -30145
rect 5252 -30145 5282 -30125
rect 5252 -30185 5302 -30145
rect 5142 -30255 5302 -30185
rect 5142 -30295 5192 -30255
rect 5162 -30315 5192 -30295
rect 5252 -30295 5302 -30255
rect 5252 -30315 5282 -30295
rect 5362 -30345 5422 -30085
rect 5352 -30355 5422 -30345
rect 5022 -30365 5102 -30355
rect 5022 -30425 5032 -30365
rect 5092 -30375 5102 -30365
rect 5342 -30365 5422 -30355
rect 5342 -30375 5352 -30365
rect 5092 -30425 5352 -30375
rect 5412 -30425 5422 -30365
rect 5022 -30435 5422 -30425
rect 5480 -30015 5880 -30005
rect 5480 -30075 5490 -30015
rect 5550 -30065 5810 -30015
rect 5550 -30075 5560 -30065
rect 5480 -30085 5560 -30075
rect 5800 -30075 5810 -30065
rect 5870 -30075 5880 -30015
rect 5800 -30085 5880 -30075
rect 5480 -30355 5540 -30085
rect 5620 -30145 5650 -30125
rect 5600 -30185 5650 -30145
rect 5710 -30145 5740 -30125
rect 5710 -30185 5760 -30145
rect 5600 -30255 5760 -30185
rect 5600 -30295 5650 -30255
rect 5620 -30315 5650 -30295
rect 5710 -30295 5760 -30255
rect 5710 -30315 5740 -30295
rect 5820 -30345 5880 -30085
rect 5810 -30355 5880 -30345
rect 5480 -30365 5560 -30355
rect 5480 -30425 5490 -30365
rect 5550 -30375 5560 -30365
rect 5800 -30365 5880 -30355
rect 5800 -30375 5810 -30365
rect 5550 -30425 5810 -30375
rect 5870 -30425 5880 -30365
rect 5480 -30435 5880 -30425
rect 5936 -30015 6336 -30005
rect 5936 -30075 5946 -30015
rect 6006 -30065 6266 -30015
rect 6006 -30075 6016 -30065
rect 5936 -30085 6016 -30075
rect 6256 -30075 6266 -30065
rect 6326 -30075 6336 -30015
rect 6256 -30085 6336 -30075
rect 5936 -30355 5996 -30085
rect 6076 -30145 6106 -30125
rect 6056 -30185 6106 -30145
rect 6166 -30145 6196 -30125
rect 6166 -30185 6216 -30145
rect 6056 -30255 6216 -30185
rect 6056 -30295 6106 -30255
rect 6076 -30315 6106 -30295
rect 6166 -30295 6216 -30255
rect 6166 -30315 6196 -30295
rect 6276 -30345 6336 -30085
rect 6266 -30355 6336 -30345
rect 5936 -30365 6016 -30355
rect 5936 -30425 5946 -30365
rect 6006 -30375 6016 -30365
rect 6256 -30365 6336 -30355
rect 6256 -30375 6266 -30365
rect 6006 -30425 6266 -30375
rect 6326 -30425 6336 -30365
rect 5936 -30435 6336 -30425
rect 6392 -30015 6792 -30005
rect 6392 -30075 6402 -30015
rect 6462 -30065 6722 -30015
rect 6462 -30075 6472 -30065
rect 6392 -30085 6472 -30075
rect 6712 -30075 6722 -30065
rect 6782 -30075 6792 -30015
rect 6712 -30085 6792 -30075
rect 6392 -30355 6452 -30085
rect 6532 -30145 6562 -30125
rect 6512 -30185 6562 -30145
rect 6622 -30145 6652 -30125
rect 6622 -30185 6672 -30145
rect 6512 -30255 6672 -30185
rect 6512 -30295 6562 -30255
rect 6532 -30315 6562 -30295
rect 6622 -30295 6672 -30255
rect 6622 -30315 6652 -30295
rect 6732 -30345 6792 -30085
rect 6722 -30355 6792 -30345
rect 6392 -30365 6472 -30355
rect 6392 -30425 6402 -30365
rect 6462 -30375 6472 -30365
rect 6712 -30365 6792 -30355
rect 6712 -30375 6722 -30365
rect 6462 -30425 6722 -30375
rect 6782 -30425 6792 -30365
rect 6392 -30435 6792 -30425
rect 6850 -30015 7250 -30005
rect 6850 -30075 6860 -30015
rect 6920 -30065 7180 -30015
rect 6920 -30075 6930 -30065
rect 6850 -30085 6930 -30075
rect 7170 -30075 7180 -30065
rect 7240 -30075 7250 -30015
rect 7170 -30085 7250 -30075
rect 6850 -30355 6910 -30085
rect 6990 -30145 7020 -30125
rect 6970 -30185 7020 -30145
rect 7080 -30145 7110 -30125
rect 7080 -30185 7130 -30145
rect 6970 -30255 7130 -30185
rect 6970 -30295 7020 -30255
rect 6990 -30315 7020 -30295
rect 7080 -30295 7130 -30255
rect 7080 -30315 7110 -30295
rect 7190 -30345 7250 -30085
rect 7180 -30355 7250 -30345
rect 6850 -30365 6930 -30355
rect 6850 -30425 6860 -30365
rect 6920 -30375 6930 -30365
rect 7170 -30365 7250 -30355
rect 7170 -30375 7180 -30365
rect 6920 -30425 7180 -30375
rect 7240 -30425 7250 -30365
rect 6850 -30435 7250 -30425
rect 7306 -30015 7706 -30005
rect 7306 -30075 7316 -30015
rect 7376 -30065 7636 -30015
rect 7376 -30075 7386 -30065
rect 7306 -30085 7386 -30075
rect 7626 -30075 7636 -30065
rect 7696 -30075 7706 -30015
rect 7626 -30085 7706 -30075
rect 7306 -30355 7366 -30085
rect 7446 -30145 7476 -30125
rect 7426 -30185 7476 -30145
rect 7536 -30145 7566 -30125
rect 7536 -30185 7586 -30145
rect 7426 -30255 7586 -30185
rect 7426 -30295 7476 -30255
rect 7446 -30315 7476 -30295
rect 7536 -30295 7586 -30255
rect 7536 -30315 7566 -30295
rect 7646 -30345 7706 -30085
rect 7636 -30355 7706 -30345
rect 7306 -30365 7386 -30355
rect 7306 -30425 7316 -30365
rect 7376 -30375 7386 -30365
rect 7626 -30365 7706 -30355
rect 7626 -30375 7636 -30365
rect 7376 -30425 7636 -30375
rect 7696 -30425 7706 -30365
rect 7306 -30435 7706 -30425
rect 7762 -30015 8162 -30005
rect 7762 -30075 7772 -30015
rect 7832 -30065 8092 -30015
rect 7832 -30075 7842 -30065
rect 7762 -30085 7842 -30075
rect 8082 -30075 8092 -30065
rect 8152 -30075 8162 -30015
rect 8082 -30085 8162 -30075
rect 7762 -30355 7822 -30085
rect 7902 -30145 7932 -30125
rect 7882 -30185 7932 -30145
rect 7992 -30145 8022 -30125
rect 7992 -30185 8042 -30145
rect 7882 -30255 8042 -30185
rect 7882 -30295 7932 -30255
rect 7902 -30315 7932 -30295
rect 7992 -30295 8042 -30255
rect 7992 -30315 8022 -30295
rect 8102 -30345 8162 -30085
rect 8092 -30355 8162 -30345
rect 7762 -30365 7842 -30355
rect 7762 -30425 7772 -30365
rect 7832 -30375 7842 -30365
rect 8082 -30365 8162 -30355
rect 8082 -30375 8092 -30365
rect 7832 -30425 8092 -30375
rect 8152 -30425 8162 -30365
rect 7762 -30435 8162 -30425
rect 8236 -30015 8636 -30005
rect 8236 -30075 8246 -30015
rect 8306 -30065 8566 -30015
rect 8306 -30075 8316 -30065
rect 8236 -30085 8316 -30075
rect 8556 -30075 8566 -30065
rect 8626 -30075 8636 -30015
rect 8556 -30085 8636 -30075
rect 8236 -30355 8296 -30085
rect 8376 -30145 8406 -30125
rect 8356 -30185 8406 -30145
rect 8466 -30145 8496 -30125
rect 8466 -30185 8516 -30145
rect 8356 -30255 8516 -30185
rect 8356 -30295 8406 -30255
rect 8376 -30315 8406 -30295
rect 8466 -30295 8516 -30255
rect 8466 -30315 8496 -30295
rect 8576 -30345 8636 -30085
rect 8566 -30355 8636 -30345
rect 8236 -30365 8316 -30355
rect 8236 -30425 8246 -30365
rect 8306 -30375 8316 -30365
rect 8556 -30365 8636 -30355
rect 8556 -30375 8566 -30365
rect 8306 -30425 8566 -30375
rect 8626 -30425 8636 -30365
rect 8236 -30435 8636 -30425
rect 8692 -30015 9092 -30005
rect 8692 -30075 8702 -30015
rect 8762 -30065 9022 -30015
rect 8762 -30075 8772 -30065
rect 8692 -30085 8772 -30075
rect 9012 -30075 9022 -30065
rect 9082 -30075 9092 -30015
rect 9012 -30085 9092 -30075
rect 8692 -30355 8752 -30085
rect 8832 -30145 8862 -30125
rect 8812 -30185 8862 -30145
rect 8922 -30145 8952 -30125
rect 8922 -30185 8972 -30145
rect 8812 -30255 8972 -30185
rect 8812 -30295 8862 -30255
rect 8832 -30315 8862 -30295
rect 8922 -30295 8972 -30255
rect 8922 -30315 8952 -30295
rect 9032 -30345 9092 -30085
rect 9022 -30355 9092 -30345
rect 8692 -30365 8772 -30355
rect 8692 -30425 8702 -30365
rect 8762 -30375 8772 -30365
rect 9012 -30365 9092 -30355
rect 9012 -30375 9022 -30365
rect 8762 -30425 9022 -30375
rect 9082 -30425 9092 -30365
rect 8692 -30435 9092 -30425
rect 9150 -30015 9550 -30005
rect 9150 -30075 9160 -30015
rect 9220 -30065 9480 -30015
rect 9220 -30075 9230 -30065
rect 9150 -30085 9230 -30075
rect 9470 -30075 9480 -30065
rect 9540 -30075 9550 -30015
rect 9470 -30085 9550 -30075
rect 9150 -30355 9210 -30085
rect 9290 -30145 9320 -30125
rect 9270 -30185 9320 -30145
rect 9380 -30145 9410 -30125
rect 9380 -30185 9430 -30145
rect 9270 -30255 9430 -30185
rect 9270 -30295 9320 -30255
rect 9290 -30315 9320 -30295
rect 9380 -30295 9430 -30255
rect 9380 -30315 9410 -30295
rect 9490 -30345 9550 -30085
rect 9480 -30355 9550 -30345
rect 9150 -30365 9230 -30355
rect 9150 -30425 9160 -30365
rect 9220 -30375 9230 -30365
rect 9470 -30365 9550 -30355
rect 9470 -30375 9480 -30365
rect 9220 -30425 9480 -30375
rect 9540 -30425 9550 -30365
rect 9150 -30435 9550 -30425
rect 9606 -30015 10006 -30005
rect 9606 -30075 9616 -30015
rect 9676 -30065 9936 -30015
rect 9676 -30075 9686 -30065
rect 9606 -30085 9686 -30075
rect 9926 -30075 9936 -30065
rect 9996 -30075 10006 -30015
rect 9926 -30085 10006 -30075
rect 9606 -30355 9666 -30085
rect 9746 -30145 9776 -30125
rect 9726 -30185 9776 -30145
rect 9836 -30145 9866 -30125
rect 9836 -30185 9886 -30145
rect 9726 -30255 9886 -30185
rect 9726 -30295 9776 -30255
rect 9746 -30315 9776 -30295
rect 9836 -30295 9886 -30255
rect 9836 -30315 9866 -30295
rect 9946 -30345 10006 -30085
rect 9936 -30355 10006 -30345
rect 9606 -30365 9686 -30355
rect 9606 -30425 9616 -30365
rect 9676 -30375 9686 -30365
rect 9926 -30365 10006 -30355
rect 9926 -30375 9936 -30365
rect 9676 -30425 9936 -30375
rect 9996 -30425 10006 -30365
rect 9606 -30435 10006 -30425
rect 10062 -30015 10462 -30005
rect 10062 -30075 10072 -30015
rect 10132 -30065 10392 -30015
rect 10132 -30075 10142 -30065
rect 10062 -30085 10142 -30075
rect 10382 -30075 10392 -30065
rect 10452 -30075 10462 -30015
rect 10382 -30085 10462 -30075
rect 10062 -30355 10122 -30085
rect 10202 -30145 10232 -30125
rect 10182 -30185 10232 -30145
rect 10292 -30145 10322 -30125
rect 10292 -30185 10342 -30145
rect 10182 -30255 10342 -30185
rect 10182 -30295 10232 -30255
rect 10202 -30315 10232 -30295
rect 10292 -30295 10342 -30255
rect 10292 -30315 10322 -30295
rect 10402 -30345 10462 -30085
rect 10392 -30355 10462 -30345
rect 10062 -30365 10142 -30355
rect 10062 -30425 10072 -30365
rect 10132 -30375 10142 -30365
rect 10382 -30365 10462 -30355
rect 10382 -30375 10392 -30365
rect 10132 -30425 10392 -30375
rect 10452 -30425 10462 -30365
rect 10062 -30435 10462 -30425
rect 10520 -30015 10920 -30005
rect 10520 -30075 10530 -30015
rect 10590 -30065 10850 -30015
rect 10590 -30075 10600 -30065
rect 10520 -30085 10600 -30075
rect 10840 -30075 10850 -30065
rect 10910 -30075 10920 -30015
rect 10840 -30085 10920 -30075
rect 10520 -30355 10580 -30085
rect 10660 -30145 10690 -30125
rect 10640 -30185 10690 -30145
rect 10750 -30145 10780 -30125
rect 10750 -30185 10800 -30145
rect 10640 -30255 10800 -30185
rect 10640 -30295 10690 -30255
rect 10660 -30315 10690 -30295
rect 10750 -30295 10800 -30255
rect 10750 -30315 10780 -30295
rect 10860 -30345 10920 -30085
rect 10850 -30355 10920 -30345
rect 10520 -30365 10600 -30355
rect 10520 -30425 10530 -30365
rect 10590 -30375 10600 -30365
rect 10840 -30365 10920 -30355
rect 10840 -30375 10850 -30365
rect 10590 -30425 10850 -30375
rect 10910 -30425 10920 -30365
rect 10520 -30435 10920 -30425
rect 10976 -30015 11376 -30005
rect 10976 -30075 10986 -30015
rect 11046 -30065 11306 -30015
rect 11046 -30075 11056 -30065
rect 10976 -30085 11056 -30075
rect 11296 -30075 11306 -30065
rect 11366 -30075 11376 -30015
rect 11296 -30085 11376 -30075
rect 10976 -30355 11036 -30085
rect 11116 -30145 11146 -30125
rect 11096 -30185 11146 -30145
rect 11206 -30145 11236 -30125
rect 11206 -30185 11256 -30145
rect 11096 -30255 11256 -30185
rect 11096 -30295 11146 -30255
rect 11116 -30315 11146 -30295
rect 11206 -30295 11256 -30255
rect 11206 -30315 11236 -30295
rect 11316 -30345 11376 -30085
rect 11306 -30355 11376 -30345
rect 10976 -30365 11056 -30355
rect 10976 -30425 10986 -30365
rect 11046 -30375 11056 -30365
rect 11296 -30365 11376 -30355
rect 11296 -30375 11306 -30365
rect 11046 -30425 11306 -30375
rect 11366 -30425 11376 -30365
rect 10976 -30435 11376 -30425
rect 11432 -30015 11832 -30005
rect 11432 -30075 11442 -30015
rect 11502 -30065 11762 -30015
rect 11502 -30075 11512 -30065
rect 11432 -30085 11512 -30075
rect 11752 -30075 11762 -30065
rect 11822 -30075 11832 -30015
rect 11752 -30085 11832 -30075
rect 11432 -30355 11492 -30085
rect 11572 -30145 11602 -30125
rect 11552 -30185 11602 -30145
rect 11662 -30145 11692 -30125
rect 11662 -30185 11712 -30145
rect 11552 -30255 11712 -30185
rect 11552 -30295 11602 -30255
rect 11572 -30315 11602 -30295
rect 11662 -30295 11712 -30255
rect 11662 -30315 11692 -30295
rect 11772 -30345 11832 -30085
rect 11762 -30355 11832 -30345
rect 11432 -30365 11512 -30355
rect 11432 -30425 11442 -30365
rect 11502 -30375 11512 -30365
rect 11752 -30365 11832 -30355
rect 11752 -30375 11762 -30365
rect 11502 -30425 11762 -30375
rect 11822 -30425 11832 -30365
rect 11432 -30435 11832 -30425
rect 11890 -30015 12290 -30005
rect 11890 -30075 11900 -30015
rect 11960 -30065 12220 -30015
rect 11960 -30075 11970 -30065
rect 11890 -30085 11970 -30075
rect 12210 -30075 12220 -30065
rect 12280 -30075 12290 -30015
rect 12210 -30085 12290 -30075
rect 11890 -30355 11950 -30085
rect 12030 -30145 12060 -30125
rect 12010 -30185 12060 -30145
rect 12120 -30145 12150 -30125
rect 12120 -30185 12170 -30145
rect 12010 -30255 12170 -30185
rect 12010 -30295 12060 -30255
rect 12030 -30315 12060 -30295
rect 12120 -30295 12170 -30255
rect 12120 -30315 12150 -30295
rect 12230 -30345 12290 -30085
rect 12220 -30355 12290 -30345
rect 11890 -30365 11970 -30355
rect 11890 -30425 11900 -30365
rect 11960 -30375 11970 -30365
rect 12210 -30365 12290 -30355
rect 12210 -30375 12220 -30365
rect 11960 -30425 12220 -30375
rect 12280 -30425 12290 -30365
rect 11890 -30435 12290 -30425
rect 12346 -30015 12746 -30005
rect 12346 -30075 12356 -30015
rect 12416 -30065 12676 -30015
rect 12416 -30075 12426 -30065
rect 12346 -30085 12426 -30075
rect 12666 -30075 12676 -30065
rect 12736 -30075 12746 -30015
rect 12666 -30085 12746 -30075
rect 12346 -30355 12406 -30085
rect 12486 -30145 12516 -30125
rect 12466 -30185 12516 -30145
rect 12576 -30145 12606 -30125
rect 12576 -30185 12626 -30145
rect 12466 -30255 12626 -30185
rect 12466 -30295 12516 -30255
rect 12486 -30315 12516 -30295
rect 12576 -30295 12626 -30255
rect 12576 -30315 12606 -30295
rect 12686 -30345 12746 -30085
rect 12676 -30355 12746 -30345
rect 12346 -30365 12426 -30355
rect 12346 -30425 12356 -30365
rect 12416 -30375 12426 -30365
rect 12666 -30365 12746 -30355
rect 12666 -30375 12676 -30365
rect 12416 -30425 12676 -30375
rect 12736 -30425 12746 -30365
rect 12346 -30435 12746 -30425
rect 12802 -30015 13202 -30005
rect 12802 -30075 12812 -30015
rect 12872 -30065 13132 -30015
rect 12872 -30075 12882 -30065
rect 12802 -30085 12882 -30075
rect 13122 -30075 13132 -30065
rect 13192 -30075 13202 -30015
rect 13122 -30085 13202 -30075
rect 12802 -30355 12862 -30085
rect 12942 -30145 12972 -30125
rect 12922 -30185 12972 -30145
rect 13032 -30145 13062 -30125
rect 13032 -30185 13082 -30145
rect 12922 -30255 13082 -30185
rect 12922 -30295 12972 -30255
rect 12942 -30315 12972 -30295
rect 13032 -30295 13082 -30255
rect 13032 -30315 13062 -30295
rect 13142 -30345 13202 -30085
rect 13132 -30355 13202 -30345
rect 12802 -30365 12882 -30355
rect 12802 -30425 12812 -30365
rect 12872 -30375 12882 -30365
rect 13122 -30365 13202 -30355
rect 13122 -30375 13132 -30365
rect 12872 -30425 13132 -30375
rect 13192 -30425 13202 -30365
rect 12802 -30435 13202 -30425
rect 13260 -30015 13660 -30005
rect 13260 -30075 13270 -30015
rect 13330 -30065 13590 -30015
rect 13330 -30075 13340 -30065
rect 13260 -30085 13340 -30075
rect 13580 -30075 13590 -30065
rect 13650 -30075 13660 -30015
rect 13580 -30085 13660 -30075
rect 13260 -30355 13320 -30085
rect 13400 -30145 13430 -30125
rect 13380 -30185 13430 -30145
rect 13490 -30145 13520 -30125
rect 13490 -30185 13540 -30145
rect 13380 -30255 13540 -30185
rect 13380 -30295 13430 -30255
rect 13400 -30315 13430 -30295
rect 13490 -30295 13540 -30255
rect 13490 -30315 13520 -30295
rect 13600 -30345 13660 -30085
rect 13590 -30355 13660 -30345
rect 13260 -30365 13340 -30355
rect 13260 -30425 13270 -30365
rect 13330 -30375 13340 -30365
rect 13580 -30365 13660 -30355
rect 13580 -30375 13590 -30365
rect 13330 -30425 13590 -30375
rect 13650 -30425 13660 -30365
rect 13260 -30435 13660 -30425
rect 13716 -30015 14116 -30005
rect 13716 -30075 13726 -30015
rect 13786 -30065 14046 -30015
rect 13786 -30075 13796 -30065
rect 13716 -30085 13796 -30075
rect 14036 -30075 14046 -30065
rect 14106 -30075 14116 -30015
rect 14036 -30085 14116 -30075
rect 13716 -30355 13776 -30085
rect 13856 -30145 13886 -30125
rect 13836 -30185 13886 -30145
rect 13946 -30145 13976 -30125
rect 13946 -30185 13996 -30145
rect 13836 -30255 13996 -30185
rect 13836 -30295 13886 -30255
rect 13856 -30315 13886 -30295
rect 13946 -30295 13996 -30255
rect 13946 -30315 13976 -30295
rect 14056 -30345 14116 -30085
rect 14046 -30355 14116 -30345
rect 13716 -30365 13796 -30355
rect 13716 -30425 13726 -30365
rect 13786 -30375 13796 -30365
rect 14036 -30365 14116 -30355
rect 14036 -30375 14046 -30365
rect 13786 -30425 14046 -30375
rect 14106 -30425 14116 -30365
rect 13716 -30435 14116 -30425
rect 14172 -30015 14572 -30005
rect 14172 -30075 14182 -30015
rect 14242 -30065 14502 -30015
rect 14242 -30075 14252 -30065
rect 14172 -30085 14252 -30075
rect 14492 -30075 14502 -30065
rect 14562 -30075 14572 -30015
rect 14492 -30085 14572 -30075
rect 14172 -30355 14232 -30085
rect 14312 -30145 14342 -30125
rect 14292 -30185 14342 -30145
rect 14402 -30145 14432 -30125
rect 14402 -30185 14452 -30145
rect 14292 -30255 14452 -30185
rect 14292 -30295 14342 -30255
rect 14312 -30315 14342 -30295
rect 14402 -30295 14452 -30255
rect 14402 -30315 14432 -30295
rect 14512 -30345 14572 -30085
rect 14502 -30355 14572 -30345
rect 14172 -30365 14252 -30355
rect 14172 -30425 14182 -30365
rect 14242 -30375 14252 -30365
rect 14492 -30365 14572 -30355
rect 14492 -30375 14502 -30365
rect 14242 -30425 14502 -30375
rect 14562 -30425 14572 -30365
rect 14172 -30435 14572 -30425
rect 14630 -30015 15030 -30005
rect 14630 -30075 14640 -30015
rect 14700 -30065 14960 -30015
rect 14700 -30075 14710 -30065
rect 14630 -30085 14710 -30075
rect 14950 -30075 14960 -30065
rect 15020 -30075 15030 -30015
rect 14950 -30085 15030 -30075
rect 14630 -30355 14690 -30085
rect 14770 -30145 14800 -30125
rect 14750 -30185 14800 -30145
rect 14860 -30145 14890 -30125
rect 14860 -30185 14910 -30145
rect 14750 -30255 14910 -30185
rect 14750 -30295 14800 -30255
rect 14770 -30315 14800 -30295
rect 14860 -30295 14910 -30255
rect 14860 -30315 14890 -30295
rect 14970 -30345 15030 -30085
rect 14960 -30355 15030 -30345
rect 14630 -30365 14710 -30355
rect 14630 -30425 14640 -30365
rect 14700 -30375 14710 -30365
rect 14950 -30365 15030 -30355
rect 14950 -30375 14960 -30365
rect 14700 -30425 14960 -30375
rect 15020 -30425 15030 -30365
rect 14630 -30435 15030 -30425
rect 15086 -30015 15486 -30005
rect 15086 -30075 15096 -30015
rect 15156 -30065 15416 -30015
rect 15156 -30075 15166 -30065
rect 15086 -30085 15166 -30075
rect 15406 -30075 15416 -30065
rect 15476 -30075 15486 -30015
rect 15406 -30085 15486 -30075
rect 15086 -30355 15146 -30085
rect 15226 -30145 15256 -30125
rect 15206 -30185 15256 -30145
rect 15316 -30145 15346 -30125
rect 15316 -30185 15366 -30145
rect 15206 -30255 15366 -30185
rect 15206 -30295 15256 -30255
rect 15226 -30315 15256 -30295
rect 15316 -30295 15366 -30255
rect 15316 -30315 15346 -30295
rect 15426 -30345 15486 -30085
rect 15416 -30355 15486 -30345
rect 15086 -30365 15166 -30355
rect 15086 -30425 15096 -30365
rect 15156 -30375 15166 -30365
rect 15406 -30365 15486 -30355
rect 15406 -30375 15416 -30365
rect 15156 -30425 15416 -30375
rect 15476 -30425 15486 -30365
rect 15086 -30435 15486 -30425
rect 0 -30531 400 -30521
rect 0 -30591 10 -30531
rect 70 -30581 330 -30531
rect 70 -30591 80 -30581
rect 0 -30601 80 -30591
rect 320 -30591 330 -30581
rect 390 -30591 400 -30531
rect 320 -30601 400 -30591
rect 0 -30871 60 -30601
rect 140 -30661 170 -30641
rect 120 -30701 170 -30661
rect 230 -30661 260 -30641
rect 230 -30701 280 -30661
rect 120 -30771 280 -30701
rect 120 -30811 170 -30771
rect 140 -30831 170 -30811
rect 230 -30811 280 -30771
rect 230 -30831 260 -30811
rect 340 -30861 400 -30601
rect 330 -30871 400 -30861
rect 0 -30881 80 -30871
rect 0 -30941 10 -30881
rect 70 -30891 80 -30881
rect 320 -30881 400 -30871
rect 320 -30891 330 -30881
rect 70 -30941 330 -30891
rect 390 -30941 400 -30881
rect 0 -30951 400 -30941
rect 456 -30531 856 -30521
rect 456 -30591 466 -30531
rect 526 -30581 786 -30531
rect 526 -30591 536 -30581
rect 456 -30601 536 -30591
rect 776 -30591 786 -30581
rect 846 -30591 856 -30531
rect 776 -30601 856 -30591
rect 456 -30871 516 -30601
rect 596 -30661 626 -30641
rect 576 -30701 626 -30661
rect 686 -30661 716 -30641
rect 686 -30701 736 -30661
rect 576 -30771 736 -30701
rect 576 -30811 626 -30771
rect 596 -30831 626 -30811
rect 686 -30811 736 -30771
rect 686 -30831 716 -30811
rect 796 -30861 856 -30601
rect 786 -30871 856 -30861
rect 456 -30881 536 -30871
rect 456 -30941 466 -30881
rect 526 -30891 536 -30881
rect 776 -30881 856 -30871
rect 776 -30891 786 -30881
rect 526 -30941 786 -30891
rect 846 -30941 856 -30881
rect 456 -30951 856 -30941
rect 912 -30531 1312 -30521
rect 912 -30591 922 -30531
rect 982 -30581 1242 -30531
rect 982 -30591 992 -30581
rect 912 -30601 992 -30591
rect 1232 -30591 1242 -30581
rect 1302 -30591 1312 -30531
rect 1232 -30601 1312 -30591
rect 912 -30871 972 -30601
rect 1052 -30661 1082 -30641
rect 1032 -30701 1082 -30661
rect 1142 -30661 1172 -30641
rect 1142 -30701 1192 -30661
rect 1032 -30771 1192 -30701
rect 1032 -30811 1082 -30771
rect 1052 -30831 1082 -30811
rect 1142 -30811 1192 -30771
rect 1142 -30831 1172 -30811
rect 1252 -30861 1312 -30601
rect 1242 -30871 1312 -30861
rect 912 -30881 992 -30871
rect 912 -30941 922 -30881
rect 982 -30891 992 -30881
rect 1232 -30881 1312 -30871
rect 1232 -30891 1242 -30881
rect 982 -30941 1242 -30891
rect 1302 -30941 1312 -30881
rect 912 -30951 1312 -30941
rect 1370 -30531 1770 -30521
rect 1370 -30591 1380 -30531
rect 1440 -30581 1700 -30531
rect 1440 -30591 1450 -30581
rect 1370 -30601 1450 -30591
rect 1690 -30591 1700 -30581
rect 1760 -30591 1770 -30531
rect 1690 -30601 1770 -30591
rect 1370 -30871 1430 -30601
rect 1510 -30661 1540 -30641
rect 1490 -30701 1540 -30661
rect 1600 -30661 1630 -30641
rect 1600 -30701 1650 -30661
rect 1490 -30771 1650 -30701
rect 1490 -30811 1540 -30771
rect 1510 -30831 1540 -30811
rect 1600 -30811 1650 -30771
rect 1600 -30831 1630 -30811
rect 1710 -30861 1770 -30601
rect 1700 -30871 1770 -30861
rect 1370 -30881 1450 -30871
rect 1370 -30941 1380 -30881
rect 1440 -30891 1450 -30881
rect 1690 -30881 1770 -30871
rect 1690 -30891 1700 -30881
rect 1440 -30941 1700 -30891
rect 1760 -30941 1770 -30881
rect 1370 -30951 1770 -30941
rect 1826 -30531 2226 -30521
rect 1826 -30591 1836 -30531
rect 1896 -30581 2156 -30531
rect 1896 -30591 1906 -30581
rect 1826 -30601 1906 -30591
rect 2146 -30591 2156 -30581
rect 2216 -30591 2226 -30531
rect 2146 -30601 2226 -30591
rect 1826 -30871 1886 -30601
rect 1966 -30661 1996 -30641
rect 1946 -30701 1996 -30661
rect 2056 -30661 2086 -30641
rect 2056 -30701 2106 -30661
rect 1946 -30771 2106 -30701
rect 1946 -30811 1996 -30771
rect 1966 -30831 1996 -30811
rect 2056 -30811 2106 -30771
rect 2056 -30831 2086 -30811
rect 2166 -30861 2226 -30601
rect 2156 -30871 2226 -30861
rect 1826 -30881 1906 -30871
rect 1826 -30941 1836 -30881
rect 1896 -30891 1906 -30881
rect 2146 -30881 2226 -30871
rect 2146 -30891 2156 -30881
rect 1896 -30941 2156 -30891
rect 2216 -30941 2226 -30881
rect 1826 -30951 2226 -30941
rect 2282 -30531 2682 -30521
rect 2282 -30591 2292 -30531
rect 2352 -30581 2612 -30531
rect 2352 -30591 2362 -30581
rect 2282 -30601 2362 -30591
rect 2602 -30591 2612 -30581
rect 2672 -30591 2682 -30531
rect 2602 -30601 2682 -30591
rect 2282 -30871 2342 -30601
rect 2422 -30661 2452 -30641
rect 2402 -30701 2452 -30661
rect 2512 -30661 2542 -30641
rect 2512 -30701 2562 -30661
rect 2402 -30771 2562 -30701
rect 2402 -30811 2452 -30771
rect 2422 -30831 2452 -30811
rect 2512 -30811 2562 -30771
rect 2512 -30831 2542 -30811
rect 2622 -30861 2682 -30601
rect 2612 -30871 2682 -30861
rect 2282 -30881 2362 -30871
rect 2282 -30941 2292 -30881
rect 2352 -30891 2362 -30881
rect 2602 -30881 2682 -30871
rect 2602 -30891 2612 -30881
rect 2352 -30941 2612 -30891
rect 2672 -30941 2682 -30881
rect 2282 -30951 2682 -30941
rect 2740 -30531 3140 -30521
rect 2740 -30591 2750 -30531
rect 2810 -30581 3070 -30531
rect 2810 -30591 2820 -30581
rect 2740 -30601 2820 -30591
rect 3060 -30591 3070 -30581
rect 3130 -30591 3140 -30531
rect 3060 -30601 3140 -30591
rect 2740 -30871 2800 -30601
rect 2880 -30661 2910 -30641
rect 2860 -30701 2910 -30661
rect 2970 -30661 3000 -30641
rect 2970 -30701 3020 -30661
rect 2860 -30771 3020 -30701
rect 2860 -30811 2910 -30771
rect 2880 -30831 2910 -30811
rect 2970 -30811 3020 -30771
rect 2970 -30831 3000 -30811
rect 3080 -30861 3140 -30601
rect 3070 -30871 3140 -30861
rect 2740 -30881 2820 -30871
rect 2740 -30941 2750 -30881
rect 2810 -30891 2820 -30881
rect 3060 -30881 3140 -30871
rect 3060 -30891 3070 -30881
rect 2810 -30941 3070 -30891
rect 3130 -30941 3140 -30881
rect 2740 -30951 3140 -30941
rect 3196 -30531 3596 -30521
rect 3196 -30591 3206 -30531
rect 3266 -30581 3526 -30531
rect 3266 -30591 3276 -30581
rect 3196 -30601 3276 -30591
rect 3516 -30591 3526 -30581
rect 3586 -30591 3596 -30531
rect 3516 -30601 3596 -30591
rect 3196 -30871 3256 -30601
rect 3336 -30661 3366 -30641
rect 3316 -30701 3366 -30661
rect 3426 -30661 3456 -30641
rect 3426 -30701 3476 -30661
rect 3316 -30771 3476 -30701
rect 3316 -30811 3366 -30771
rect 3336 -30831 3366 -30811
rect 3426 -30811 3476 -30771
rect 3426 -30831 3456 -30811
rect 3536 -30861 3596 -30601
rect 3526 -30871 3596 -30861
rect 3196 -30881 3276 -30871
rect 3196 -30941 3206 -30881
rect 3266 -30891 3276 -30881
rect 3516 -30881 3596 -30871
rect 3516 -30891 3526 -30881
rect 3266 -30941 3526 -30891
rect 3586 -30941 3596 -30881
rect 3196 -30951 3596 -30941
rect 3652 -30531 4052 -30521
rect 3652 -30591 3662 -30531
rect 3722 -30581 3982 -30531
rect 3722 -30591 3732 -30581
rect 3652 -30601 3732 -30591
rect 3972 -30591 3982 -30581
rect 4042 -30591 4052 -30531
rect 3972 -30601 4052 -30591
rect 3652 -30871 3712 -30601
rect 3792 -30661 3822 -30641
rect 3772 -30701 3822 -30661
rect 3882 -30661 3912 -30641
rect 3882 -30701 3932 -30661
rect 3772 -30771 3932 -30701
rect 3772 -30811 3822 -30771
rect 3792 -30831 3822 -30811
rect 3882 -30811 3932 -30771
rect 3882 -30831 3912 -30811
rect 3992 -30861 4052 -30601
rect 3982 -30871 4052 -30861
rect 3652 -30881 3732 -30871
rect 3652 -30941 3662 -30881
rect 3722 -30891 3732 -30881
rect 3972 -30881 4052 -30871
rect 3972 -30891 3982 -30881
rect 3722 -30941 3982 -30891
rect 4042 -30941 4052 -30881
rect 3652 -30951 4052 -30941
rect 4110 -30531 4510 -30521
rect 4110 -30591 4120 -30531
rect 4180 -30581 4440 -30531
rect 4180 -30591 4190 -30581
rect 4110 -30601 4190 -30591
rect 4430 -30591 4440 -30581
rect 4500 -30591 4510 -30531
rect 4430 -30601 4510 -30591
rect 4110 -30871 4170 -30601
rect 4250 -30661 4280 -30641
rect 4230 -30701 4280 -30661
rect 4340 -30661 4370 -30641
rect 4340 -30701 4390 -30661
rect 4230 -30771 4390 -30701
rect 4230 -30811 4280 -30771
rect 4250 -30831 4280 -30811
rect 4340 -30811 4390 -30771
rect 4340 -30831 4370 -30811
rect 4450 -30861 4510 -30601
rect 4440 -30871 4510 -30861
rect 4110 -30881 4190 -30871
rect 4110 -30941 4120 -30881
rect 4180 -30891 4190 -30881
rect 4430 -30881 4510 -30871
rect 4430 -30891 4440 -30881
rect 4180 -30941 4440 -30891
rect 4500 -30941 4510 -30881
rect 4110 -30951 4510 -30941
rect 4566 -30531 4966 -30521
rect 4566 -30591 4576 -30531
rect 4636 -30581 4896 -30531
rect 4636 -30591 4646 -30581
rect 4566 -30601 4646 -30591
rect 4886 -30591 4896 -30581
rect 4956 -30591 4966 -30531
rect 4886 -30601 4966 -30591
rect 4566 -30871 4626 -30601
rect 4706 -30661 4736 -30641
rect 4686 -30701 4736 -30661
rect 4796 -30661 4826 -30641
rect 4796 -30701 4846 -30661
rect 4686 -30771 4846 -30701
rect 4686 -30811 4736 -30771
rect 4706 -30831 4736 -30811
rect 4796 -30811 4846 -30771
rect 4796 -30831 4826 -30811
rect 4906 -30861 4966 -30601
rect 4896 -30871 4966 -30861
rect 4566 -30881 4646 -30871
rect 4566 -30941 4576 -30881
rect 4636 -30891 4646 -30881
rect 4886 -30881 4966 -30871
rect 4886 -30891 4896 -30881
rect 4636 -30941 4896 -30891
rect 4956 -30941 4966 -30881
rect 4566 -30951 4966 -30941
rect 5022 -30531 5422 -30521
rect 5022 -30591 5032 -30531
rect 5092 -30581 5352 -30531
rect 5092 -30591 5102 -30581
rect 5022 -30601 5102 -30591
rect 5342 -30591 5352 -30581
rect 5412 -30591 5422 -30531
rect 5342 -30601 5422 -30591
rect 5022 -30871 5082 -30601
rect 5162 -30661 5192 -30641
rect 5142 -30701 5192 -30661
rect 5252 -30661 5282 -30641
rect 5252 -30701 5302 -30661
rect 5142 -30771 5302 -30701
rect 5142 -30811 5192 -30771
rect 5162 -30831 5192 -30811
rect 5252 -30811 5302 -30771
rect 5252 -30831 5282 -30811
rect 5362 -30861 5422 -30601
rect 5352 -30871 5422 -30861
rect 5022 -30881 5102 -30871
rect 5022 -30941 5032 -30881
rect 5092 -30891 5102 -30881
rect 5342 -30881 5422 -30871
rect 5342 -30891 5352 -30881
rect 5092 -30941 5352 -30891
rect 5412 -30941 5422 -30881
rect 5022 -30951 5422 -30941
rect 5480 -30531 5880 -30521
rect 5480 -30591 5490 -30531
rect 5550 -30581 5810 -30531
rect 5550 -30591 5560 -30581
rect 5480 -30601 5560 -30591
rect 5800 -30591 5810 -30581
rect 5870 -30591 5880 -30531
rect 5800 -30601 5880 -30591
rect 5480 -30871 5540 -30601
rect 5620 -30661 5650 -30641
rect 5600 -30701 5650 -30661
rect 5710 -30661 5740 -30641
rect 5710 -30701 5760 -30661
rect 5600 -30771 5760 -30701
rect 5600 -30811 5650 -30771
rect 5620 -30831 5650 -30811
rect 5710 -30811 5760 -30771
rect 5710 -30831 5740 -30811
rect 5820 -30861 5880 -30601
rect 5810 -30871 5880 -30861
rect 5480 -30881 5560 -30871
rect 5480 -30941 5490 -30881
rect 5550 -30891 5560 -30881
rect 5800 -30881 5880 -30871
rect 5800 -30891 5810 -30881
rect 5550 -30941 5810 -30891
rect 5870 -30941 5880 -30881
rect 5480 -30951 5880 -30941
rect 5936 -30531 6336 -30521
rect 5936 -30591 5946 -30531
rect 6006 -30581 6266 -30531
rect 6006 -30591 6016 -30581
rect 5936 -30601 6016 -30591
rect 6256 -30591 6266 -30581
rect 6326 -30591 6336 -30531
rect 6256 -30601 6336 -30591
rect 5936 -30871 5996 -30601
rect 6076 -30661 6106 -30641
rect 6056 -30701 6106 -30661
rect 6166 -30661 6196 -30641
rect 6166 -30701 6216 -30661
rect 6056 -30771 6216 -30701
rect 6056 -30811 6106 -30771
rect 6076 -30831 6106 -30811
rect 6166 -30811 6216 -30771
rect 6166 -30831 6196 -30811
rect 6276 -30861 6336 -30601
rect 6266 -30871 6336 -30861
rect 5936 -30881 6016 -30871
rect 5936 -30941 5946 -30881
rect 6006 -30891 6016 -30881
rect 6256 -30881 6336 -30871
rect 6256 -30891 6266 -30881
rect 6006 -30941 6266 -30891
rect 6326 -30941 6336 -30881
rect 5936 -30951 6336 -30941
rect 6392 -30531 6792 -30521
rect 6392 -30591 6402 -30531
rect 6462 -30581 6722 -30531
rect 6462 -30591 6472 -30581
rect 6392 -30601 6472 -30591
rect 6712 -30591 6722 -30581
rect 6782 -30591 6792 -30531
rect 6712 -30601 6792 -30591
rect 6392 -30871 6452 -30601
rect 6532 -30661 6562 -30641
rect 6512 -30701 6562 -30661
rect 6622 -30661 6652 -30641
rect 6622 -30701 6672 -30661
rect 6512 -30771 6672 -30701
rect 6512 -30811 6562 -30771
rect 6532 -30831 6562 -30811
rect 6622 -30811 6672 -30771
rect 6622 -30831 6652 -30811
rect 6732 -30861 6792 -30601
rect 6722 -30871 6792 -30861
rect 6392 -30881 6472 -30871
rect 6392 -30941 6402 -30881
rect 6462 -30891 6472 -30881
rect 6712 -30881 6792 -30871
rect 6712 -30891 6722 -30881
rect 6462 -30941 6722 -30891
rect 6782 -30941 6792 -30881
rect 6392 -30951 6792 -30941
rect 6850 -30531 7250 -30521
rect 6850 -30591 6860 -30531
rect 6920 -30581 7180 -30531
rect 6920 -30591 6930 -30581
rect 6850 -30601 6930 -30591
rect 7170 -30591 7180 -30581
rect 7240 -30591 7250 -30531
rect 7170 -30601 7250 -30591
rect 6850 -30871 6910 -30601
rect 6990 -30661 7020 -30641
rect 6970 -30701 7020 -30661
rect 7080 -30661 7110 -30641
rect 7080 -30701 7130 -30661
rect 6970 -30771 7130 -30701
rect 6970 -30811 7020 -30771
rect 6990 -30831 7020 -30811
rect 7080 -30811 7130 -30771
rect 7080 -30831 7110 -30811
rect 7190 -30861 7250 -30601
rect 7180 -30871 7250 -30861
rect 6850 -30881 6930 -30871
rect 6850 -30941 6860 -30881
rect 6920 -30891 6930 -30881
rect 7170 -30881 7250 -30871
rect 7170 -30891 7180 -30881
rect 6920 -30941 7180 -30891
rect 7240 -30941 7250 -30881
rect 6850 -30951 7250 -30941
rect 7306 -30531 7706 -30521
rect 7306 -30591 7316 -30531
rect 7376 -30581 7636 -30531
rect 7376 -30591 7386 -30581
rect 7306 -30601 7386 -30591
rect 7626 -30591 7636 -30581
rect 7696 -30591 7706 -30531
rect 7626 -30601 7706 -30591
rect 7306 -30871 7366 -30601
rect 7446 -30661 7476 -30641
rect 7426 -30701 7476 -30661
rect 7536 -30661 7566 -30641
rect 7536 -30701 7586 -30661
rect 7426 -30771 7586 -30701
rect 7426 -30811 7476 -30771
rect 7446 -30831 7476 -30811
rect 7536 -30811 7586 -30771
rect 7536 -30831 7566 -30811
rect 7646 -30861 7706 -30601
rect 7636 -30871 7706 -30861
rect 7306 -30881 7386 -30871
rect 7306 -30941 7316 -30881
rect 7376 -30891 7386 -30881
rect 7626 -30881 7706 -30871
rect 7626 -30891 7636 -30881
rect 7376 -30941 7636 -30891
rect 7696 -30941 7706 -30881
rect 7306 -30951 7706 -30941
rect 7762 -30531 8162 -30521
rect 7762 -30591 7772 -30531
rect 7832 -30581 8092 -30531
rect 7832 -30591 7842 -30581
rect 7762 -30601 7842 -30591
rect 8082 -30591 8092 -30581
rect 8152 -30591 8162 -30531
rect 8082 -30601 8162 -30591
rect 7762 -30871 7822 -30601
rect 7902 -30661 7932 -30641
rect 7882 -30701 7932 -30661
rect 7992 -30661 8022 -30641
rect 7992 -30701 8042 -30661
rect 7882 -30771 8042 -30701
rect 7882 -30811 7932 -30771
rect 7902 -30831 7932 -30811
rect 7992 -30811 8042 -30771
rect 7992 -30831 8022 -30811
rect 8102 -30861 8162 -30601
rect 8092 -30871 8162 -30861
rect 7762 -30881 7842 -30871
rect 7762 -30941 7772 -30881
rect 7832 -30891 7842 -30881
rect 8082 -30881 8162 -30871
rect 8082 -30891 8092 -30881
rect 7832 -30941 8092 -30891
rect 8152 -30941 8162 -30881
rect 7762 -30951 8162 -30941
rect 8236 -30531 8636 -30521
rect 8236 -30591 8246 -30531
rect 8306 -30581 8566 -30531
rect 8306 -30591 8316 -30581
rect 8236 -30601 8316 -30591
rect 8556 -30591 8566 -30581
rect 8626 -30591 8636 -30531
rect 8556 -30601 8636 -30591
rect 8236 -30871 8296 -30601
rect 8376 -30661 8406 -30641
rect 8356 -30701 8406 -30661
rect 8466 -30661 8496 -30641
rect 8466 -30701 8516 -30661
rect 8356 -30771 8516 -30701
rect 8356 -30811 8406 -30771
rect 8376 -30831 8406 -30811
rect 8466 -30811 8516 -30771
rect 8466 -30831 8496 -30811
rect 8576 -30861 8636 -30601
rect 8566 -30871 8636 -30861
rect 8236 -30881 8316 -30871
rect 8236 -30941 8246 -30881
rect 8306 -30891 8316 -30881
rect 8556 -30881 8636 -30871
rect 8556 -30891 8566 -30881
rect 8306 -30941 8566 -30891
rect 8626 -30941 8636 -30881
rect 8236 -30951 8636 -30941
rect 8692 -30531 9092 -30521
rect 8692 -30591 8702 -30531
rect 8762 -30581 9022 -30531
rect 8762 -30591 8772 -30581
rect 8692 -30601 8772 -30591
rect 9012 -30591 9022 -30581
rect 9082 -30591 9092 -30531
rect 9012 -30601 9092 -30591
rect 8692 -30871 8752 -30601
rect 8832 -30661 8862 -30641
rect 8812 -30701 8862 -30661
rect 8922 -30661 8952 -30641
rect 8922 -30701 8972 -30661
rect 8812 -30771 8972 -30701
rect 8812 -30811 8862 -30771
rect 8832 -30831 8862 -30811
rect 8922 -30811 8972 -30771
rect 8922 -30831 8952 -30811
rect 9032 -30861 9092 -30601
rect 9022 -30871 9092 -30861
rect 8692 -30881 8772 -30871
rect 8692 -30941 8702 -30881
rect 8762 -30891 8772 -30881
rect 9012 -30881 9092 -30871
rect 9012 -30891 9022 -30881
rect 8762 -30941 9022 -30891
rect 9082 -30941 9092 -30881
rect 8692 -30951 9092 -30941
rect 9150 -30531 9550 -30521
rect 9150 -30591 9160 -30531
rect 9220 -30581 9480 -30531
rect 9220 -30591 9230 -30581
rect 9150 -30601 9230 -30591
rect 9470 -30591 9480 -30581
rect 9540 -30591 9550 -30531
rect 9470 -30601 9550 -30591
rect 9150 -30871 9210 -30601
rect 9290 -30661 9320 -30641
rect 9270 -30701 9320 -30661
rect 9380 -30661 9410 -30641
rect 9380 -30701 9430 -30661
rect 9270 -30771 9430 -30701
rect 9270 -30811 9320 -30771
rect 9290 -30831 9320 -30811
rect 9380 -30811 9430 -30771
rect 9380 -30831 9410 -30811
rect 9490 -30861 9550 -30601
rect 9480 -30871 9550 -30861
rect 9150 -30881 9230 -30871
rect 9150 -30941 9160 -30881
rect 9220 -30891 9230 -30881
rect 9470 -30881 9550 -30871
rect 9470 -30891 9480 -30881
rect 9220 -30941 9480 -30891
rect 9540 -30941 9550 -30881
rect 9150 -30951 9550 -30941
rect 9606 -30531 10006 -30521
rect 9606 -30591 9616 -30531
rect 9676 -30581 9936 -30531
rect 9676 -30591 9686 -30581
rect 9606 -30601 9686 -30591
rect 9926 -30591 9936 -30581
rect 9996 -30591 10006 -30531
rect 9926 -30601 10006 -30591
rect 9606 -30871 9666 -30601
rect 9746 -30661 9776 -30641
rect 9726 -30701 9776 -30661
rect 9836 -30661 9866 -30641
rect 9836 -30701 9886 -30661
rect 9726 -30771 9886 -30701
rect 9726 -30811 9776 -30771
rect 9746 -30831 9776 -30811
rect 9836 -30811 9886 -30771
rect 9836 -30831 9866 -30811
rect 9946 -30861 10006 -30601
rect 9936 -30871 10006 -30861
rect 9606 -30881 9686 -30871
rect 9606 -30941 9616 -30881
rect 9676 -30891 9686 -30881
rect 9926 -30881 10006 -30871
rect 9926 -30891 9936 -30881
rect 9676 -30941 9936 -30891
rect 9996 -30941 10006 -30881
rect 9606 -30951 10006 -30941
rect 10062 -30531 10462 -30521
rect 10062 -30591 10072 -30531
rect 10132 -30581 10392 -30531
rect 10132 -30591 10142 -30581
rect 10062 -30601 10142 -30591
rect 10382 -30591 10392 -30581
rect 10452 -30591 10462 -30531
rect 10382 -30601 10462 -30591
rect 10062 -30871 10122 -30601
rect 10202 -30661 10232 -30641
rect 10182 -30701 10232 -30661
rect 10292 -30661 10322 -30641
rect 10292 -30701 10342 -30661
rect 10182 -30771 10342 -30701
rect 10182 -30811 10232 -30771
rect 10202 -30831 10232 -30811
rect 10292 -30811 10342 -30771
rect 10292 -30831 10322 -30811
rect 10402 -30861 10462 -30601
rect 10392 -30871 10462 -30861
rect 10062 -30881 10142 -30871
rect 10062 -30941 10072 -30881
rect 10132 -30891 10142 -30881
rect 10382 -30881 10462 -30871
rect 10382 -30891 10392 -30881
rect 10132 -30941 10392 -30891
rect 10452 -30941 10462 -30881
rect 10062 -30951 10462 -30941
rect 10520 -30531 10920 -30521
rect 10520 -30591 10530 -30531
rect 10590 -30581 10850 -30531
rect 10590 -30591 10600 -30581
rect 10520 -30601 10600 -30591
rect 10840 -30591 10850 -30581
rect 10910 -30591 10920 -30531
rect 10840 -30601 10920 -30591
rect 10520 -30871 10580 -30601
rect 10660 -30661 10690 -30641
rect 10640 -30701 10690 -30661
rect 10750 -30661 10780 -30641
rect 10750 -30701 10800 -30661
rect 10640 -30771 10800 -30701
rect 10640 -30811 10690 -30771
rect 10660 -30831 10690 -30811
rect 10750 -30811 10800 -30771
rect 10750 -30831 10780 -30811
rect 10860 -30861 10920 -30601
rect 10850 -30871 10920 -30861
rect 10520 -30881 10600 -30871
rect 10520 -30941 10530 -30881
rect 10590 -30891 10600 -30881
rect 10840 -30881 10920 -30871
rect 10840 -30891 10850 -30881
rect 10590 -30941 10850 -30891
rect 10910 -30941 10920 -30881
rect 10520 -30951 10920 -30941
rect 10976 -30531 11376 -30521
rect 10976 -30591 10986 -30531
rect 11046 -30581 11306 -30531
rect 11046 -30591 11056 -30581
rect 10976 -30601 11056 -30591
rect 11296 -30591 11306 -30581
rect 11366 -30591 11376 -30531
rect 11296 -30601 11376 -30591
rect 10976 -30871 11036 -30601
rect 11116 -30661 11146 -30641
rect 11096 -30701 11146 -30661
rect 11206 -30661 11236 -30641
rect 11206 -30701 11256 -30661
rect 11096 -30771 11256 -30701
rect 11096 -30811 11146 -30771
rect 11116 -30831 11146 -30811
rect 11206 -30811 11256 -30771
rect 11206 -30831 11236 -30811
rect 11316 -30861 11376 -30601
rect 11306 -30871 11376 -30861
rect 10976 -30881 11056 -30871
rect 10976 -30941 10986 -30881
rect 11046 -30891 11056 -30881
rect 11296 -30881 11376 -30871
rect 11296 -30891 11306 -30881
rect 11046 -30941 11306 -30891
rect 11366 -30941 11376 -30881
rect 10976 -30951 11376 -30941
rect 11432 -30531 11832 -30521
rect 11432 -30591 11442 -30531
rect 11502 -30581 11762 -30531
rect 11502 -30591 11512 -30581
rect 11432 -30601 11512 -30591
rect 11752 -30591 11762 -30581
rect 11822 -30591 11832 -30531
rect 11752 -30601 11832 -30591
rect 11432 -30871 11492 -30601
rect 11572 -30661 11602 -30641
rect 11552 -30701 11602 -30661
rect 11662 -30661 11692 -30641
rect 11662 -30701 11712 -30661
rect 11552 -30771 11712 -30701
rect 11552 -30811 11602 -30771
rect 11572 -30831 11602 -30811
rect 11662 -30811 11712 -30771
rect 11662 -30831 11692 -30811
rect 11772 -30861 11832 -30601
rect 11762 -30871 11832 -30861
rect 11432 -30881 11512 -30871
rect 11432 -30941 11442 -30881
rect 11502 -30891 11512 -30881
rect 11752 -30881 11832 -30871
rect 11752 -30891 11762 -30881
rect 11502 -30941 11762 -30891
rect 11822 -30941 11832 -30881
rect 11432 -30951 11832 -30941
rect 11890 -30531 12290 -30521
rect 11890 -30591 11900 -30531
rect 11960 -30581 12220 -30531
rect 11960 -30591 11970 -30581
rect 11890 -30601 11970 -30591
rect 12210 -30591 12220 -30581
rect 12280 -30591 12290 -30531
rect 12210 -30601 12290 -30591
rect 11890 -30871 11950 -30601
rect 12030 -30661 12060 -30641
rect 12010 -30701 12060 -30661
rect 12120 -30661 12150 -30641
rect 12120 -30701 12170 -30661
rect 12010 -30771 12170 -30701
rect 12010 -30811 12060 -30771
rect 12030 -30831 12060 -30811
rect 12120 -30811 12170 -30771
rect 12120 -30831 12150 -30811
rect 12230 -30861 12290 -30601
rect 12220 -30871 12290 -30861
rect 11890 -30881 11970 -30871
rect 11890 -30941 11900 -30881
rect 11960 -30891 11970 -30881
rect 12210 -30881 12290 -30871
rect 12210 -30891 12220 -30881
rect 11960 -30941 12220 -30891
rect 12280 -30941 12290 -30881
rect 11890 -30951 12290 -30941
rect 12346 -30531 12746 -30521
rect 12346 -30591 12356 -30531
rect 12416 -30581 12676 -30531
rect 12416 -30591 12426 -30581
rect 12346 -30601 12426 -30591
rect 12666 -30591 12676 -30581
rect 12736 -30591 12746 -30531
rect 12666 -30601 12746 -30591
rect 12346 -30871 12406 -30601
rect 12486 -30661 12516 -30641
rect 12466 -30701 12516 -30661
rect 12576 -30661 12606 -30641
rect 12576 -30701 12626 -30661
rect 12466 -30771 12626 -30701
rect 12466 -30811 12516 -30771
rect 12486 -30831 12516 -30811
rect 12576 -30811 12626 -30771
rect 12576 -30831 12606 -30811
rect 12686 -30861 12746 -30601
rect 12676 -30871 12746 -30861
rect 12346 -30881 12426 -30871
rect 12346 -30941 12356 -30881
rect 12416 -30891 12426 -30881
rect 12666 -30881 12746 -30871
rect 12666 -30891 12676 -30881
rect 12416 -30941 12676 -30891
rect 12736 -30941 12746 -30881
rect 12346 -30951 12746 -30941
rect 12802 -30531 13202 -30521
rect 12802 -30591 12812 -30531
rect 12872 -30581 13132 -30531
rect 12872 -30591 12882 -30581
rect 12802 -30601 12882 -30591
rect 13122 -30591 13132 -30581
rect 13192 -30591 13202 -30531
rect 13122 -30601 13202 -30591
rect 12802 -30871 12862 -30601
rect 12942 -30661 12972 -30641
rect 12922 -30701 12972 -30661
rect 13032 -30661 13062 -30641
rect 13032 -30701 13082 -30661
rect 12922 -30771 13082 -30701
rect 12922 -30811 12972 -30771
rect 12942 -30831 12972 -30811
rect 13032 -30811 13082 -30771
rect 13032 -30831 13062 -30811
rect 13142 -30861 13202 -30601
rect 13132 -30871 13202 -30861
rect 12802 -30881 12882 -30871
rect 12802 -30941 12812 -30881
rect 12872 -30891 12882 -30881
rect 13122 -30881 13202 -30871
rect 13122 -30891 13132 -30881
rect 12872 -30941 13132 -30891
rect 13192 -30941 13202 -30881
rect 12802 -30951 13202 -30941
rect 13260 -30531 13660 -30521
rect 13260 -30591 13270 -30531
rect 13330 -30581 13590 -30531
rect 13330 -30591 13340 -30581
rect 13260 -30601 13340 -30591
rect 13580 -30591 13590 -30581
rect 13650 -30591 13660 -30531
rect 13580 -30601 13660 -30591
rect 13260 -30871 13320 -30601
rect 13400 -30661 13430 -30641
rect 13380 -30701 13430 -30661
rect 13490 -30661 13520 -30641
rect 13490 -30701 13540 -30661
rect 13380 -30771 13540 -30701
rect 13380 -30811 13430 -30771
rect 13400 -30831 13430 -30811
rect 13490 -30811 13540 -30771
rect 13490 -30831 13520 -30811
rect 13600 -30861 13660 -30601
rect 13590 -30871 13660 -30861
rect 13260 -30881 13340 -30871
rect 13260 -30941 13270 -30881
rect 13330 -30891 13340 -30881
rect 13580 -30881 13660 -30871
rect 13580 -30891 13590 -30881
rect 13330 -30941 13590 -30891
rect 13650 -30941 13660 -30881
rect 13260 -30951 13660 -30941
rect 13716 -30531 14116 -30521
rect 13716 -30591 13726 -30531
rect 13786 -30581 14046 -30531
rect 13786 -30591 13796 -30581
rect 13716 -30601 13796 -30591
rect 14036 -30591 14046 -30581
rect 14106 -30591 14116 -30531
rect 14036 -30601 14116 -30591
rect 13716 -30871 13776 -30601
rect 13856 -30661 13886 -30641
rect 13836 -30701 13886 -30661
rect 13946 -30661 13976 -30641
rect 13946 -30701 13996 -30661
rect 13836 -30771 13996 -30701
rect 13836 -30811 13886 -30771
rect 13856 -30831 13886 -30811
rect 13946 -30811 13996 -30771
rect 13946 -30831 13976 -30811
rect 14056 -30861 14116 -30601
rect 14046 -30871 14116 -30861
rect 13716 -30881 13796 -30871
rect 13716 -30941 13726 -30881
rect 13786 -30891 13796 -30881
rect 14036 -30881 14116 -30871
rect 14036 -30891 14046 -30881
rect 13786 -30941 14046 -30891
rect 14106 -30941 14116 -30881
rect 13716 -30951 14116 -30941
rect 14172 -30531 14572 -30521
rect 14172 -30591 14182 -30531
rect 14242 -30581 14502 -30531
rect 14242 -30591 14252 -30581
rect 14172 -30601 14252 -30591
rect 14492 -30591 14502 -30581
rect 14562 -30591 14572 -30531
rect 14492 -30601 14572 -30591
rect 14172 -30871 14232 -30601
rect 14312 -30661 14342 -30641
rect 14292 -30701 14342 -30661
rect 14402 -30661 14432 -30641
rect 14402 -30701 14452 -30661
rect 14292 -30771 14452 -30701
rect 14292 -30811 14342 -30771
rect 14312 -30831 14342 -30811
rect 14402 -30811 14452 -30771
rect 14402 -30831 14432 -30811
rect 14512 -30861 14572 -30601
rect 14502 -30871 14572 -30861
rect 14172 -30881 14252 -30871
rect 14172 -30941 14182 -30881
rect 14242 -30891 14252 -30881
rect 14492 -30881 14572 -30871
rect 14492 -30891 14502 -30881
rect 14242 -30941 14502 -30891
rect 14562 -30941 14572 -30881
rect 14172 -30951 14572 -30941
rect 14630 -30531 15030 -30521
rect 14630 -30591 14640 -30531
rect 14700 -30581 14960 -30531
rect 14700 -30591 14710 -30581
rect 14630 -30601 14710 -30591
rect 14950 -30591 14960 -30581
rect 15020 -30591 15030 -30531
rect 14950 -30601 15030 -30591
rect 14630 -30871 14690 -30601
rect 14770 -30661 14800 -30641
rect 14750 -30701 14800 -30661
rect 14860 -30661 14890 -30641
rect 14860 -30701 14910 -30661
rect 14750 -30771 14910 -30701
rect 14750 -30811 14800 -30771
rect 14770 -30831 14800 -30811
rect 14860 -30811 14910 -30771
rect 14860 -30831 14890 -30811
rect 14970 -30861 15030 -30601
rect 14960 -30871 15030 -30861
rect 14630 -30881 14710 -30871
rect 14630 -30941 14640 -30881
rect 14700 -30891 14710 -30881
rect 14950 -30881 15030 -30871
rect 14950 -30891 14960 -30881
rect 14700 -30941 14960 -30891
rect 15020 -30941 15030 -30881
rect 14630 -30951 15030 -30941
rect 15086 -30531 15486 -30521
rect 15086 -30591 15096 -30531
rect 15156 -30581 15416 -30531
rect 15156 -30591 15166 -30581
rect 15086 -30601 15166 -30591
rect 15406 -30591 15416 -30581
rect 15476 -30591 15486 -30531
rect 15406 -30601 15486 -30591
rect 15086 -30871 15146 -30601
rect 15226 -30661 15256 -30641
rect 15206 -30701 15256 -30661
rect 15316 -30661 15346 -30641
rect 15316 -30701 15366 -30661
rect 15206 -30771 15366 -30701
rect 15206 -30811 15256 -30771
rect 15226 -30831 15256 -30811
rect 15316 -30811 15366 -30771
rect 15316 -30831 15346 -30811
rect 15426 -30861 15486 -30601
rect 15416 -30871 15486 -30861
rect 15086 -30881 15166 -30871
rect 15086 -30941 15096 -30881
rect 15156 -30891 15166 -30881
rect 15406 -30881 15486 -30871
rect 15406 -30891 15416 -30881
rect 15156 -30941 15416 -30891
rect 15476 -30941 15486 -30881
rect 15086 -30951 15486 -30941
rect 0 -31023 400 -31013
rect 0 -31083 10 -31023
rect 70 -31073 330 -31023
rect 70 -31083 80 -31073
rect 0 -31093 80 -31083
rect 320 -31083 330 -31073
rect 390 -31083 400 -31023
rect 320 -31093 400 -31083
rect 0 -31363 60 -31093
rect 140 -31153 170 -31133
rect 120 -31193 170 -31153
rect 230 -31153 260 -31133
rect 230 -31193 280 -31153
rect 120 -31263 280 -31193
rect 120 -31303 170 -31263
rect 140 -31323 170 -31303
rect 230 -31303 280 -31263
rect 230 -31323 260 -31303
rect 340 -31353 400 -31093
rect 330 -31363 400 -31353
rect 0 -31373 80 -31363
rect 0 -31433 10 -31373
rect 70 -31383 80 -31373
rect 320 -31373 400 -31363
rect 320 -31383 330 -31373
rect 70 -31433 330 -31383
rect 390 -31433 400 -31373
rect 0 -31443 400 -31433
rect 456 -31023 856 -31013
rect 456 -31083 466 -31023
rect 526 -31073 786 -31023
rect 526 -31083 536 -31073
rect 456 -31093 536 -31083
rect 776 -31083 786 -31073
rect 846 -31083 856 -31023
rect 776 -31093 856 -31083
rect 456 -31363 516 -31093
rect 596 -31153 626 -31133
rect 576 -31193 626 -31153
rect 686 -31153 716 -31133
rect 686 -31193 736 -31153
rect 576 -31263 736 -31193
rect 576 -31303 626 -31263
rect 596 -31323 626 -31303
rect 686 -31303 736 -31263
rect 686 -31323 716 -31303
rect 796 -31353 856 -31093
rect 786 -31363 856 -31353
rect 456 -31373 536 -31363
rect 456 -31433 466 -31373
rect 526 -31383 536 -31373
rect 776 -31373 856 -31363
rect 776 -31383 786 -31373
rect 526 -31433 786 -31383
rect 846 -31433 856 -31373
rect 456 -31443 856 -31433
rect 912 -31023 1312 -31013
rect 912 -31083 922 -31023
rect 982 -31073 1242 -31023
rect 982 -31083 992 -31073
rect 912 -31093 992 -31083
rect 1232 -31083 1242 -31073
rect 1302 -31083 1312 -31023
rect 1232 -31093 1312 -31083
rect 912 -31363 972 -31093
rect 1052 -31153 1082 -31133
rect 1032 -31193 1082 -31153
rect 1142 -31153 1172 -31133
rect 1142 -31193 1192 -31153
rect 1032 -31263 1192 -31193
rect 1032 -31303 1082 -31263
rect 1052 -31323 1082 -31303
rect 1142 -31303 1192 -31263
rect 1142 -31323 1172 -31303
rect 1252 -31353 1312 -31093
rect 1242 -31363 1312 -31353
rect 912 -31373 992 -31363
rect 912 -31433 922 -31373
rect 982 -31383 992 -31373
rect 1232 -31373 1312 -31363
rect 1232 -31383 1242 -31373
rect 982 -31433 1242 -31383
rect 1302 -31433 1312 -31373
rect 912 -31443 1312 -31433
rect 1370 -31023 1770 -31013
rect 1370 -31083 1380 -31023
rect 1440 -31073 1700 -31023
rect 1440 -31083 1450 -31073
rect 1370 -31093 1450 -31083
rect 1690 -31083 1700 -31073
rect 1760 -31083 1770 -31023
rect 1690 -31093 1770 -31083
rect 1370 -31363 1430 -31093
rect 1510 -31153 1540 -31133
rect 1490 -31193 1540 -31153
rect 1600 -31153 1630 -31133
rect 1600 -31193 1650 -31153
rect 1490 -31263 1650 -31193
rect 1490 -31303 1540 -31263
rect 1510 -31323 1540 -31303
rect 1600 -31303 1650 -31263
rect 1600 -31323 1630 -31303
rect 1710 -31353 1770 -31093
rect 1700 -31363 1770 -31353
rect 1370 -31373 1450 -31363
rect 1370 -31433 1380 -31373
rect 1440 -31383 1450 -31373
rect 1690 -31373 1770 -31363
rect 1690 -31383 1700 -31373
rect 1440 -31433 1700 -31383
rect 1760 -31433 1770 -31373
rect 1370 -31443 1770 -31433
rect 1826 -31023 2226 -31013
rect 1826 -31083 1836 -31023
rect 1896 -31073 2156 -31023
rect 1896 -31083 1906 -31073
rect 1826 -31093 1906 -31083
rect 2146 -31083 2156 -31073
rect 2216 -31083 2226 -31023
rect 2146 -31093 2226 -31083
rect 1826 -31363 1886 -31093
rect 1966 -31153 1996 -31133
rect 1946 -31193 1996 -31153
rect 2056 -31153 2086 -31133
rect 2056 -31193 2106 -31153
rect 1946 -31263 2106 -31193
rect 1946 -31303 1996 -31263
rect 1966 -31323 1996 -31303
rect 2056 -31303 2106 -31263
rect 2056 -31323 2086 -31303
rect 2166 -31353 2226 -31093
rect 2156 -31363 2226 -31353
rect 1826 -31373 1906 -31363
rect 1826 -31433 1836 -31373
rect 1896 -31383 1906 -31373
rect 2146 -31373 2226 -31363
rect 2146 -31383 2156 -31373
rect 1896 -31433 2156 -31383
rect 2216 -31433 2226 -31373
rect 1826 -31443 2226 -31433
rect 2282 -31023 2682 -31013
rect 2282 -31083 2292 -31023
rect 2352 -31073 2612 -31023
rect 2352 -31083 2362 -31073
rect 2282 -31093 2362 -31083
rect 2602 -31083 2612 -31073
rect 2672 -31083 2682 -31023
rect 2602 -31093 2682 -31083
rect 2282 -31363 2342 -31093
rect 2422 -31153 2452 -31133
rect 2402 -31193 2452 -31153
rect 2512 -31153 2542 -31133
rect 2512 -31193 2562 -31153
rect 2402 -31263 2562 -31193
rect 2402 -31303 2452 -31263
rect 2422 -31323 2452 -31303
rect 2512 -31303 2562 -31263
rect 2512 -31323 2542 -31303
rect 2622 -31353 2682 -31093
rect 2612 -31363 2682 -31353
rect 2282 -31373 2362 -31363
rect 2282 -31433 2292 -31373
rect 2352 -31383 2362 -31373
rect 2602 -31373 2682 -31363
rect 2602 -31383 2612 -31373
rect 2352 -31433 2612 -31383
rect 2672 -31433 2682 -31373
rect 2282 -31443 2682 -31433
rect 2740 -31023 3140 -31013
rect 2740 -31083 2750 -31023
rect 2810 -31073 3070 -31023
rect 2810 -31083 2820 -31073
rect 2740 -31093 2820 -31083
rect 3060 -31083 3070 -31073
rect 3130 -31083 3140 -31023
rect 3060 -31093 3140 -31083
rect 2740 -31363 2800 -31093
rect 2880 -31153 2910 -31133
rect 2860 -31193 2910 -31153
rect 2970 -31153 3000 -31133
rect 2970 -31193 3020 -31153
rect 2860 -31263 3020 -31193
rect 2860 -31303 2910 -31263
rect 2880 -31323 2910 -31303
rect 2970 -31303 3020 -31263
rect 2970 -31323 3000 -31303
rect 3080 -31353 3140 -31093
rect 3070 -31363 3140 -31353
rect 2740 -31373 2820 -31363
rect 2740 -31433 2750 -31373
rect 2810 -31383 2820 -31373
rect 3060 -31373 3140 -31363
rect 3060 -31383 3070 -31373
rect 2810 -31433 3070 -31383
rect 3130 -31433 3140 -31373
rect 2740 -31443 3140 -31433
rect 3196 -31023 3596 -31013
rect 3196 -31083 3206 -31023
rect 3266 -31073 3526 -31023
rect 3266 -31083 3276 -31073
rect 3196 -31093 3276 -31083
rect 3516 -31083 3526 -31073
rect 3586 -31083 3596 -31023
rect 3516 -31093 3596 -31083
rect 3196 -31363 3256 -31093
rect 3336 -31153 3366 -31133
rect 3316 -31193 3366 -31153
rect 3426 -31153 3456 -31133
rect 3426 -31193 3476 -31153
rect 3316 -31263 3476 -31193
rect 3316 -31303 3366 -31263
rect 3336 -31323 3366 -31303
rect 3426 -31303 3476 -31263
rect 3426 -31323 3456 -31303
rect 3536 -31353 3596 -31093
rect 3526 -31363 3596 -31353
rect 3196 -31373 3276 -31363
rect 3196 -31433 3206 -31373
rect 3266 -31383 3276 -31373
rect 3516 -31373 3596 -31363
rect 3516 -31383 3526 -31373
rect 3266 -31433 3526 -31383
rect 3586 -31433 3596 -31373
rect 3196 -31443 3596 -31433
rect 3652 -31023 4052 -31013
rect 3652 -31083 3662 -31023
rect 3722 -31073 3982 -31023
rect 3722 -31083 3732 -31073
rect 3652 -31093 3732 -31083
rect 3972 -31083 3982 -31073
rect 4042 -31083 4052 -31023
rect 3972 -31093 4052 -31083
rect 3652 -31363 3712 -31093
rect 3792 -31153 3822 -31133
rect 3772 -31193 3822 -31153
rect 3882 -31153 3912 -31133
rect 3882 -31193 3932 -31153
rect 3772 -31263 3932 -31193
rect 3772 -31303 3822 -31263
rect 3792 -31323 3822 -31303
rect 3882 -31303 3932 -31263
rect 3882 -31323 3912 -31303
rect 3992 -31353 4052 -31093
rect 3982 -31363 4052 -31353
rect 3652 -31373 3732 -31363
rect 3652 -31433 3662 -31373
rect 3722 -31383 3732 -31373
rect 3972 -31373 4052 -31363
rect 3972 -31383 3982 -31373
rect 3722 -31433 3982 -31383
rect 4042 -31433 4052 -31373
rect 3652 -31443 4052 -31433
rect 4110 -31023 4510 -31013
rect 4110 -31083 4120 -31023
rect 4180 -31073 4440 -31023
rect 4180 -31083 4190 -31073
rect 4110 -31093 4190 -31083
rect 4430 -31083 4440 -31073
rect 4500 -31083 4510 -31023
rect 4430 -31093 4510 -31083
rect 4110 -31363 4170 -31093
rect 4250 -31153 4280 -31133
rect 4230 -31193 4280 -31153
rect 4340 -31153 4370 -31133
rect 4340 -31193 4390 -31153
rect 4230 -31263 4390 -31193
rect 4230 -31303 4280 -31263
rect 4250 -31323 4280 -31303
rect 4340 -31303 4390 -31263
rect 4340 -31323 4370 -31303
rect 4450 -31353 4510 -31093
rect 4440 -31363 4510 -31353
rect 4110 -31373 4190 -31363
rect 4110 -31433 4120 -31373
rect 4180 -31383 4190 -31373
rect 4430 -31373 4510 -31363
rect 4430 -31383 4440 -31373
rect 4180 -31433 4440 -31383
rect 4500 -31433 4510 -31373
rect 4110 -31443 4510 -31433
rect 4566 -31023 4966 -31013
rect 4566 -31083 4576 -31023
rect 4636 -31073 4896 -31023
rect 4636 -31083 4646 -31073
rect 4566 -31093 4646 -31083
rect 4886 -31083 4896 -31073
rect 4956 -31083 4966 -31023
rect 4886 -31093 4966 -31083
rect 4566 -31363 4626 -31093
rect 4706 -31153 4736 -31133
rect 4686 -31193 4736 -31153
rect 4796 -31153 4826 -31133
rect 4796 -31193 4846 -31153
rect 4686 -31263 4846 -31193
rect 4686 -31303 4736 -31263
rect 4706 -31323 4736 -31303
rect 4796 -31303 4846 -31263
rect 4796 -31323 4826 -31303
rect 4906 -31353 4966 -31093
rect 4896 -31363 4966 -31353
rect 4566 -31373 4646 -31363
rect 4566 -31433 4576 -31373
rect 4636 -31383 4646 -31373
rect 4886 -31373 4966 -31363
rect 4886 -31383 4896 -31373
rect 4636 -31433 4896 -31383
rect 4956 -31433 4966 -31373
rect 4566 -31443 4966 -31433
rect 5022 -31023 5422 -31013
rect 5022 -31083 5032 -31023
rect 5092 -31073 5352 -31023
rect 5092 -31083 5102 -31073
rect 5022 -31093 5102 -31083
rect 5342 -31083 5352 -31073
rect 5412 -31083 5422 -31023
rect 5342 -31093 5422 -31083
rect 5022 -31363 5082 -31093
rect 5162 -31153 5192 -31133
rect 5142 -31193 5192 -31153
rect 5252 -31153 5282 -31133
rect 5252 -31193 5302 -31153
rect 5142 -31263 5302 -31193
rect 5142 -31303 5192 -31263
rect 5162 -31323 5192 -31303
rect 5252 -31303 5302 -31263
rect 5252 -31323 5282 -31303
rect 5362 -31353 5422 -31093
rect 5352 -31363 5422 -31353
rect 5022 -31373 5102 -31363
rect 5022 -31433 5032 -31373
rect 5092 -31383 5102 -31373
rect 5342 -31373 5422 -31363
rect 5342 -31383 5352 -31373
rect 5092 -31433 5352 -31383
rect 5412 -31433 5422 -31373
rect 5022 -31443 5422 -31433
rect 5480 -31023 5880 -31013
rect 5480 -31083 5490 -31023
rect 5550 -31073 5810 -31023
rect 5550 -31083 5560 -31073
rect 5480 -31093 5560 -31083
rect 5800 -31083 5810 -31073
rect 5870 -31083 5880 -31023
rect 5800 -31093 5880 -31083
rect 5480 -31363 5540 -31093
rect 5620 -31153 5650 -31133
rect 5600 -31193 5650 -31153
rect 5710 -31153 5740 -31133
rect 5710 -31193 5760 -31153
rect 5600 -31263 5760 -31193
rect 5600 -31303 5650 -31263
rect 5620 -31323 5650 -31303
rect 5710 -31303 5760 -31263
rect 5710 -31323 5740 -31303
rect 5820 -31353 5880 -31093
rect 5810 -31363 5880 -31353
rect 5480 -31373 5560 -31363
rect 5480 -31433 5490 -31373
rect 5550 -31383 5560 -31373
rect 5800 -31373 5880 -31363
rect 5800 -31383 5810 -31373
rect 5550 -31433 5810 -31383
rect 5870 -31433 5880 -31373
rect 5480 -31443 5880 -31433
rect 5936 -31023 6336 -31013
rect 5936 -31083 5946 -31023
rect 6006 -31073 6266 -31023
rect 6006 -31083 6016 -31073
rect 5936 -31093 6016 -31083
rect 6256 -31083 6266 -31073
rect 6326 -31083 6336 -31023
rect 6256 -31093 6336 -31083
rect 5936 -31363 5996 -31093
rect 6076 -31153 6106 -31133
rect 6056 -31193 6106 -31153
rect 6166 -31153 6196 -31133
rect 6166 -31193 6216 -31153
rect 6056 -31263 6216 -31193
rect 6056 -31303 6106 -31263
rect 6076 -31323 6106 -31303
rect 6166 -31303 6216 -31263
rect 6166 -31323 6196 -31303
rect 6276 -31353 6336 -31093
rect 6266 -31363 6336 -31353
rect 5936 -31373 6016 -31363
rect 5936 -31433 5946 -31373
rect 6006 -31383 6016 -31373
rect 6256 -31373 6336 -31363
rect 6256 -31383 6266 -31373
rect 6006 -31433 6266 -31383
rect 6326 -31433 6336 -31373
rect 5936 -31443 6336 -31433
rect 6392 -31023 6792 -31013
rect 6392 -31083 6402 -31023
rect 6462 -31073 6722 -31023
rect 6462 -31083 6472 -31073
rect 6392 -31093 6472 -31083
rect 6712 -31083 6722 -31073
rect 6782 -31083 6792 -31023
rect 6712 -31093 6792 -31083
rect 6392 -31363 6452 -31093
rect 6532 -31153 6562 -31133
rect 6512 -31193 6562 -31153
rect 6622 -31153 6652 -31133
rect 6622 -31193 6672 -31153
rect 6512 -31263 6672 -31193
rect 6512 -31303 6562 -31263
rect 6532 -31323 6562 -31303
rect 6622 -31303 6672 -31263
rect 6622 -31323 6652 -31303
rect 6732 -31353 6792 -31093
rect 6722 -31363 6792 -31353
rect 6392 -31373 6472 -31363
rect 6392 -31433 6402 -31373
rect 6462 -31383 6472 -31373
rect 6712 -31373 6792 -31363
rect 6712 -31383 6722 -31373
rect 6462 -31433 6722 -31383
rect 6782 -31433 6792 -31373
rect 6392 -31443 6792 -31433
rect 6850 -31023 7250 -31013
rect 6850 -31083 6860 -31023
rect 6920 -31073 7180 -31023
rect 6920 -31083 6930 -31073
rect 6850 -31093 6930 -31083
rect 7170 -31083 7180 -31073
rect 7240 -31083 7250 -31023
rect 7170 -31093 7250 -31083
rect 6850 -31363 6910 -31093
rect 6990 -31153 7020 -31133
rect 6970 -31193 7020 -31153
rect 7080 -31153 7110 -31133
rect 7080 -31193 7130 -31153
rect 6970 -31263 7130 -31193
rect 6970 -31303 7020 -31263
rect 6990 -31323 7020 -31303
rect 7080 -31303 7130 -31263
rect 7080 -31323 7110 -31303
rect 7190 -31353 7250 -31093
rect 7180 -31363 7250 -31353
rect 6850 -31373 6930 -31363
rect 6850 -31433 6860 -31373
rect 6920 -31383 6930 -31373
rect 7170 -31373 7250 -31363
rect 7170 -31383 7180 -31373
rect 6920 -31433 7180 -31383
rect 7240 -31433 7250 -31373
rect 6850 -31443 7250 -31433
rect 7306 -31023 7706 -31013
rect 7306 -31083 7316 -31023
rect 7376 -31073 7636 -31023
rect 7376 -31083 7386 -31073
rect 7306 -31093 7386 -31083
rect 7626 -31083 7636 -31073
rect 7696 -31083 7706 -31023
rect 7626 -31093 7706 -31083
rect 7306 -31363 7366 -31093
rect 7446 -31153 7476 -31133
rect 7426 -31193 7476 -31153
rect 7536 -31153 7566 -31133
rect 7536 -31193 7586 -31153
rect 7426 -31263 7586 -31193
rect 7426 -31303 7476 -31263
rect 7446 -31323 7476 -31303
rect 7536 -31303 7586 -31263
rect 7536 -31323 7566 -31303
rect 7646 -31353 7706 -31093
rect 7636 -31363 7706 -31353
rect 7306 -31373 7386 -31363
rect 7306 -31433 7316 -31373
rect 7376 -31383 7386 -31373
rect 7626 -31373 7706 -31363
rect 7626 -31383 7636 -31373
rect 7376 -31433 7636 -31383
rect 7696 -31433 7706 -31373
rect 7306 -31443 7706 -31433
rect 7762 -31023 8162 -31013
rect 7762 -31083 7772 -31023
rect 7832 -31073 8092 -31023
rect 7832 -31083 7842 -31073
rect 7762 -31093 7842 -31083
rect 8082 -31083 8092 -31073
rect 8152 -31083 8162 -31023
rect 8082 -31093 8162 -31083
rect 7762 -31363 7822 -31093
rect 7902 -31153 7932 -31133
rect 7882 -31193 7932 -31153
rect 7992 -31153 8022 -31133
rect 7992 -31193 8042 -31153
rect 7882 -31263 8042 -31193
rect 7882 -31303 7932 -31263
rect 7902 -31323 7932 -31303
rect 7992 -31303 8042 -31263
rect 7992 -31323 8022 -31303
rect 8102 -31353 8162 -31093
rect 8092 -31363 8162 -31353
rect 7762 -31373 7842 -31363
rect 7762 -31433 7772 -31373
rect 7832 -31383 7842 -31373
rect 8082 -31373 8162 -31363
rect 8082 -31383 8092 -31373
rect 7832 -31433 8092 -31383
rect 8152 -31433 8162 -31373
rect 7762 -31443 8162 -31433
rect 8236 -31023 8636 -31013
rect 8236 -31083 8246 -31023
rect 8306 -31073 8566 -31023
rect 8306 -31083 8316 -31073
rect 8236 -31093 8316 -31083
rect 8556 -31083 8566 -31073
rect 8626 -31083 8636 -31023
rect 8556 -31093 8636 -31083
rect 8236 -31363 8296 -31093
rect 8376 -31153 8406 -31133
rect 8356 -31193 8406 -31153
rect 8466 -31153 8496 -31133
rect 8466 -31193 8516 -31153
rect 8356 -31263 8516 -31193
rect 8356 -31303 8406 -31263
rect 8376 -31323 8406 -31303
rect 8466 -31303 8516 -31263
rect 8466 -31323 8496 -31303
rect 8576 -31353 8636 -31093
rect 8566 -31363 8636 -31353
rect 8236 -31373 8316 -31363
rect 8236 -31433 8246 -31373
rect 8306 -31383 8316 -31373
rect 8556 -31373 8636 -31363
rect 8556 -31383 8566 -31373
rect 8306 -31433 8566 -31383
rect 8626 -31433 8636 -31373
rect 8236 -31443 8636 -31433
rect 8692 -31023 9092 -31013
rect 8692 -31083 8702 -31023
rect 8762 -31073 9022 -31023
rect 8762 -31083 8772 -31073
rect 8692 -31093 8772 -31083
rect 9012 -31083 9022 -31073
rect 9082 -31083 9092 -31023
rect 9012 -31093 9092 -31083
rect 8692 -31363 8752 -31093
rect 8832 -31153 8862 -31133
rect 8812 -31193 8862 -31153
rect 8922 -31153 8952 -31133
rect 8922 -31193 8972 -31153
rect 8812 -31263 8972 -31193
rect 8812 -31303 8862 -31263
rect 8832 -31323 8862 -31303
rect 8922 -31303 8972 -31263
rect 8922 -31323 8952 -31303
rect 9032 -31353 9092 -31093
rect 9022 -31363 9092 -31353
rect 8692 -31373 8772 -31363
rect 8692 -31433 8702 -31373
rect 8762 -31383 8772 -31373
rect 9012 -31373 9092 -31363
rect 9012 -31383 9022 -31373
rect 8762 -31433 9022 -31383
rect 9082 -31433 9092 -31373
rect 8692 -31443 9092 -31433
rect 9150 -31023 9550 -31013
rect 9150 -31083 9160 -31023
rect 9220 -31073 9480 -31023
rect 9220 -31083 9230 -31073
rect 9150 -31093 9230 -31083
rect 9470 -31083 9480 -31073
rect 9540 -31083 9550 -31023
rect 9470 -31093 9550 -31083
rect 9150 -31363 9210 -31093
rect 9290 -31153 9320 -31133
rect 9270 -31193 9320 -31153
rect 9380 -31153 9410 -31133
rect 9380 -31193 9430 -31153
rect 9270 -31263 9430 -31193
rect 9270 -31303 9320 -31263
rect 9290 -31323 9320 -31303
rect 9380 -31303 9430 -31263
rect 9380 -31323 9410 -31303
rect 9490 -31353 9550 -31093
rect 9480 -31363 9550 -31353
rect 9150 -31373 9230 -31363
rect 9150 -31433 9160 -31373
rect 9220 -31383 9230 -31373
rect 9470 -31373 9550 -31363
rect 9470 -31383 9480 -31373
rect 9220 -31433 9480 -31383
rect 9540 -31433 9550 -31373
rect 9150 -31443 9550 -31433
rect 9606 -31023 10006 -31013
rect 9606 -31083 9616 -31023
rect 9676 -31073 9936 -31023
rect 9676 -31083 9686 -31073
rect 9606 -31093 9686 -31083
rect 9926 -31083 9936 -31073
rect 9996 -31083 10006 -31023
rect 9926 -31093 10006 -31083
rect 9606 -31363 9666 -31093
rect 9746 -31153 9776 -31133
rect 9726 -31193 9776 -31153
rect 9836 -31153 9866 -31133
rect 9836 -31193 9886 -31153
rect 9726 -31263 9886 -31193
rect 9726 -31303 9776 -31263
rect 9746 -31323 9776 -31303
rect 9836 -31303 9886 -31263
rect 9836 -31323 9866 -31303
rect 9946 -31353 10006 -31093
rect 9936 -31363 10006 -31353
rect 9606 -31373 9686 -31363
rect 9606 -31433 9616 -31373
rect 9676 -31383 9686 -31373
rect 9926 -31373 10006 -31363
rect 9926 -31383 9936 -31373
rect 9676 -31433 9936 -31383
rect 9996 -31433 10006 -31373
rect 9606 -31443 10006 -31433
rect 10062 -31023 10462 -31013
rect 10062 -31083 10072 -31023
rect 10132 -31073 10392 -31023
rect 10132 -31083 10142 -31073
rect 10062 -31093 10142 -31083
rect 10382 -31083 10392 -31073
rect 10452 -31083 10462 -31023
rect 10382 -31093 10462 -31083
rect 10062 -31363 10122 -31093
rect 10202 -31153 10232 -31133
rect 10182 -31193 10232 -31153
rect 10292 -31153 10322 -31133
rect 10292 -31193 10342 -31153
rect 10182 -31263 10342 -31193
rect 10182 -31303 10232 -31263
rect 10202 -31323 10232 -31303
rect 10292 -31303 10342 -31263
rect 10292 -31323 10322 -31303
rect 10402 -31353 10462 -31093
rect 10392 -31363 10462 -31353
rect 10062 -31373 10142 -31363
rect 10062 -31433 10072 -31373
rect 10132 -31383 10142 -31373
rect 10382 -31373 10462 -31363
rect 10382 -31383 10392 -31373
rect 10132 -31433 10392 -31383
rect 10452 -31433 10462 -31373
rect 10062 -31443 10462 -31433
rect 10520 -31023 10920 -31013
rect 10520 -31083 10530 -31023
rect 10590 -31073 10850 -31023
rect 10590 -31083 10600 -31073
rect 10520 -31093 10600 -31083
rect 10840 -31083 10850 -31073
rect 10910 -31083 10920 -31023
rect 10840 -31093 10920 -31083
rect 10520 -31363 10580 -31093
rect 10660 -31153 10690 -31133
rect 10640 -31193 10690 -31153
rect 10750 -31153 10780 -31133
rect 10750 -31193 10800 -31153
rect 10640 -31263 10800 -31193
rect 10640 -31303 10690 -31263
rect 10660 -31323 10690 -31303
rect 10750 -31303 10800 -31263
rect 10750 -31323 10780 -31303
rect 10860 -31353 10920 -31093
rect 10850 -31363 10920 -31353
rect 10520 -31373 10600 -31363
rect 10520 -31433 10530 -31373
rect 10590 -31383 10600 -31373
rect 10840 -31373 10920 -31363
rect 10840 -31383 10850 -31373
rect 10590 -31433 10850 -31383
rect 10910 -31433 10920 -31373
rect 10520 -31443 10920 -31433
rect 10976 -31023 11376 -31013
rect 10976 -31083 10986 -31023
rect 11046 -31073 11306 -31023
rect 11046 -31083 11056 -31073
rect 10976 -31093 11056 -31083
rect 11296 -31083 11306 -31073
rect 11366 -31083 11376 -31023
rect 11296 -31093 11376 -31083
rect 10976 -31363 11036 -31093
rect 11116 -31153 11146 -31133
rect 11096 -31193 11146 -31153
rect 11206 -31153 11236 -31133
rect 11206 -31193 11256 -31153
rect 11096 -31263 11256 -31193
rect 11096 -31303 11146 -31263
rect 11116 -31323 11146 -31303
rect 11206 -31303 11256 -31263
rect 11206 -31323 11236 -31303
rect 11316 -31353 11376 -31093
rect 11306 -31363 11376 -31353
rect 10976 -31373 11056 -31363
rect 10976 -31433 10986 -31373
rect 11046 -31383 11056 -31373
rect 11296 -31373 11376 -31363
rect 11296 -31383 11306 -31373
rect 11046 -31433 11306 -31383
rect 11366 -31433 11376 -31373
rect 10976 -31443 11376 -31433
rect 11432 -31023 11832 -31013
rect 11432 -31083 11442 -31023
rect 11502 -31073 11762 -31023
rect 11502 -31083 11512 -31073
rect 11432 -31093 11512 -31083
rect 11752 -31083 11762 -31073
rect 11822 -31083 11832 -31023
rect 11752 -31093 11832 -31083
rect 11432 -31363 11492 -31093
rect 11572 -31153 11602 -31133
rect 11552 -31193 11602 -31153
rect 11662 -31153 11692 -31133
rect 11662 -31193 11712 -31153
rect 11552 -31263 11712 -31193
rect 11552 -31303 11602 -31263
rect 11572 -31323 11602 -31303
rect 11662 -31303 11712 -31263
rect 11662 -31323 11692 -31303
rect 11772 -31353 11832 -31093
rect 11762 -31363 11832 -31353
rect 11432 -31373 11512 -31363
rect 11432 -31433 11442 -31373
rect 11502 -31383 11512 -31373
rect 11752 -31373 11832 -31363
rect 11752 -31383 11762 -31373
rect 11502 -31433 11762 -31383
rect 11822 -31433 11832 -31373
rect 11432 -31443 11832 -31433
rect 11890 -31023 12290 -31013
rect 11890 -31083 11900 -31023
rect 11960 -31073 12220 -31023
rect 11960 -31083 11970 -31073
rect 11890 -31093 11970 -31083
rect 12210 -31083 12220 -31073
rect 12280 -31083 12290 -31023
rect 12210 -31093 12290 -31083
rect 11890 -31363 11950 -31093
rect 12030 -31153 12060 -31133
rect 12010 -31193 12060 -31153
rect 12120 -31153 12150 -31133
rect 12120 -31193 12170 -31153
rect 12010 -31263 12170 -31193
rect 12010 -31303 12060 -31263
rect 12030 -31323 12060 -31303
rect 12120 -31303 12170 -31263
rect 12120 -31323 12150 -31303
rect 12230 -31353 12290 -31093
rect 12220 -31363 12290 -31353
rect 11890 -31373 11970 -31363
rect 11890 -31433 11900 -31373
rect 11960 -31383 11970 -31373
rect 12210 -31373 12290 -31363
rect 12210 -31383 12220 -31373
rect 11960 -31433 12220 -31383
rect 12280 -31433 12290 -31373
rect 11890 -31443 12290 -31433
rect 12346 -31023 12746 -31013
rect 12346 -31083 12356 -31023
rect 12416 -31073 12676 -31023
rect 12416 -31083 12426 -31073
rect 12346 -31093 12426 -31083
rect 12666 -31083 12676 -31073
rect 12736 -31083 12746 -31023
rect 12666 -31093 12746 -31083
rect 12346 -31363 12406 -31093
rect 12486 -31153 12516 -31133
rect 12466 -31193 12516 -31153
rect 12576 -31153 12606 -31133
rect 12576 -31193 12626 -31153
rect 12466 -31263 12626 -31193
rect 12466 -31303 12516 -31263
rect 12486 -31323 12516 -31303
rect 12576 -31303 12626 -31263
rect 12576 -31323 12606 -31303
rect 12686 -31353 12746 -31093
rect 12676 -31363 12746 -31353
rect 12346 -31373 12426 -31363
rect 12346 -31433 12356 -31373
rect 12416 -31383 12426 -31373
rect 12666 -31373 12746 -31363
rect 12666 -31383 12676 -31373
rect 12416 -31433 12676 -31383
rect 12736 -31433 12746 -31373
rect 12346 -31443 12746 -31433
rect 12802 -31023 13202 -31013
rect 12802 -31083 12812 -31023
rect 12872 -31073 13132 -31023
rect 12872 -31083 12882 -31073
rect 12802 -31093 12882 -31083
rect 13122 -31083 13132 -31073
rect 13192 -31083 13202 -31023
rect 13122 -31093 13202 -31083
rect 12802 -31363 12862 -31093
rect 12942 -31153 12972 -31133
rect 12922 -31193 12972 -31153
rect 13032 -31153 13062 -31133
rect 13032 -31193 13082 -31153
rect 12922 -31263 13082 -31193
rect 12922 -31303 12972 -31263
rect 12942 -31323 12972 -31303
rect 13032 -31303 13082 -31263
rect 13032 -31323 13062 -31303
rect 13142 -31353 13202 -31093
rect 13132 -31363 13202 -31353
rect 12802 -31373 12882 -31363
rect 12802 -31433 12812 -31373
rect 12872 -31383 12882 -31373
rect 13122 -31373 13202 -31363
rect 13122 -31383 13132 -31373
rect 12872 -31433 13132 -31383
rect 13192 -31433 13202 -31373
rect 12802 -31443 13202 -31433
rect 13260 -31023 13660 -31013
rect 13260 -31083 13270 -31023
rect 13330 -31073 13590 -31023
rect 13330 -31083 13340 -31073
rect 13260 -31093 13340 -31083
rect 13580 -31083 13590 -31073
rect 13650 -31083 13660 -31023
rect 13580 -31093 13660 -31083
rect 13260 -31363 13320 -31093
rect 13400 -31153 13430 -31133
rect 13380 -31193 13430 -31153
rect 13490 -31153 13520 -31133
rect 13490 -31193 13540 -31153
rect 13380 -31263 13540 -31193
rect 13380 -31303 13430 -31263
rect 13400 -31323 13430 -31303
rect 13490 -31303 13540 -31263
rect 13490 -31323 13520 -31303
rect 13600 -31353 13660 -31093
rect 13590 -31363 13660 -31353
rect 13260 -31373 13340 -31363
rect 13260 -31433 13270 -31373
rect 13330 -31383 13340 -31373
rect 13580 -31373 13660 -31363
rect 13580 -31383 13590 -31373
rect 13330 -31433 13590 -31383
rect 13650 -31433 13660 -31373
rect 13260 -31443 13660 -31433
rect 13716 -31023 14116 -31013
rect 13716 -31083 13726 -31023
rect 13786 -31073 14046 -31023
rect 13786 -31083 13796 -31073
rect 13716 -31093 13796 -31083
rect 14036 -31083 14046 -31073
rect 14106 -31083 14116 -31023
rect 14036 -31093 14116 -31083
rect 13716 -31363 13776 -31093
rect 13856 -31153 13886 -31133
rect 13836 -31193 13886 -31153
rect 13946 -31153 13976 -31133
rect 13946 -31193 13996 -31153
rect 13836 -31263 13996 -31193
rect 13836 -31303 13886 -31263
rect 13856 -31323 13886 -31303
rect 13946 -31303 13996 -31263
rect 13946 -31323 13976 -31303
rect 14056 -31353 14116 -31093
rect 14046 -31363 14116 -31353
rect 13716 -31373 13796 -31363
rect 13716 -31433 13726 -31373
rect 13786 -31383 13796 -31373
rect 14036 -31373 14116 -31363
rect 14036 -31383 14046 -31373
rect 13786 -31433 14046 -31383
rect 14106 -31433 14116 -31373
rect 13716 -31443 14116 -31433
rect 14172 -31023 14572 -31013
rect 14172 -31083 14182 -31023
rect 14242 -31073 14502 -31023
rect 14242 -31083 14252 -31073
rect 14172 -31093 14252 -31083
rect 14492 -31083 14502 -31073
rect 14562 -31083 14572 -31023
rect 14492 -31093 14572 -31083
rect 14172 -31363 14232 -31093
rect 14312 -31153 14342 -31133
rect 14292 -31193 14342 -31153
rect 14402 -31153 14432 -31133
rect 14402 -31193 14452 -31153
rect 14292 -31263 14452 -31193
rect 14292 -31303 14342 -31263
rect 14312 -31323 14342 -31303
rect 14402 -31303 14452 -31263
rect 14402 -31323 14432 -31303
rect 14512 -31353 14572 -31093
rect 14502 -31363 14572 -31353
rect 14172 -31373 14252 -31363
rect 14172 -31433 14182 -31373
rect 14242 -31383 14252 -31373
rect 14492 -31373 14572 -31363
rect 14492 -31383 14502 -31373
rect 14242 -31433 14502 -31383
rect 14562 -31433 14572 -31373
rect 14172 -31443 14572 -31433
rect 14630 -31023 15030 -31013
rect 14630 -31083 14640 -31023
rect 14700 -31073 14960 -31023
rect 14700 -31083 14710 -31073
rect 14630 -31093 14710 -31083
rect 14950 -31083 14960 -31073
rect 15020 -31083 15030 -31023
rect 14950 -31093 15030 -31083
rect 14630 -31363 14690 -31093
rect 14770 -31153 14800 -31133
rect 14750 -31193 14800 -31153
rect 14860 -31153 14890 -31133
rect 14860 -31193 14910 -31153
rect 14750 -31263 14910 -31193
rect 14750 -31303 14800 -31263
rect 14770 -31323 14800 -31303
rect 14860 -31303 14910 -31263
rect 14860 -31323 14890 -31303
rect 14970 -31353 15030 -31093
rect 14960 -31363 15030 -31353
rect 14630 -31373 14710 -31363
rect 14630 -31433 14640 -31373
rect 14700 -31383 14710 -31373
rect 14950 -31373 15030 -31363
rect 14950 -31383 14960 -31373
rect 14700 -31433 14960 -31383
rect 15020 -31433 15030 -31373
rect 14630 -31443 15030 -31433
rect 15086 -31023 15486 -31013
rect 15086 -31083 15096 -31023
rect 15156 -31073 15416 -31023
rect 15156 -31083 15166 -31073
rect 15086 -31093 15166 -31083
rect 15406 -31083 15416 -31073
rect 15476 -31083 15486 -31023
rect 15406 -31093 15486 -31083
rect 15086 -31363 15146 -31093
rect 15226 -31153 15256 -31133
rect 15206 -31193 15256 -31153
rect 15316 -31153 15346 -31133
rect 15316 -31193 15366 -31153
rect 15206 -31263 15366 -31193
rect 15206 -31303 15256 -31263
rect 15226 -31323 15256 -31303
rect 15316 -31303 15366 -31263
rect 15316 -31323 15346 -31303
rect 15426 -31353 15486 -31093
rect 15416 -31363 15486 -31353
rect 15086 -31373 15166 -31363
rect 15086 -31433 15096 -31373
rect 15156 -31383 15166 -31373
rect 15406 -31373 15486 -31363
rect 15406 -31383 15416 -31373
rect 15156 -31433 15416 -31383
rect 15476 -31433 15486 -31373
rect 15086 -31443 15486 -31433
rect 0 -31525 400 -31515
rect 0 -31585 10 -31525
rect 70 -31575 330 -31525
rect 70 -31585 80 -31575
rect 0 -31595 80 -31585
rect 320 -31585 330 -31575
rect 390 -31585 400 -31525
rect 320 -31595 400 -31585
rect 0 -31865 60 -31595
rect 140 -31655 170 -31635
rect 120 -31695 170 -31655
rect 230 -31655 260 -31635
rect 230 -31695 280 -31655
rect 120 -31765 280 -31695
rect 120 -31805 170 -31765
rect 140 -31825 170 -31805
rect 230 -31805 280 -31765
rect 230 -31825 260 -31805
rect 340 -31855 400 -31595
rect 330 -31865 400 -31855
rect 0 -31875 80 -31865
rect 0 -31935 10 -31875
rect 70 -31885 80 -31875
rect 320 -31875 400 -31865
rect 320 -31885 330 -31875
rect 70 -31935 330 -31885
rect 390 -31935 400 -31875
rect 0 -31945 400 -31935
rect 456 -31525 856 -31515
rect 456 -31585 466 -31525
rect 526 -31575 786 -31525
rect 526 -31585 536 -31575
rect 456 -31595 536 -31585
rect 776 -31585 786 -31575
rect 846 -31585 856 -31525
rect 776 -31595 856 -31585
rect 456 -31865 516 -31595
rect 596 -31655 626 -31635
rect 576 -31695 626 -31655
rect 686 -31655 716 -31635
rect 686 -31695 736 -31655
rect 576 -31765 736 -31695
rect 576 -31805 626 -31765
rect 596 -31825 626 -31805
rect 686 -31805 736 -31765
rect 686 -31825 716 -31805
rect 796 -31855 856 -31595
rect 786 -31865 856 -31855
rect 456 -31875 536 -31865
rect 456 -31935 466 -31875
rect 526 -31885 536 -31875
rect 776 -31875 856 -31865
rect 776 -31885 786 -31875
rect 526 -31935 786 -31885
rect 846 -31935 856 -31875
rect 456 -31945 856 -31935
rect 912 -31525 1312 -31515
rect 912 -31585 922 -31525
rect 982 -31575 1242 -31525
rect 982 -31585 992 -31575
rect 912 -31595 992 -31585
rect 1232 -31585 1242 -31575
rect 1302 -31585 1312 -31525
rect 1232 -31595 1312 -31585
rect 912 -31865 972 -31595
rect 1052 -31655 1082 -31635
rect 1032 -31695 1082 -31655
rect 1142 -31655 1172 -31635
rect 1142 -31695 1192 -31655
rect 1032 -31765 1192 -31695
rect 1032 -31805 1082 -31765
rect 1052 -31825 1082 -31805
rect 1142 -31805 1192 -31765
rect 1142 -31825 1172 -31805
rect 1252 -31855 1312 -31595
rect 1242 -31865 1312 -31855
rect 912 -31875 992 -31865
rect 912 -31935 922 -31875
rect 982 -31885 992 -31875
rect 1232 -31875 1312 -31865
rect 1232 -31885 1242 -31875
rect 982 -31935 1242 -31885
rect 1302 -31935 1312 -31875
rect 912 -31945 1312 -31935
rect 1370 -31525 1770 -31515
rect 1370 -31585 1380 -31525
rect 1440 -31575 1700 -31525
rect 1440 -31585 1450 -31575
rect 1370 -31595 1450 -31585
rect 1690 -31585 1700 -31575
rect 1760 -31585 1770 -31525
rect 1690 -31595 1770 -31585
rect 1370 -31865 1430 -31595
rect 1510 -31655 1540 -31635
rect 1490 -31695 1540 -31655
rect 1600 -31655 1630 -31635
rect 1600 -31695 1650 -31655
rect 1490 -31765 1650 -31695
rect 1490 -31805 1540 -31765
rect 1510 -31825 1540 -31805
rect 1600 -31805 1650 -31765
rect 1600 -31825 1630 -31805
rect 1710 -31855 1770 -31595
rect 1700 -31865 1770 -31855
rect 1370 -31875 1450 -31865
rect 1370 -31935 1380 -31875
rect 1440 -31885 1450 -31875
rect 1690 -31875 1770 -31865
rect 1690 -31885 1700 -31875
rect 1440 -31935 1700 -31885
rect 1760 -31935 1770 -31875
rect 1370 -31945 1770 -31935
rect 1826 -31525 2226 -31515
rect 1826 -31585 1836 -31525
rect 1896 -31575 2156 -31525
rect 1896 -31585 1906 -31575
rect 1826 -31595 1906 -31585
rect 2146 -31585 2156 -31575
rect 2216 -31585 2226 -31525
rect 2146 -31595 2226 -31585
rect 1826 -31865 1886 -31595
rect 1966 -31655 1996 -31635
rect 1946 -31695 1996 -31655
rect 2056 -31655 2086 -31635
rect 2056 -31695 2106 -31655
rect 1946 -31765 2106 -31695
rect 1946 -31805 1996 -31765
rect 1966 -31825 1996 -31805
rect 2056 -31805 2106 -31765
rect 2056 -31825 2086 -31805
rect 2166 -31855 2226 -31595
rect 2156 -31865 2226 -31855
rect 1826 -31875 1906 -31865
rect 1826 -31935 1836 -31875
rect 1896 -31885 1906 -31875
rect 2146 -31875 2226 -31865
rect 2146 -31885 2156 -31875
rect 1896 -31935 2156 -31885
rect 2216 -31935 2226 -31875
rect 1826 -31945 2226 -31935
rect 2282 -31525 2682 -31515
rect 2282 -31585 2292 -31525
rect 2352 -31575 2612 -31525
rect 2352 -31585 2362 -31575
rect 2282 -31595 2362 -31585
rect 2602 -31585 2612 -31575
rect 2672 -31585 2682 -31525
rect 2602 -31595 2682 -31585
rect 2282 -31865 2342 -31595
rect 2422 -31655 2452 -31635
rect 2402 -31695 2452 -31655
rect 2512 -31655 2542 -31635
rect 2512 -31695 2562 -31655
rect 2402 -31765 2562 -31695
rect 2402 -31805 2452 -31765
rect 2422 -31825 2452 -31805
rect 2512 -31805 2562 -31765
rect 2512 -31825 2542 -31805
rect 2622 -31855 2682 -31595
rect 2612 -31865 2682 -31855
rect 2282 -31875 2362 -31865
rect 2282 -31935 2292 -31875
rect 2352 -31885 2362 -31875
rect 2602 -31875 2682 -31865
rect 2602 -31885 2612 -31875
rect 2352 -31935 2612 -31885
rect 2672 -31935 2682 -31875
rect 2282 -31945 2682 -31935
rect 2740 -31525 3140 -31515
rect 2740 -31585 2750 -31525
rect 2810 -31575 3070 -31525
rect 2810 -31585 2820 -31575
rect 2740 -31595 2820 -31585
rect 3060 -31585 3070 -31575
rect 3130 -31585 3140 -31525
rect 3060 -31595 3140 -31585
rect 2740 -31865 2800 -31595
rect 2880 -31655 2910 -31635
rect 2860 -31695 2910 -31655
rect 2970 -31655 3000 -31635
rect 2970 -31695 3020 -31655
rect 2860 -31765 3020 -31695
rect 2860 -31805 2910 -31765
rect 2880 -31825 2910 -31805
rect 2970 -31805 3020 -31765
rect 2970 -31825 3000 -31805
rect 3080 -31855 3140 -31595
rect 3070 -31865 3140 -31855
rect 2740 -31875 2820 -31865
rect 2740 -31935 2750 -31875
rect 2810 -31885 2820 -31875
rect 3060 -31875 3140 -31865
rect 3060 -31885 3070 -31875
rect 2810 -31935 3070 -31885
rect 3130 -31935 3140 -31875
rect 2740 -31945 3140 -31935
rect 3196 -31525 3596 -31515
rect 3196 -31585 3206 -31525
rect 3266 -31575 3526 -31525
rect 3266 -31585 3276 -31575
rect 3196 -31595 3276 -31585
rect 3516 -31585 3526 -31575
rect 3586 -31585 3596 -31525
rect 3516 -31595 3596 -31585
rect 3196 -31865 3256 -31595
rect 3336 -31655 3366 -31635
rect 3316 -31695 3366 -31655
rect 3426 -31655 3456 -31635
rect 3426 -31695 3476 -31655
rect 3316 -31765 3476 -31695
rect 3316 -31805 3366 -31765
rect 3336 -31825 3366 -31805
rect 3426 -31805 3476 -31765
rect 3426 -31825 3456 -31805
rect 3536 -31855 3596 -31595
rect 3526 -31865 3596 -31855
rect 3196 -31875 3276 -31865
rect 3196 -31935 3206 -31875
rect 3266 -31885 3276 -31875
rect 3516 -31875 3596 -31865
rect 3516 -31885 3526 -31875
rect 3266 -31935 3526 -31885
rect 3586 -31935 3596 -31875
rect 3196 -31945 3596 -31935
rect 3652 -31525 4052 -31515
rect 3652 -31585 3662 -31525
rect 3722 -31575 3982 -31525
rect 3722 -31585 3732 -31575
rect 3652 -31595 3732 -31585
rect 3972 -31585 3982 -31575
rect 4042 -31585 4052 -31525
rect 3972 -31595 4052 -31585
rect 3652 -31865 3712 -31595
rect 3792 -31655 3822 -31635
rect 3772 -31695 3822 -31655
rect 3882 -31655 3912 -31635
rect 3882 -31695 3932 -31655
rect 3772 -31765 3932 -31695
rect 3772 -31805 3822 -31765
rect 3792 -31825 3822 -31805
rect 3882 -31805 3932 -31765
rect 3882 -31825 3912 -31805
rect 3992 -31855 4052 -31595
rect 3982 -31865 4052 -31855
rect 3652 -31875 3732 -31865
rect 3652 -31935 3662 -31875
rect 3722 -31885 3732 -31875
rect 3972 -31875 4052 -31865
rect 3972 -31885 3982 -31875
rect 3722 -31935 3982 -31885
rect 4042 -31935 4052 -31875
rect 3652 -31945 4052 -31935
rect 4110 -31525 4510 -31515
rect 4110 -31585 4120 -31525
rect 4180 -31575 4440 -31525
rect 4180 -31585 4190 -31575
rect 4110 -31595 4190 -31585
rect 4430 -31585 4440 -31575
rect 4500 -31585 4510 -31525
rect 4430 -31595 4510 -31585
rect 4110 -31865 4170 -31595
rect 4250 -31655 4280 -31635
rect 4230 -31695 4280 -31655
rect 4340 -31655 4370 -31635
rect 4340 -31695 4390 -31655
rect 4230 -31765 4390 -31695
rect 4230 -31805 4280 -31765
rect 4250 -31825 4280 -31805
rect 4340 -31805 4390 -31765
rect 4340 -31825 4370 -31805
rect 4450 -31855 4510 -31595
rect 4440 -31865 4510 -31855
rect 4110 -31875 4190 -31865
rect 4110 -31935 4120 -31875
rect 4180 -31885 4190 -31875
rect 4430 -31875 4510 -31865
rect 4430 -31885 4440 -31875
rect 4180 -31935 4440 -31885
rect 4500 -31935 4510 -31875
rect 4110 -31945 4510 -31935
rect 4566 -31525 4966 -31515
rect 4566 -31585 4576 -31525
rect 4636 -31575 4896 -31525
rect 4636 -31585 4646 -31575
rect 4566 -31595 4646 -31585
rect 4886 -31585 4896 -31575
rect 4956 -31585 4966 -31525
rect 4886 -31595 4966 -31585
rect 4566 -31865 4626 -31595
rect 4706 -31655 4736 -31635
rect 4686 -31695 4736 -31655
rect 4796 -31655 4826 -31635
rect 4796 -31695 4846 -31655
rect 4686 -31765 4846 -31695
rect 4686 -31805 4736 -31765
rect 4706 -31825 4736 -31805
rect 4796 -31805 4846 -31765
rect 4796 -31825 4826 -31805
rect 4906 -31855 4966 -31595
rect 4896 -31865 4966 -31855
rect 4566 -31875 4646 -31865
rect 4566 -31935 4576 -31875
rect 4636 -31885 4646 -31875
rect 4886 -31875 4966 -31865
rect 4886 -31885 4896 -31875
rect 4636 -31935 4896 -31885
rect 4956 -31935 4966 -31875
rect 4566 -31945 4966 -31935
rect 5022 -31525 5422 -31515
rect 5022 -31585 5032 -31525
rect 5092 -31575 5352 -31525
rect 5092 -31585 5102 -31575
rect 5022 -31595 5102 -31585
rect 5342 -31585 5352 -31575
rect 5412 -31585 5422 -31525
rect 5342 -31595 5422 -31585
rect 5022 -31865 5082 -31595
rect 5162 -31655 5192 -31635
rect 5142 -31695 5192 -31655
rect 5252 -31655 5282 -31635
rect 5252 -31695 5302 -31655
rect 5142 -31765 5302 -31695
rect 5142 -31805 5192 -31765
rect 5162 -31825 5192 -31805
rect 5252 -31805 5302 -31765
rect 5252 -31825 5282 -31805
rect 5362 -31855 5422 -31595
rect 5352 -31865 5422 -31855
rect 5022 -31875 5102 -31865
rect 5022 -31935 5032 -31875
rect 5092 -31885 5102 -31875
rect 5342 -31875 5422 -31865
rect 5342 -31885 5352 -31875
rect 5092 -31935 5352 -31885
rect 5412 -31935 5422 -31875
rect 5022 -31945 5422 -31935
rect 5480 -31525 5880 -31515
rect 5480 -31585 5490 -31525
rect 5550 -31575 5810 -31525
rect 5550 -31585 5560 -31575
rect 5480 -31595 5560 -31585
rect 5800 -31585 5810 -31575
rect 5870 -31585 5880 -31525
rect 5800 -31595 5880 -31585
rect 5480 -31865 5540 -31595
rect 5620 -31655 5650 -31635
rect 5600 -31695 5650 -31655
rect 5710 -31655 5740 -31635
rect 5710 -31695 5760 -31655
rect 5600 -31765 5760 -31695
rect 5600 -31805 5650 -31765
rect 5620 -31825 5650 -31805
rect 5710 -31805 5760 -31765
rect 5710 -31825 5740 -31805
rect 5820 -31855 5880 -31595
rect 5810 -31865 5880 -31855
rect 5480 -31875 5560 -31865
rect 5480 -31935 5490 -31875
rect 5550 -31885 5560 -31875
rect 5800 -31875 5880 -31865
rect 5800 -31885 5810 -31875
rect 5550 -31935 5810 -31885
rect 5870 -31935 5880 -31875
rect 5480 -31945 5880 -31935
rect 5936 -31525 6336 -31515
rect 5936 -31585 5946 -31525
rect 6006 -31575 6266 -31525
rect 6006 -31585 6016 -31575
rect 5936 -31595 6016 -31585
rect 6256 -31585 6266 -31575
rect 6326 -31585 6336 -31525
rect 6256 -31595 6336 -31585
rect 5936 -31865 5996 -31595
rect 6076 -31655 6106 -31635
rect 6056 -31695 6106 -31655
rect 6166 -31655 6196 -31635
rect 6166 -31695 6216 -31655
rect 6056 -31765 6216 -31695
rect 6056 -31805 6106 -31765
rect 6076 -31825 6106 -31805
rect 6166 -31805 6216 -31765
rect 6166 -31825 6196 -31805
rect 6276 -31855 6336 -31595
rect 6266 -31865 6336 -31855
rect 5936 -31875 6016 -31865
rect 5936 -31935 5946 -31875
rect 6006 -31885 6016 -31875
rect 6256 -31875 6336 -31865
rect 6256 -31885 6266 -31875
rect 6006 -31935 6266 -31885
rect 6326 -31935 6336 -31875
rect 5936 -31945 6336 -31935
rect 6392 -31525 6792 -31515
rect 6392 -31585 6402 -31525
rect 6462 -31575 6722 -31525
rect 6462 -31585 6472 -31575
rect 6392 -31595 6472 -31585
rect 6712 -31585 6722 -31575
rect 6782 -31585 6792 -31525
rect 6712 -31595 6792 -31585
rect 6392 -31865 6452 -31595
rect 6532 -31655 6562 -31635
rect 6512 -31695 6562 -31655
rect 6622 -31655 6652 -31635
rect 6622 -31695 6672 -31655
rect 6512 -31765 6672 -31695
rect 6512 -31805 6562 -31765
rect 6532 -31825 6562 -31805
rect 6622 -31805 6672 -31765
rect 6622 -31825 6652 -31805
rect 6732 -31855 6792 -31595
rect 6722 -31865 6792 -31855
rect 6392 -31875 6472 -31865
rect 6392 -31935 6402 -31875
rect 6462 -31885 6472 -31875
rect 6712 -31875 6792 -31865
rect 6712 -31885 6722 -31875
rect 6462 -31935 6722 -31885
rect 6782 -31935 6792 -31875
rect 6392 -31945 6792 -31935
rect 6850 -31525 7250 -31515
rect 6850 -31585 6860 -31525
rect 6920 -31575 7180 -31525
rect 6920 -31585 6930 -31575
rect 6850 -31595 6930 -31585
rect 7170 -31585 7180 -31575
rect 7240 -31585 7250 -31525
rect 7170 -31595 7250 -31585
rect 6850 -31865 6910 -31595
rect 6990 -31655 7020 -31635
rect 6970 -31695 7020 -31655
rect 7080 -31655 7110 -31635
rect 7080 -31695 7130 -31655
rect 6970 -31765 7130 -31695
rect 6970 -31805 7020 -31765
rect 6990 -31825 7020 -31805
rect 7080 -31805 7130 -31765
rect 7080 -31825 7110 -31805
rect 7190 -31855 7250 -31595
rect 7180 -31865 7250 -31855
rect 6850 -31875 6930 -31865
rect 6850 -31935 6860 -31875
rect 6920 -31885 6930 -31875
rect 7170 -31875 7250 -31865
rect 7170 -31885 7180 -31875
rect 6920 -31935 7180 -31885
rect 7240 -31935 7250 -31875
rect 6850 -31945 7250 -31935
rect 7306 -31525 7706 -31515
rect 7306 -31585 7316 -31525
rect 7376 -31575 7636 -31525
rect 7376 -31585 7386 -31575
rect 7306 -31595 7386 -31585
rect 7626 -31585 7636 -31575
rect 7696 -31585 7706 -31525
rect 7626 -31595 7706 -31585
rect 7306 -31865 7366 -31595
rect 7446 -31655 7476 -31635
rect 7426 -31695 7476 -31655
rect 7536 -31655 7566 -31635
rect 7536 -31695 7586 -31655
rect 7426 -31765 7586 -31695
rect 7426 -31805 7476 -31765
rect 7446 -31825 7476 -31805
rect 7536 -31805 7586 -31765
rect 7536 -31825 7566 -31805
rect 7646 -31855 7706 -31595
rect 7636 -31865 7706 -31855
rect 7306 -31875 7386 -31865
rect 7306 -31935 7316 -31875
rect 7376 -31885 7386 -31875
rect 7626 -31875 7706 -31865
rect 7626 -31885 7636 -31875
rect 7376 -31935 7636 -31885
rect 7696 -31935 7706 -31875
rect 7306 -31945 7706 -31935
rect 7762 -31525 8162 -31515
rect 7762 -31585 7772 -31525
rect 7832 -31575 8092 -31525
rect 7832 -31585 7842 -31575
rect 7762 -31595 7842 -31585
rect 8082 -31585 8092 -31575
rect 8152 -31585 8162 -31525
rect 8082 -31595 8162 -31585
rect 7762 -31865 7822 -31595
rect 7902 -31655 7932 -31635
rect 7882 -31695 7932 -31655
rect 7992 -31655 8022 -31635
rect 7992 -31695 8042 -31655
rect 7882 -31765 8042 -31695
rect 7882 -31805 7932 -31765
rect 7902 -31825 7932 -31805
rect 7992 -31805 8042 -31765
rect 7992 -31825 8022 -31805
rect 8102 -31855 8162 -31595
rect 8092 -31865 8162 -31855
rect 7762 -31875 7842 -31865
rect 7762 -31935 7772 -31875
rect 7832 -31885 7842 -31875
rect 8082 -31875 8162 -31865
rect 8082 -31885 8092 -31875
rect 7832 -31935 8092 -31885
rect 8152 -31935 8162 -31875
rect 7762 -31945 8162 -31935
rect 8236 -31525 8636 -31515
rect 8236 -31585 8246 -31525
rect 8306 -31575 8566 -31525
rect 8306 -31585 8316 -31575
rect 8236 -31595 8316 -31585
rect 8556 -31585 8566 -31575
rect 8626 -31585 8636 -31525
rect 8556 -31595 8636 -31585
rect 8236 -31865 8296 -31595
rect 8376 -31655 8406 -31635
rect 8356 -31695 8406 -31655
rect 8466 -31655 8496 -31635
rect 8466 -31695 8516 -31655
rect 8356 -31765 8516 -31695
rect 8356 -31805 8406 -31765
rect 8376 -31825 8406 -31805
rect 8466 -31805 8516 -31765
rect 8466 -31825 8496 -31805
rect 8576 -31855 8636 -31595
rect 8566 -31865 8636 -31855
rect 8236 -31875 8316 -31865
rect 8236 -31935 8246 -31875
rect 8306 -31885 8316 -31875
rect 8556 -31875 8636 -31865
rect 8556 -31885 8566 -31875
rect 8306 -31935 8566 -31885
rect 8626 -31935 8636 -31875
rect 8236 -31945 8636 -31935
rect 8692 -31525 9092 -31515
rect 8692 -31585 8702 -31525
rect 8762 -31575 9022 -31525
rect 8762 -31585 8772 -31575
rect 8692 -31595 8772 -31585
rect 9012 -31585 9022 -31575
rect 9082 -31585 9092 -31525
rect 9012 -31595 9092 -31585
rect 8692 -31865 8752 -31595
rect 8832 -31655 8862 -31635
rect 8812 -31695 8862 -31655
rect 8922 -31655 8952 -31635
rect 8922 -31695 8972 -31655
rect 8812 -31765 8972 -31695
rect 8812 -31805 8862 -31765
rect 8832 -31825 8862 -31805
rect 8922 -31805 8972 -31765
rect 8922 -31825 8952 -31805
rect 9032 -31855 9092 -31595
rect 9022 -31865 9092 -31855
rect 8692 -31875 8772 -31865
rect 8692 -31935 8702 -31875
rect 8762 -31885 8772 -31875
rect 9012 -31875 9092 -31865
rect 9012 -31885 9022 -31875
rect 8762 -31935 9022 -31885
rect 9082 -31935 9092 -31875
rect 8692 -31945 9092 -31935
rect 9150 -31525 9550 -31515
rect 9150 -31585 9160 -31525
rect 9220 -31575 9480 -31525
rect 9220 -31585 9230 -31575
rect 9150 -31595 9230 -31585
rect 9470 -31585 9480 -31575
rect 9540 -31585 9550 -31525
rect 9470 -31595 9550 -31585
rect 9150 -31865 9210 -31595
rect 9290 -31655 9320 -31635
rect 9270 -31695 9320 -31655
rect 9380 -31655 9410 -31635
rect 9380 -31695 9430 -31655
rect 9270 -31765 9430 -31695
rect 9270 -31805 9320 -31765
rect 9290 -31825 9320 -31805
rect 9380 -31805 9430 -31765
rect 9380 -31825 9410 -31805
rect 9490 -31855 9550 -31595
rect 9480 -31865 9550 -31855
rect 9150 -31875 9230 -31865
rect 9150 -31935 9160 -31875
rect 9220 -31885 9230 -31875
rect 9470 -31875 9550 -31865
rect 9470 -31885 9480 -31875
rect 9220 -31935 9480 -31885
rect 9540 -31935 9550 -31875
rect 9150 -31945 9550 -31935
rect 9606 -31525 10006 -31515
rect 9606 -31585 9616 -31525
rect 9676 -31575 9936 -31525
rect 9676 -31585 9686 -31575
rect 9606 -31595 9686 -31585
rect 9926 -31585 9936 -31575
rect 9996 -31585 10006 -31525
rect 9926 -31595 10006 -31585
rect 9606 -31865 9666 -31595
rect 9746 -31655 9776 -31635
rect 9726 -31695 9776 -31655
rect 9836 -31655 9866 -31635
rect 9836 -31695 9886 -31655
rect 9726 -31765 9886 -31695
rect 9726 -31805 9776 -31765
rect 9746 -31825 9776 -31805
rect 9836 -31805 9886 -31765
rect 9836 -31825 9866 -31805
rect 9946 -31855 10006 -31595
rect 9936 -31865 10006 -31855
rect 9606 -31875 9686 -31865
rect 9606 -31935 9616 -31875
rect 9676 -31885 9686 -31875
rect 9926 -31875 10006 -31865
rect 9926 -31885 9936 -31875
rect 9676 -31935 9936 -31885
rect 9996 -31935 10006 -31875
rect 9606 -31945 10006 -31935
rect 10062 -31525 10462 -31515
rect 10062 -31585 10072 -31525
rect 10132 -31575 10392 -31525
rect 10132 -31585 10142 -31575
rect 10062 -31595 10142 -31585
rect 10382 -31585 10392 -31575
rect 10452 -31585 10462 -31525
rect 10382 -31595 10462 -31585
rect 10062 -31865 10122 -31595
rect 10202 -31655 10232 -31635
rect 10182 -31695 10232 -31655
rect 10292 -31655 10322 -31635
rect 10292 -31695 10342 -31655
rect 10182 -31765 10342 -31695
rect 10182 -31805 10232 -31765
rect 10202 -31825 10232 -31805
rect 10292 -31805 10342 -31765
rect 10292 -31825 10322 -31805
rect 10402 -31855 10462 -31595
rect 10392 -31865 10462 -31855
rect 10062 -31875 10142 -31865
rect 10062 -31935 10072 -31875
rect 10132 -31885 10142 -31875
rect 10382 -31875 10462 -31865
rect 10382 -31885 10392 -31875
rect 10132 -31935 10392 -31885
rect 10452 -31935 10462 -31875
rect 10062 -31945 10462 -31935
rect 10520 -31525 10920 -31515
rect 10520 -31585 10530 -31525
rect 10590 -31575 10850 -31525
rect 10590 -31585 10600 -31575
rect 10520 -31595 10600 -31585
rect 10840 -31585 10850 -31575
rect 10910 -31585 10920 -31525
rect 10840 -31595 10920 -31585
rect 10520 -31865 10580 -31595
rect 10660 -31655 10690 -31635
rect 10640 -31695 10690 -31655
rect 10750 -31655 10780 -31635
rect 10750 -31695 10800 -31655
rect 10640 -31765 10800 -31695
rect 10640 -31805 10690 -31765
rect 10660 -31825 10690 -31805
rect 10750 -31805 10800 -31765
rect 10750 -31825 10780 -31805
rect 10860 -31855 10920 -31595
rect 10850 -31865 10920 -31855
rect 10520 -31875 10600 -31865
rect 10520 -31935 10530 -31875
rect 10590 -31885 10600 -31875
rect 10840 -31875 10920 -31865
rect 10840 -31885 10850 -31875
rect 10590 -31935 10850 -31885
rect 10910 -31935 10920 -31875
rect 10520 -31945 10920 -31935
rect 10976 -31525 11376 -31515
rect 10976 -31585 10986 -31525
rect 11046 -31575 11306 -31525
rect 11046 -31585 11056 -31575
rect 10976 -31595 11056 -31585
rect 11296 -31585 11306 -31575
rect 11366 -31585 11376 -31525
rect 11296 -31595 11376 -31585
rect 10976 -31865 11036 -31595
rect 11116 -31655 11146 -31635
rect 11096 -31695 11146 -31655
rect 11206 -31655 11236 -31635
rect 11206 -31695 11256 -31655
rect 11096 -31765 11256 -31695
rect 11096 -31805 11146 -31765
rect 11116 -31825 11146 -31805
rect 11206 -31805 11256 -31765
rect 11206 -31825 11236 -31805
rect 11316 -31855 11376 -31595
rect 11306 -31865 11376 -31855
rect 10976 -31875 11056 -31865
rect 10976 -31935 10986 -31875
rect 11046 -31885 11056 -31875
rect 11296 -31875 11376 -31865
rect 11296 -31885 11306 -31875
rect 11046 -31935 11306 -31885
rect 11366 -31935 11376 -31875
rect 10976 -31945 11376 -31935
rect 11432 -31525 11832 -31515
rect 11432 -31585 11442 -31525
rect 11502 -31575 11762 -31525
rect 11502 -31585 11512 -31575
rect 11432 -31595 11512 -31585
rect 11752 -31585 11762 -31575
rect 11822 -31585 11832 -31525
rect 11752 -31595 11832 -31585
rect 11432 -31865 11492 -31595
rect 11572 -31655 11602 -31635
rect 11552 -31695 11602 -31655
rect 11662 -31655 11692 -31635
rect 11662 -31695 11712 -31655
rect 11552 -31765 11712 -31695
rect 11552 -31805 11602 -31765
rect 11572 -31825 11602 -31805
rect 11662 -31805 11712 -31765
rect 11662 -31825 11692 -31805
rect 11772 -31855 11832 -31595
rect 11762 -31865 11832 -31855
rect 11432 -31875 11512 -31865
rect 11432 -31935 11442 -31875
rect 11502 -31885 11512 -31875
rect 11752 -31875 11832 -31865
rect 11752 -31885 11762 -31875
rect 11502 -31935 11762 -31885
rect 11822 -31935 11832 -31875
rect 11432 -31945 11832 -31935
rect 11890 -31525 12290 -31515
rect 11890 -31585 11900 -31525
rect 11960 -31575 12220 -31525
rect 11960 -31585 11970 -31575
rect 11890 -31595 11970 -31585
rect 12210 -31585 12220 -31575
rect 12280 -31585 12290 -31525
rect 12210 -31595 12290 -31585
rect 11890 -31865 11950 -31595
rect 12030 -31655 12060 -31635
rect 12010 -31695 12060 -31655
rect 12120 -31655 12150 -31635
rect 12120 -31695 12170 -31655
rect 12010 -31765 12170 -31695
rect 12010 -31805 12060 -31765
rect 12030 -31825 12060 -31805
rect 12120 -31805 12170 -31765
rect 12120 -31825 12150 -31805
rect 12230 -31855 12290 -31595
rect 12220 -31865 12290 -31855
rect 11890 -31875 11970 -31865
rect 11890 -31935 11900 -31875
rect 11960 -31885 11970 -31875
rect 12210 -31875 12290 -31865
rect 12210 -31885 12220 -31875
rect 11960 -31935 12220 -31885
rect 12280 -31935 12290 -31875
rect 11890 -31945 12290 -31935
rect 12346 -31525 12746 -31515
rect 12346 -31585 12356 -31525
rect 12416 -31575 12676 -31525
rect 12416 -31585 12426 -31575
rect 12346 -31595 12426 -31585
rect 12666 -31585 12676 -31575
rect 12736 -31585 12746 -31525
rect 12666 -31595 12746 -31585
rect 12346 -31865 12406 -31595
rect 12486 -31655 12516 -31635
rect 12466 -31695 12516 -31655
rect 12576 -31655 12606 -31635
rect 12576 -31695 12626 -31655
rect 12466 -31765 12626 -31695
rect 12466 -31805 12516 -31765
rect 12486 -31825 12516 -31805
rect 12576 -31805 12626 -31765
rect 12576 -31825 12606 -31805
rect 12686 -31855 12746 -31595
rect 12676 -31865 12746 -31855
rect 12346 -31875 12426 -31865
rect 12346 -31935 12356 -31875
rect 12416 -31885 12426 -31875
rect 12666 -31875 12746 -31865
rect 12666 -31885 12676 -31875
rect 12416 -31935 12676 -31885
rect 12736 -31935 12746 -31875
rect 12346 -31945 12746 -31935
rect 12802 -31525 13202 -31515
rect 12802 -31585 12812 -31525
rect 12872 -31575 13132 -31525
rect 12872 -31585 12882 -31575
rect 12802 -31595 12882 -31585
rect 13122 -31585 13132 -31575
rect 13192 -31585 13202 -31525
rect 13122 -31595 13202 -31585
rect 12802 -31865 12862 -31595
rect 12942 -31655 12972 -31635
rect 12922 -31695 12972 -31655
rect 13032 -31655 13062 -31635
rect 13032 -31695 13082 -31655
rect 12922 -31765 13082 -31695
rect 12922 -31805 12972 -31765
rect 12942 -31825 12972 -31805
rect 13032 -31805 13082 -31765
rect 13032 -31825 13062 -31805
rect 13142 -31855 13202 -31595
rect 13132 -31865 13202 -31855
rect 12802 -31875 12882 -31865
rect 12802 -31935 12812 -31875
rect 12872 -31885 12882 -31875
rect 13122 -31875 13202 -31865
rect 13122 -31885 13132 -31875
rect 12872 -31935 13132 -31885
rect 13192 -31935 13202 -31875
rect 12802 -31945 13202 -31935
rect 13260 -31525 13660 -31515
rect 13260 -31585 13270 -31525
rect 13330 -31575 13590 -31525
rect 13330 -31585 13340 -31575
rect 13260 -31595 13340 -31585
rect 13580 -31585 13590 -31575
rect 13650 -31585 13660 -31525
rect 13580 -31595 13660 -31585
rect 13260 -31865 13320 -31595
rect 13400 -31655 13430 -31635
rect 13380 -31695 13430 -31655
rect 13490 -31655 13520 -31635
rect 13490 -31695 13540 -31655
rect 13380 -31765 13540 -31695
rect 13380 -31805 13430 -31765
rect 13400 -31825 13430 -31805
rect 13490 -31805 13540 -31765
rect 13490 -31825 13520 -31805
rect 13600 -31855 13660 -31595
rect 13590 -31865 13660 -31855
rect 13260 -31875 13340 -31865
rect 13260 -31935 13270 -31875
rect 13330 -31885 13340 -31875
rect 13580 -31875 13660 -31865
rect 13580 -31885 13590 -31875
rect 13330 -31935 13590 -31885
rect 13650 -31935 13660 -31875
rect 13260 -31945 13660 -31935
rect 13716 -31525 14116 -31515
rect 13716 -31585 13726 -31525
rect 13786 -31575 14046 -31525
rect 13786 -31585 13796 -31575
rect 13716 -31595 13796 -31585
rect 14036 -31585 14046 -31575
rect 14106 -31585 14116 -31525
rect 14036 -31595 14116 -31585
rect 13716 -31865 13776 -31595
rect 13856 -31655 13886 -31635
rect 13836 -31695 13886 -31655
rect 13946 -31655 13976 -31635
rect 13946 -31695 13996 -31655
rect 13836 -31765 13996 -31695
rect 13836 -31805 13886 -31765
rect 13856 -31825 13886 -31805
rect 13946 -31805 13996 -31765
rect 13946 -31825 13976 -31805
rect 14056 -31855 14116 -31595
rect 14046 -31865 14116 -31855
rect 13716 -31875 13796 -31865
rect 13716 -31935 13726 -31875
rect 13786 -31885 13796 -31875
rect 14036 -31875 14116 -31865
rect 14036 -31885 14046 -31875
rect 13786 -31935 14046 -31885
rect 14106 -31935 14116 -31875
rect 13716 -31945 14116 -31935
rect 14172 -31525 14572 -31515
rect 14172 -31585 14182 -31525
rect 14242 -31575 14502 -31525
rect 14242 -31585 14252 -31575
rect 14172 -31595 14252 -31585
rect 14492 -31585 14502 -31575
rect 14562 -31585 14572 -31525
rect 14492 -31595 14572 -31585
rect 14172 -31865 14232 -31595
rect 14312 -31655 14342 -31635
rect 14292 -31695 14342 -31655
rect 14402 -31655 14432 -31635
rect 14402 -31695 14452 -31655
rect 14292 -31765 14452 -31695
rect 14292 -31805 14342 -31765
rect 14312 -31825 14342 -31805
rect 14402 -31805 14452 -31765
rect 14402 -31825 14432 -31805
rect 14512 -31855 14572 -31595
rect 14502 -31865 14572 -31855
rect 14172 -31875 14252 -31865
rect 14172 -31935 14182 -31875
rect 14242 -31885 14252 -31875
rect 14492 -31875 14572 -31865
rect 14492 -31885 14502 -31875
rect 14242 -31935 14502 -31885
rect 14562 -31935 14572 -31875
rect 14172 -31945 14572 -31935
rect 14630 -31525 15030 -31515
rect 14630 -31585 14640 -31525
rect 14700 -31575 14960 -31525
rect 14700 -31585 14710 -31575
rect 14630 -31595 14710 -31585
rect 14950 -31585 14960 -31575
rect 15020 -31585 15030 -31525
rect 14950 -31595 15030 -31585
rect 14630 -31865 14690 -31595
rect 14770 -31655 14800 -31635
rect 14750 -31695 14800 -31655
rect 14860 -31655 14890 -31635
rect 14860 -31695 14910 -31655
rect 14750 -31765 14910 -31695
rect 14750 -31805 14800 -31765
rect 14770 -31825 14800 -31805
rect 14860 -31805 14910 -31765
rect 14860 -31825 14890 -31805
rect 14970 -31855 15030 -31595
rect 14960 -31865 15030 -31855
rect 14630 -31875 14710 -31865
rect 14630 -31935 14640 -31875
rect 14700 -31885 14710 -31875
rect 14950 -31875 15030 -31865
rect 14950 -31885 14960 -31875
rect 14700 -31935 14960 -31885
rect 15020 -31935 15030 -31875
rect 14630 -31945 15030 -31935
rect 15086 -31525 15486 -31515
rect 15086 -31585 15096 -31525
rect 15156 -31575 15416 -31525
rect 15156 -31585 15166 -31575
rect 15086 -31595 15166 -31585
rect 15406 -31585 15416 -31575
rect 15476 -31585 15486 -31525
rect 15406 -31595 15486 -31585
rect 15086 -31865 15146 -31595
rect 15226 -31655 15256 -31635
rect 15206 -31695 15256 -31655
rect 15316 -31655 15346 -31635
rect 15316 -31695 15366 -31655
rect 15206 -31765 15366 -31695
rect 15206 -31805 15256 -31765
rect 15226 -31825 15256 -31805
rect 15316 -31805 15366 -31765
rect 15316 -31825 15346 -31805
rect 15426 -31855 15486 -31595
rect 15416 -31865 15486 -31855
rect 15086 -31875 15166 -31865
rect 15086 -31935 15096 -31875
rect 15156 -31885 15166 -31875
rect 15406 -31875 15486 -31865
rect 15406 -31885 15416 -31875
rect 15156 -31935 15416 -31885
rect 15476 -31935 15486 -31875
rect 15086 -31945 15486 -31935
rect 0 -32017 400 -32007
rect 0 -32077 10 -32017
rect 70 -32067 330 -32017
rect 70 -32077 80 -32067
rect 0 -32087 80 -32077
rect 320 -32077 330 -32067
rect 390 -32077 400 -32017
rect 320 -32087 400 -32077
rect 0 -32357 60 -32087
rect 140 -32147 170 -32127
rect 120 -32187 170 -32147
rect 230 -32147 260 -32127
rect 230 -32187 280 -32147
rect 120 -32257 280 -32187
rect 120 -32297 170 -32257
rect 140 -32317 170 -32297
rect 230 -32297 280 -32257
rect 230 -32317 260 -32297
rect 340 -32347 400 -32087
rect 330 -32357 400 -32347
rect 0 -32367 80 -32357
rect 0 -32427 10 -32367
rect 70 -32377 80 -32367
rect 320 -32367 400 -32357
rect 320 -32377 330 -32367
rect 70 -32427 330 -32377
rect 390 -32427 400 -32367
rect 0 -32437 400 -32427
rect 456 -32017 856 -32007
rect 456 -32077 466 -32017
rect 526 -32067 786 -32017
rect 526 -32077 536 -32067
rect 456 -32087 536 -32077
rect 776 -32077 786 -32067
rect 846 -32077 856 -32017
rect 776 -32087 856 -32077
rect 456 -32357 516 -32087
rect 596 -32147 626 -32127
rect 576 -32187 626 -32147
rect 686 -32147 716 -32127
rect 686 -32187 736 -32147
rect 576 -32257 736 -32187
rect 576 -32297 626 -32257
rect 596 -32317 626 -32297
rect 686 -32297 736 -32257
rect 686 -32317 716 -32297
rect 796 -32347 856 -32087
rect 786 -32357 856 -32347
rect 456 -32367 536 -32357
rect 456 -32427 466 -32367
rect 526 -32377 536 -32367
rect 776 -32367 856 -32357
rect 776 -32377 786 -32367
rect 526 -32427 786 -32377
rect 846 -32427 856 -32367
rect 456 -32437 856 -32427
rect 912 -32017 1312 -32007
rect 912 -32077 922 -32017
rect 982 -32067 1242 -32017
rect 982 -32077 992 -32067
rect 912 -32087 992 -32077
rect 1232 -32077 1242 -32067
rect 1302 -32077 1312 -32017
rect 1232 -32087 1312 -32077
rect 912 -32357 972 -32087
rect 1052 -32147 1082 -32127
rect 1032 -32187 1082 -32147
rect 1142 -32147 1172 -32127
rect 1142 -32187 1192 -32147
rect 1032 -32257 1192 -32187
rect 1032 -32297 1082 -32257
rect 1052 -32317 1082 -32297
rect 1142 -32297 1192 -32257
rect 1142 -32317 1172 -32297
rect 1252 -32347 1312 -32087
rect 1242 -32357 1312 -32347
rect 912 -32367 992 -32357
rect 912 -32427 922 -32367
rect 982 -32377 992 -32367
rect 1232 -32367 1312 -32357
rect 1232 -32377 1242 -32367
rect 982 -32427 1242 -32377
rect 1302 -32427 1312 -32367
rect 912 -32437 1312 -32427
rect 1370 -32017 1770 -32007
rect 1370 -32077 1380 -32017
rect 1440 -32067 1700 -32017
rect 1440 -32077 1450 -32067
rect 1370 -32087 1450 -32077
rect 1690 -32077 1700 -32067
rect 1760 -32077 1770 -32017
rect 1690 -32087 1770 -32077
rect 1370 -32357 1430 -32087
rect 1510 -32147 1540 -32127
rect 1490 -32187 1540 -32147
rect 1600 -32147 1630 -32127
rect 1600 -32187 1650 -32147
rect 1490 -32257 1650 -32187
rect 1490 -32297 1540 -32257
rect 1510 -32317 1540 -32297
rect 1600 -32297 1650 -32257
rect 1600 -32317 1630 -32297
rect 1710 -32347 1770 -32087
rect 1700 -32357 1770 -32347
rect 1370 -32367 1450 -32357
rect 1370 -32427 1380 -32367
rect 1440 -32377 1450 -32367
rect 1690 -32367 1770 -32357
rect 1690 -32377 1700 -32367
rect 1440 -32427 1700 -32377
rect 1760 -32427 1770 -32367
rect 1370 -32437 1770 -32427
rect 1826 -32017 2226 -32007
rect 1826 -32077 1836 -32017
rect 1896 -32067 2156 -32017
rect 1896 -32077 1906 -32067
rect 1826 -32087 1906 -32077
rect 2146 -32077 2156 -32067
rect 2216 -32077 2226 -32017
rect 2146 -32087 2226 -32077
rect 1826 -32357 1886 -32087
rect 1966 -32147 1996 -32127
rect 1946 -32187 1996 -32147
rect 2056 -32147 2086 -32127
rect 2056 -32187 2106 -32147
rect 1946 -32257 2106 -32187
rect 1946 -32297 1996 -32257
rect 1966 -32317 1996 -32297
rect 2056 -32297 2106 -32257
rect 2056 -32317 2086 -32297
rect 2166 -32347 2226 -32087
rect 2156 -32357 2226 -32347
rect 1826 -32367 1906 -32357
rect 1826 -32427 1836 -32367
rect 1896 -32377 1906 -32367
rect 2146 -32367 2226 -32357
rect 2146 -32377 2156 -32367
rect 1896 -32427 2156 -32377
rect 2216 -32427 2226 -32367
rect 1826 -32437 2226 -32427
rect 2282 -32017 2682 -32007
rect 2282 -32077 2292 -32017
rect 2352 -32067 2612 -32017
rect 2352 -32077 2362 -32067
rect 2282 -32087 2362 -32077
rect 2602 -32077 2612 -32067
rect 2672 -32077 2682 -32017
rect 2602 -32087 2682 -32077
rect 2282 -32357 2342 -32087
rect 2422 -32147 2452 -32127
rect 2402 -32187 2452 -32147
rect 2512 -32147 2542 -32127
rect 2512 -32187 2562 -32147
rect 2402 -32257 2562 -32187
rect 2402 -32297 2452 -32257
rect 2422 -32317 2452 -32297
rect 2512 -32297 2562 -32257
rect 2512 -32317 2542 -32297
rect 2622 -32347 2682 -32087
rect 2612 -32357 2682 -32347
rect 2282 -32367 2362 -32357
rect 2282 -32427 2292 -32367
rect 2352 -32377 2362 -32367
rect 2602 -32367 2682 -32357
rect 2602 -32377 2612 -32367
rect 2352 -32427 2612 -32377
rect 2672 -32427 2682 -32367
rect 2282 -32437 2682 -32427
rect 2740 -32017 3140 -32007
rect 2740 -32077 2750 -32017
rect 2810 -32067 3070 -32017
rect 2810 -32077 2820 -32067
rect 2740 -32087 2820 -32077
rect 3060 -32077 3070 -32067
rect 3130 -32077 3140 -32017
rect 3060 -32087 3140 -32077
rect 2740 -32357 2800 -32087
rect 2880 -32147 2910 -32127
rect 2860 -32187 2910 -32147
rect 2970 -32147 3000 -32127
rect 2970 -32187 3020 -32147
rect 2860 -32257 3020 -32187
rect 2860 -32297 2910 -32257
rect 2880 -32317 2910 -32297
rect 2970 -32297 3020 -32257
rect 2970 -32317 3000 -32297
rect 3080 -32347 3140 -32087
rect 3070 -32357 3140 -32347
rect 2740 -32367 2820 -32357
rect 2740 -32427 2750 -32367
rect 2810 -32377 2820 -32367
rect 3060 -32367 3140 -32357
rect 3060 -32377 3070 -32367
rect 2810 -32427 3070 -32377
rect 3130 -32427 3140 -32367
rect 2740 -32437 3140 -32427
rect 3196 -32017 3596 -32007
rect 3196 -32077 3206 -32017
rect 3266 -32067 3526 -32017
rect 3266 -32077 3276 -32067
rect 3196 -32087 3276 -32077
rect 3516 -32077 3526 -32067
rect 3586 -32077 3596 -32017
rect 3516 -32087 3596 -32077
rect 3196 -32357 3256 -32087
rect 3336 -32147 3366 -32127
rect 3316 -32187 3366 -32147
rect 3426 -32147 3456 -32127
rect 3426 -32187 3476 -32147
rect 3316 -32257 3476 -32187
rect 3316 -32297 3366 -32257
rect 3336 -32317 3366 -32297
rect 3426 -32297 3476 -32257
rect 3426 -32317 3456 -32297
rect 3536 -32347 3596 -32087
rect 3526 -32357 3596 -32347
rect 3196 -32367 3276 -32357
rect 3196 -32427 3206 -32367
rect 3266 -32377 3276 -32367
rect 3516 -32367 3596 -32357
rect 3516 -32377 3526 -32367
rect 3266 -32427 3526 -32377
rect 3586 -32427 3596 -32367
rect 3196 -32437 3596 -32427
rect 3652 -32017 4052 -32007
rect 3652 -32077 3662 -32017
rect 3722 -32067 3982 -32017
rect 3722 -32077 3732 -32067
rect 3652 -32087 3732 -32077
rect 3972 -32077 3982 -32067
rect 4042 -32077 4052 -32017
rect 3972 -32087 4052 -32077
rect 3652 -32357 3712 -32087
rect 3792 -32147 3822 -32127
rect 3772 -32187 3822 -32147
rect 3882 -32147 3912 -32127
rect 3882 -32187 3932 -32147
rect 3772 -32257 3932 -32187
rect 3772 -32297 3822 -32257
rect 3792 -32317 3822 -32297
rect 3882 -32297 3932 -32257
rect 3882 -32317 3912 -32297
rect 3992 -32347 4052 -32087
rect 3982 -32357 4052 -32347
rect 3652 -32367 3732 -32357
rect 3652 -32427 3662 -32367
rect 3722 -32377 3732 -32367
rect 3972 -32367 4052 -32357
rect 3972 -32377 3982 -32367
rect 3722 -32427 3982 -32377
rect 4042 -32427 4052 -32367
rect 3652 -32437 4052 -32427
rect 4110 -32017 4510 -32007
rect 4110 -32077 4120 -32017
rect 4180 -32067 4440 -32017
rect 4180 -32077 4190 -32067
rect 4110 -32087 4190 -32077
rect 4430 -32077 4440 -32067
rect 4500 -32077 4510 -32017
rect 4430 -32087 4510 -32077
rect 4110 -32357 4170 -32087
rect 4250 -32147 4280 -32127
rect 4230 -32187 4280 -32147
rect 4340 -32147 4370 -32127
rect 4340 -32187 4390 -32147
rect 4230 -32257 4390 -32187
rect 4230 -32297 4280 -32257
rect 4250 -32317 4280 -32297
rect 4340 -32297 4390 -32257
rect 4340 -32317 4370 -32297
rect 4450 -32347 4510 -32087
rect 4440 -32357 4510 -32347
rect 4110 -32367 4190 -32357
rect 4110 -32427 4120 -32367
rect 4180 -32377 4190 -32367
rect 4430 -32367 4510 -32357
rect 4430 -32377 4440 -32367
rect 4180 -32427 4440 -32377
rect 4500 -32427 4510 -32367
rect 4110 -32437 4510 -32427
rect 4566 -32017 4966 -32007
rect 4566 -32077 4576 -32017
rect 4636 -32067 4896 -32017
rect 4636 -32077 4646 -32067
rect 4566 -32087 4646 -32077
rect 4886 -32077 4896 -32067
rect 4956 -32077 4966 -32017
rect 4886 -32087 4966 -32077
rect 4566 -32357 4626 -32087
rect 4706 -32147 4736 -32127
rect 4686 -32187 4736 -32147
rect 4796 -32147 4826 -32127
rect 4796 -32187 4846 -32147
rect 4686 -32257 4846 -32187
rect 4686 -32297 4736 -32257
rect 4706 -32317 4736 -32297
rect 4796 -32297 4846 -32257
rect 4796 -32317 4826 -32297
rect 4906 -32347 4966 -32087
rect 4896 -32357 4966 -32347
rect 4566 -32367 4646 -32357
rect 4566 -32427 4576 -32367
rect 4636 -32377 4646 -32367
rect 4886 -32367 4966 -32357
rect 4886 -32377 4896 -32367
rect 4636 -32427 4896 -32377
rect 4956 -32427 4966 -32367
rect 4566 -32437 4966 -32427
rect 5022 -32017 5422 -32007
rect 5022 -32077 5032 -32017
rect 5092 -32067 5352 -32017
rect 5092 -32077 5102 -32067
rect 5022 -32087 5102 -32077
rect 5342 -32077 5352 -32067
rect 5412 -32077 5422 -32017
rect 5342 -32087 5422 -32077
rect 5022 -32357 5082 -32087
rect 5162 -32147 5192 -32127
rect 5142 -32187 5192 -32147
rect 5252 -32147 5282 -32127
rect 5252 -32187 5302 -32147
rect 5142 -32257 5302 -32187
rect 5142 -32297 5192 -32257
rect 5162 -32317 5192 -32297
rect 5252 -32297 5302 -32257
rect 5252 -32317 5282 -32297
rect 5362 -32347 5422 -32087
rect 5352 -32357 5422 -32347
rect 5022 -32367 5102 -32357
rect 5022 -32427 5032 -32367
rect 5092 -32377 5102 -32367
rect 5342 -32367 5422 -32357
rect 5342 -32377 5352 -32367
rect 5092 -32427 5352 -32377
rect 5412 -32427 5422 -32367
rect 5022 -32437 5422 -32427
rect 5480 -32017 5880 -32007
rect 5480 -32077 5490 -32017
rect 5550 -32067 5810 -32017
rect 5550 -32077 5560 -32067
rect 5480 -32087 5560 -32077
rect 5800 -32077 5810 -32067
rect 5870 -32077 5880 -32017
rect 5800 -32087 5880 -32077
rect 5480 -32357 5540 -32087
rect 5620 -32147 5650 -32127
rect 5600 -32187 5650 -32147
rect 5710 -32147 5740 -32127
rect 5710 -32187 5760 -32147
rect 5600 -32257 5760 -32187
rect 5600 -32297 5650 -32257
rect 5620 -32317 5650 -32297
rect 5710 -32297 5760 -32257
rect 5710 -32317 5740 -32297
rect 5820 -32347 5880 -32087
rect 5810 -32357 5880 -32347
rect 5480 -32367 5560 -32357
rect 5480 -32427 5490 -32367
rect 5550 -32377 5560 -32367
rect 5800 -32367 5880 -32357
rect 5800 -32377 5810 -32367
rect 5550 -32427 5810 -32377
rect 5870 -32427 5880 -32367
rect 5480 -32437 5880 -32427
rect 5936 -32017 6336 -32007
rect 5936 -32077 5946 -32017
rect 6006 -32067 6266 -32017
rect 6006 -32077 6016 -32067
rect 5936 -32087 6016 -32077
rect 6256 -32077 6266 -32067
rect 6326 -32077 6336 -32017
rect 6256 -32087 6336 -32077
rect 5936 -32357 5996 -32087
rect 6076 -32147 6106 -32127
rect 6056 -32187 6106 -32147
rect 6166 -32147 6196 -32127
rect 6166 -32187 6216 -32147
rect 6056 -32257 6216 -32187
rect 6056 -32297 6106 -32257
rect 6076 -32317 6106 -32297
rect 6166 -32297 6216 -32257
rect 6166 -32317 6196 -32297
rect 6276 -32347 6336 -32087
rect 6266 -32357 6336 -32347
rect 5936 -32367 6016 -32357
rect 5936 -32427 5946 -32367
rect 6006 -32377 6016 -32367
rect 6256 -32367 6336 -32357
rect 6256 -32377 6266 -32367
rect 6006 -32427 6266 -32377
rect 6326 -32427 6336 -32367
rect 5936 -32437 6336 -32427
rect 6392 -32017 6792 -32007
rect 6392 -32077 6402 -32017
rect 6462 -32067 6722 -32017
rect 6462 -32077 6472 -32067
rect 6392 -32087 6472 -32077
rect 6712 -32077 6722 -32067
rect 6782 -32077 6792 -32017
rect 6712 -32087 6792 -32077
rect 6392 -32357 6452 -32087
rect 6532 -32147 6562 -32127
rect 6512 -32187 6562 -32147
rect 6622 -32147 6652 -32127
rect 6622 -32187 6672 -32147
rect 6512 -32257 6672 -32187
rect 6512 -32297 6562 -32257
rect 6532 -32317 6562 -32297
rect 6622 -32297 6672 -32257
rect 6622 -32317 6652 -32297
rect 6732 -32347 6792 -32087
rect 6722 -32357 6792 -32347
rect 6392 -32367 6472 -32357
rect 6392 -32427 6402 -32367
rect 6462 -32377 6472 -32367
rect 6712 -32367 6792 -32357
rect 6712 -32377 6722 -32367
rect 6462 -32427 6722 -32377
rect 6782 -32427 6792 -32367
rect 6392 -32437 6792 -32427
rect 6850 -32017 7250 -32007
rect 6850 -32077 6860 -32017
rect 6920 -32067 7180 -32017
rect 6920 -32077 6930 -32067
rect 6850 -32087 6930 -32077
rect 7170 -32077 7180 -32067
rect 7240 -32077 7250 -32017
rect 7170 -32087 7250 -32077
rect 6850 -32357 6910 -32087
rect 6990 -32147 7020 -32127
rect 6970 -32187 7020 -32147
rect 7080 -32147 7110 -32127
rect 7080 -32187 7130 -32147
rect 6970 -32257 7130 -32187
rect 6970 -32297 7020 -32257
rect 6990 -32317 7020 -32297
rect 7080 -32297 7130 -32257
rect 7080 -32317 7110 -32297
rect 7190 -32347 7250 -32087
rect 7180 -32357 7250 -32347
rect 6850 -32367 6930 -32357
rect 6850 -32427 6860 -32367
rect 6920 -32377 6930 -32367
rect 7170 -32367 7250 -32357
rect 7170 -32377 7180 -32367
rect 6920 -32427 7180 -32377
rect 7240 -32427 7250 -32367
rect 6850 -32437 7250 -32427
rect 7306 -32017 7706 -32007
rect 7306 -32077 7316 -32017
rect 7376 -32067 7636 -32017
rect 7376 -32077 7386 -32067
rect 7306 -32087 7386 -32077
rect 7626 -32077 7636 -32067
rect 7696 -32077 7706 -32017
rect 7626 -32087 7706 -32077
rect 7306 -32357 7366 -32087
rect 7446 -32147 7476 -32127
rect 7426 -32187 7476 -32147
rect 7536 -32147 7566 -32127
rect 7536 -32187 7586 -32147
rect 7426 -32257 7586 -32187
rect 7426 -32297 7476 -32257
rect 7446 -32317 7476 -32297
rect 7536 -32297 7586 -32257
rect 7536 -32317 7566 -32297
rect 7646 -32347 7706 -32087
rect 7636 -32357 7706 -32347
rect 7306 -32367 7386 -32357
rect 7306 -32427 7316 -32367
rect 7376 -32377 7386 -32367
rect 7626 -32367 7706 -32357
rect 7626 -32377 7636 -32367
rect 7376 -32427 7636 -32377
rect 7696 -32427 7706 -32367
rect 7306 -32437 7706 -32427
rect 7762 -32017 8162 -32007
rect 7762 -32077 7772 -32017
rect 7832 -32067 8092 -32017
rect 7832 -32077 7842 -32067
rect 7762 -32087 7842 -32077
rect 8082 -32077 8092 -32067
rect 8152 -32077 8162 -32017
rect 8082 -32087 8162 -32077
rect 7762 -32357 7822 -32087
rect 7902 -32147 7932 -32127
rect 7882 -32187 7932 -32147
rect 7992 -32147 8022 -32127
rect 7992 -32187 8042 -32147
rect 7882 -32257 8042 -32187
rect 7882 -32297 7932 -32257
rect 7902 -32317 7932 -32297
rect 7992 -32297 8042 -32257
rect 7992 -32317 8022 -32297
rect 8102 -32347 8162 -32087
rect 8092 -32357 8162 -32347
rect 7762 -32367 7842 -32357
rect 7762 -32427 7772 -32367
rect 7832 -32377 7842 -32367
rect 8082 -32367 8162 -32357
rect 8082 -32377 8092 -32367
rect 7832 -32427 8092 -32377
rect 8152 -32427 8162 -32367
rect 7762 -32437 8162 -32427
rect 8236 -32017 8636 -32007
rect 8236 -32077 8246 -32017
rect 8306 -32067 8566 -32017
rect 8306 -32077 8316 -32067
rect 8236 -32087 8316 -32077
rect 8556 -32077 8566 -32067
rect 8626 -32077 8636 -32017
rect 8556 -32087 8636 -32077
rect 8236 -32357 8296 -32087
rect 8376 -32147 8406 -32127
rect 8356 -32187 8406 -32147
rect 8466 -32147 8496 -32127
rect 8466 -32187 8516 -32147
rect 8356 -32257 8516 -32187
rect 8356 -32297 8406 -32257
rect 8376 -32317 8406 -32297
rect 8466 -32297 8516 -32257
rect 8466 -32317 8496 -32297
rect 8576 -32347 8636 -32087
rect 8566 -32357 8636 -32347
rect 8236 -32367 8316 -32357
rect 8236 -32427 8246 -32367
rect 8306 -32377 8316 -32367
rect 8556 -32367 8636 -32357
rect 8556 -32377 8566 -32367
rect 8306 -32427 8566 -32377
rect 8626 -32427 8636 -32367
rect 8236 -32437 8636 -32427
rect 8692 -32017 9092 -32007
rect 8692 -32077 8702 -32017
rect 8762 -32067 9022 -32017
rect 8762 -32077 8772 -32067
rect 8692 -32087 8772 -32077
rect 9012 -32077 9022 -32067
rect 9082 -32077 9092 -32017
rect 9012 -32087 9092 -32077
rect 8692 -32357 8752 -32087
rect 8832 -32147 8862 -32127
rect 8812 -32187 8862 -32147
rect 8922 -32147 8952 -32127
rect 8922 -32187 8972 -32147
rect 8812 -32257 8972 -32187
rect 8812 -32297 8862 -32257
rect 8832 -32317 8862 -32297
rect 8922 -32297 8972 -32257
rect 8922 -32317 8952 -32297
rect 9032 -32347 9092 -32087
rect 9022 -32357 9092 -32347
rect 8692 -32367 8772 -32357
rect 8692 -32427 8702 -32367
rect 8762 -32377 8772 -32367
rect 9012 -32367 9092 -32357
rect 9012 -32377 9022 -32367
rect 8762 -32427 9022 -32377
rect 9082 -32427 9092 -32367
rect 8692 -32437 9092 -32427
rect 9150 -32017 9550 -32007
rect 9150 -32077 9160 -32017
rect 9220 -32067 9480 -32017
rect 9220 -32077 9230 -32067
rect 9150 -32087 9230 -32077
rect 9470 -32077 9480 -32067
rect 9540 -32077 9550 -32017
rect 9470 -32087 9550 -32077
rect 9150 -32357 9210 -32087
rect 9290 -32147 9320 -32127
rect 9270 -32187 9320 -32147
rect 9380 -32147 9410 -32127
rect 9380 -32187 9430 -32147
rect 9270 -32257 9430 -32187
rect 9270 -32297 9320 -32257
rect 9290 -32317 9320 -32297
rect 9380 -32297 9430 -32257
rect 9380 -32317 9410 -32297
rect 9490 -32347 9550 -32087
rect 9480 -32357 9550 -32347
rect 9150 -32367 9230 -32357
rect 9150 -32427 9160 -32367
rect 9220 -32377 9230 -32367
rect 9470 -32367 9550 -32357
rect 9470 -32377 9480 -32367
rect 9220 -32427 9480 -32377
rect 9540 -32427 9550 -32367
rect 9150 -32437 9550 -32427
rect 9606 -32017 10006 -32007
rect 9606 -32077 9616 -32017
rect 9676 -32067 9936 -32017
rect 9676 -32077 9686 -32067
rect 9606 -32087 9686 -32077
rect 9926 -32077 9936 -32067
rect 9996 -32077 10006 -32017
rect 9926 -32087 10006 -32077
rect 9606 -32357 9666 -32087
rect 9746 -32147 9776 -32127
rect 9726 -32187 9776 -32147
rect 9836 -32147 9866 -32127
rect 9836 -32187 9886 -32147
rect 9726 -32257 9886 -32187
rect 9726 -32297 9776 -32257
rect 9746 -32317 9776 -32297
rect 9836 -32297 9886 -32257
rect 9836 -32317 9866 -32297
rect 9946 -32347 10006 -32087
rect 9936 -32357 10006 -32347
rect 9606 -32367 9686 -32357
rect 9606 -32427 9616 -32367
rect 9676 -32377 9686 -32367
rect 9926 -32367 10006 -32357
rect 9926 -32377 9936 -32367
rect 9676 -32427 9936 -32377
rect 9996 -32427 10006 -32367
rect 9606 -32437 10006 -32427
rect 10062 -32017 10462 -32007
rect 10062 -32077 10072 -32017
rect 10132 -32067 10392 -32017
rect 10132 -32077 10142 -32067
rect 10062 -32087 10142 -32077
rect 10382 -32077 10392 -32067
rect 10452 -32077 10462 -32017
rect 10382 -32087 10462 -32077
rect 10062 -32357 10122 -32087
rect 10202 -32147 10232 -32127
rect 10182 -32187 10232 -32147
rect 10292 -32147 10322 -32127
rect 10292 -32187 10342 -32147
rect 10182 -32257 10342 -32187
rect 10182 -32297 10232 -32257
rect 10202 -32317 10232 -32297
rect 10292 -32297 10342 -32257
rect 10292 -32317 10322 -32297
rect 10402 -32347 10462 -32087
rect 10392 -32357 10462 -32347
rect 10062 -32367 10142 -32357
rect 10062 -32427 10072 -32367
rect 10132 -32377 10142 -32367
rect 10382 -32367 10462 -32357
rect 10382 -32377 10392 -32367
rect 10132 -32427 10392 -32377
rect 10452 -32427 10462 -32367
rect 10062 -32437 10462 -32427
rect 10520 -32017 10920 -32007
rect 10520 -32077 10530 -32017
rect 10590 -32067 10850 -32017
rect 10590 -32077 10600 -32067
rect 10520 -32087 10600 -32077
rect 10840 -32077 10850 -32067
rect 10910 -32077 10920 -32017
rect 10840 -32087 10920 -32077
rect 10520 -32357 10580 -32087
rect 10660 -32147 10690 -32127
rect 10640 -32187 10690 -32147
rect 10750 -32147 10780 -32127
rect 10750 -32187 10800 -32147
rect 10640 -32257 10800 -32187
rect 10640 -32297 10690 -32257
rect 10660 -32317 10690 -32297
rect 10750 -32297 10800 -32257
rect 10750 -32317 10780 -32297
rect 10860 -32347 10920 -32087
rect 10850 -32357 10920 -32347
rect 10520 -32367 10600 -32357
rect 10520 -32427 10530 -32367
rect 10590 -32377 10600 -32367
rect 10840 -32367 10920 -32357
rect 10840 -32377 10850 -32367
rect 10590 -32427 10850 -32377
rect 10910 -32427 10920 -32367
rect 10520 -32437 10920 -32427
rect 10976 -32017 11376 -32007
rect 10976 -32077 10986 -32017
rect 11046 -32067 11306 -32017
rect 11046 -32077 11056 -32067
rect 10976 -32087 11056 -32077
rect 11296 -32077 11306 -32067
rect 11366 -32077 11376 -32017
rect 11296 -32087 11376 -32077
rect 10976 -32357 11036 -32087
rect 11116 -32147 11146 -32127
rect 11096 -32187 11146 -32147
rect 11206 -32147 11236 -32127
rect 11206 -32187 11256 -32147
rect 11096 -32257 11256 -32187
rect 11096 -32297 11146 -32257
rect 11116 -32317 11146 -32297
rect 11206 -32297 11256 -32257
rect 11206 -32317 11236 -32297
rect 11316 -32347 11376 -32087
rect 11306 -32357 11376 -32347
rect 10976 -32367 11056 -32357
rect 10976 -32427 10986 -32367
rect 11046 -32377 11056 -32367
rect 11296 -32367 11376 -32357
rect 11296 -32377 11306 -32367
rect 11046 -32427 11306 -32377
rect 11366 -32427 11376 -32367
rect 10976 -32437 11376 -32427
rect 11432 -32017 11832 -32007
rect 11432 -32077 11442 -32017
rect 11502 -32067 11762 -32017
rect 11502 -32077 11512 -32067
rect 11432 -32087 11512 -32077
rect 11752 -32077 11762 -32067
rect 11822 -32077 11832 -32017
rect 11752 -32087 11832 -32077
rect 11432 -32357 11492 -32087
rect 11572 -32147 11602 -32127
rect 11552 -32187 11602 -32147
rect 11662 -32147 11692 -32127
rect 11662 -32187 11712 -32147
rect 11552 -32257 11712 -32187
rect 11552 -32297 11602 -32257
rect 11572 -32317 11602 -32297
rect 11662 -32297 11712 -32257
rect 11662 -32317 11692 -32297
rect 11772 -32347 11832 -32087
rect 11762 -32357 11832 -32347
rect 11432 -32367 11512 -32357
rect 11432 -32427 11442 -32367
rect 11502 -32377 11512 -32367
rect 11752 -32367 11832 -32357
rect 11752 -32377 11762 -32367
rect 11502 -32427 11762 -32377
rect 11822 -32427 11832 -32367
rect 11432 -32437 11832 -32427
rect 11890 -32017 12290 -32007
rect 11890 -32077 11900 -32017
rect 11960 -32067 12220 -32017
rect 11960 -32077 11970 -32067
rect 11890 -32087 11970 -32077
rect 12210 -32077 12220 -32067
rect 12280 -32077 12290 -32017
rect 12210 -32087 12290 -32077
rect 11890 -32357 11950 -32087
rect 12030 -32147 12060 -32127
rect 12010 -32187 12060 -32147
rect 12120 -32147 12150 -32127
rect 12120 -32187 12170 -32147
rect 12010 -32257 12170 -32187
rect 12010 -32297 12060 -32257
rect 12030 -32317 12060 -32297
rect 12120 -32297 12170 -32257
rect 12120 -32317 12150 -32297
rect 12230 -32347 12290 -32087
rect 12220 -32357 12290 -32347
rect 11890 -32367 11970 -32357
rect 11890 -32427 11900 -32367
rect 11960 -32377 11970 -32367
rect 12210 -32367 12290 -32357
rect 12210 -32377 12220 -32367
rect 11960 -32427 12220 -32377
rect 12280 -32427 12290 -32367
rect 11890 -32437 12290 -32427
rect 12346 -32017 12746 -32007
rect 12346 -32077 12356 -32017
rect 12416 -32067 12676 -32017
rect 12416 -32077 12426 -32067
rect 12346 -32087 12426 -32077
rect 12666 -32077 12676 -32067
rect 12736 -32077 12746 -32017
rect 12666 -32087 12746 -32077
rect 12346 -32357 12406 -32087
rect 12486 -32147 12516 -32127
rect 12466 -32187 12516 -32147
rect 12576 -32147 12606 -32127
rect 12576 -32187 12626 -32147
rect 12466 -32257 12626 -32187
rect 12466 -32297 12516 -32257
rect 12486 -32317 12516 -32297
rect 12576 -32297 12626 -32257
rect 12576 -32317 12606 -32297
rect 12686 -32347 12746 -32087
rect 12676 -32357 12746 -32347
rect 12346 -32367 12426 -32357
rect 12346 -32427 12356 -32367
rect 12416 -32377 12426 -32367
rect 12666 -32367 12746 -32357
rect 12666 -32377 12676 -32367
rect 12416 -32427 12676 -32377
rect 12736 -32427 12746 -32367
rect 12346 -32437 12746 -32427
rect 12802 -32017 13202 -32007
rect 12802 -32077 12812 -32017
rect 12872 -32067 13132 -32017
rect 12872 -32077 12882 -32067
rect 12802 -32087 12882 -32077
rect 13122 -32077 13132 -32067
rect 13192 -32077 13202 -32017
rect 13122 -32087 13202 -32077
rect 12802 -32357 12862 -32087
rect 12942 -32147 12972 -32127
rect 12922 -32187 12972 -32147
rect 13032 -32147 13062 -32127
rect 13032 -32187 13082 -32147
rect 12922 -32257 13082 -32187
rect 12922 -32297 12972 -32257
rect 12942 -32317 12972 -32297
rect 13032 -32297 13082 -32257
rect 13032 -32317 13062 -32297
rect 13142 -32347 13202 -32087
rect 13132 -32357 13202 -32347
rect 12802 -32367 12882 -32357
rect 12802 -32427 12812 -32367
rect 12872 -32377 12882 -32367
rect 13122 -32367 13202 -32357
rect 13122 -32377 13132 -32367
rect 12872 -32427 13132 -32377
rect 13192 -32427 13202 -32367
rect 12802 -32437 13202 -32427
rect 13260 -32017 13660 -32007
rect 13260 -32077 13270 -32017
rect 13330 -32067 13590 -32017
rect 13330 -32077 13340 -32067
rect 13260 -32087 13340 -32077
rect 13580 -32077 13590 -32067
rect 13650 -32077 13660 -32017
rect 13580 -32087 13660 -32077
rect 13260 -32357 13320 -32087
rect 13400 -32147 13430 -32127
rect 13380 -32187 13430 -32147
rect 13490 -32147 13520 -32127
rect 13490 -32187 13540 -32147
rect 13380 -32257 13540 -32187
rect 13380 -32297 13430 -32257
rect 13400 -32317 13430 -32297
rect 13490 -32297 13540 -32257
rect 13490 -32317 13520 -32297
rect 13600 -32347 13660 -32087
rect 13590 -32357 13660 -32347
rect 13260 -32367 13340 -32357
rect 13260 -32427 13270 -32367
rect 13330 -32377 13340 -32367
rect 13580 -32367 13660 -32357
rect 13580 -32377 13590 -32367
rect 13330 -32427 13590 -32377
rect 13650 -32427 13660 -32367
rect 13260 -32437 13660 -32427
rect 13716 -32017 14116 -32007
rect 13716 -32077 13726 -32017
rect 13786 -32067 14046 -32017
rect 13786 -32077 13796 -32067
rect 13716 -32087 13796 -32077
rect 14036 -32077 14046 -32067
rect 14106 -32077 14116 -32017
rect 14036 -32087 14116 -32077
rect 13716 -32357 13776 -32087
rect 13856 -32147 13886 -32127
rect 13836 -32187 13886 -32147
rect 13946 -32147 13976 -32127
rect 13946 -32187 13996 -32147
rect 13836 -32257 13996 -32187
rect 13836 -32297 13886 -32257
rect 13856 -32317 13886 -32297
rect 13946 -32297 13996 -32257
rect 13946 -32317 13976 -32297
rect 14056 -32347 14116 -32087
rect 14046 -32357 14116 -32347
rect 13716 -32367 13796 -32357
rect 13716 -32427 13726 -32367
rect 13786 -32377 13796 -32367
rect 14036 -32367 14116 -32357
rect 14036 -32377 14046 -32367
rect 13786 -32427 14046 -32377
rect 14106 -32427 14116 -32367
rect 13716 -32437 14116 -32427
rect 14172 -32017 14572 -32007
rect 14172 -32077 14182 -32017
rect 14242 -32067 14502 -32017
rect 14242 -32077 14252 -32067
rect 14172 -32087 14252 -32077
rect 14492 -32077 14502 -32067
rect 14562 -32077 14572 -32017
rect 14492 -32087 14572 -32077
rect 14172 -32357 14232 -32087
rect 14312 -32147 14342 -32127
rect 14292 -32187 14342 -32147
rect 14402 -32147 14432 -32127
rect 14402 -32187 14452 -32147
rect 14292 -32257 14452 -32187
rect 14292 -32297 14342 -32257
rect 14312 -32317 14342 -32297
rect 14402 -32297 14452 -32257
rect 14402 -32317 14432 -32297
rect 14512 -32347 14572 -32087
rect 14502 -32357 14572 -32347
rect 14172 -32367 14252 -32357
rect 14172 -32427 14182 -32367
rect 14242 -32377 14252 -32367
rect 14492 -32367 14572 -32357
rect 14492 -32377 14502 -32367
rect 14242 -32427 14502 -32377
rect 14562 -32427 14572 -32367
rect 14172 -32437 14572 -32427
rect 14630 -32017 15030 -32007
rect 14630 -32077 14640 -32017
rect 14700 -32067 14960 -32017
rect 14700 -32077 14710 -32067
rect 14630 -32087 14710 -32077
rect 14950 -32077 14960 -32067
rect 15020 -32077 15030 -32017
rect 14950 -32087 15030 -32077
rect 14630 -32357 14690 -32087
rect 14770 -32147 14800 -32127
rect 14750 -32187 14800 -32147
rect 14860 -32147 14890 -32127
rect 14860 -32187 14910 -32147
rect 14750 -32257 14910 -32187
rect 14750 -32297 14800 -32257
rect 14770 -32317 14800 -32297
rect 14860 -32297 14910 -32257
rect 14860 -32317 14890 -32297
rect 14970 -32347 15030 -32087
rect 14960 -32357 15030 -32347
rect 14630 -32367 14710 -32357
rect 14630 -32427 14640 -32367
rect 14700 -32377 14710 -32367
rect 14950 -32367 15030 -32357
rect 14950 -32377 14960 -32367
rect 14700 -32427 14960 -32377
rect 15020 -32427 15030 -32367
rect 14630 -32437 15030 -32427
rect 15086 -32017 15486 -32007
rect 15086 -32077 15096 -32017
rect 15156 -32067 15416 -32017
rect 15156 -32077 15166 -32067
rect 15086 -32087 15166 -32077
rect 15406 -32077 15416 -32067
rect 15476 -32077 15486 -32017
rect 15406 -32087 15486 -32077
rect 15086 -32357 15146 -32087
rect 15226 -32147 15256 -32127
rect 15206 -32187 15256 -32147
rect 15316 -32147 15346 -32127
rect 15316 -32187 15366 -32147
rect 15206 -32257 15366 -32187
rect 15206 -32297 15256 -32257
rect 15226 -32317 15256 -32297
rect 15316 -32297 15366 -32257
rect 15316 -32317 15346 -32297
rect 15426 -32347 15486 -32087
rect 15416 -32357 15486 -32347
rect 15086 -32367 15166 -32357
rect 15086 -32427 15096 -32367
rect 15156 -32377 15166 -32367
rect 15406 -32367 15486 -32357
rect 15406 -32377 15416 -32367
rect 15156 -32427 15416 -32377
rect 15476 -32427 15486 -32367
rect 15086 -32437 15486 -32427
<< via3 >>
rect 89 590 150 651
rect 250 590 311 651
rect 15127 551 15201 611
rect 15358 551 15432 611
rect 1540 270 1600 330
rect 1540 140 1600 200
rect 1996 270 2056 330
rect 1996 140 2056 200
rect 2452 270 2512 330
rect 2452 140 2512 200
rect 2910 270 2970 330
rect 2910 140 2970 200
rect 3366 270 3426 330
rect 3366 140 3426 200
rect 3822 270 3882 330
rect 3822 140 3882 200
rect 4280 270 4340 330
rect 4280 140 4340 200
rect 4736 270 4796 330
rect 4736 140 4796 200
rect 5192 270 5252 330
rect 5192 140 5252 200
rect 5650 270 5710 330
rect 5650 140 5710 200
rect 6106 270 6166 330
rect 6106 140 6166 200
rect 6562 270 6622 330
rect 6562 140 6622 200
rect 7020 270 7080 330
rect 7020 140 7080 200
rect 7476 270 7536 330
rect 7476 140 7536 200
rect 7932 270 7992 330
rect 7932 140 7992 200
rect 8406 270 8466 330
rect 8406 140 8466 200
rect 8862 270 8922 330
rect 8862 140 8922 200
rect 9320 270 9380 330
rect 9320 140 9380 200
rect 9776 270 9836 330
rect 9776 140 9836 200
rect 10232 270 10292 330
rect 10232 140 10292 200
rect 10690 270 10750 330
rect 10690 140 10750 200
rect 11146 270 11206 330
rect 11146 140 11206 200
rect 11602 270 11662 330
rect 11602 140 11662 200
rect 12060 270 12120 330
rect 12060 140 12120 200
rect 12516 270 12576 330
rect 12516 140 12576 200
rect 12972 270 13032 330
rect 12972 140 13032 200
rect 13430 270 13490 330
rect 13430 140 13490 200
rect 13886 270 13946 330
rect 13886 140 13946 200
rect 14342 270 14402 330
rect 14342 140 14402 200
rect 14800 270 14860 330
rect 14800 140 14860 200
rect 15256 270 15316 330
rect 15256 140 15316 200
rect 170 -222 230 -162
rect 170 -352 230 -292
rect 626 -222 686 -162
rect 626 -352 686 -292
rect 1082 -222 1142 -162
rect 1082 -352 1142 -292
rect 1540 -222 1600 -162
rect 1540 -352 1600 -292
rect 1996 -222 2056 -162
rect 1996 -352 2056 -292
rect 2452 -222 2512 -162
rect 2452 -352 2512 -292
rect 2910 -222 2970 -162
rect 2910 -352 2970 -292
rect 3366 -222 3426 -162
rect 3366 -352 3426 -292
rect 3822 -222 3882 -162
rect 3822 -352 3882 -292
rect 4280 -222 4340 -162
rect 4280 -352 4340 -292
rect 4736 -222 4796 -162
rect 4736 -352 4796 -292
rect 5192 -222 5252 -162
rect 5192 -352 5252 -292
rect 5650 -222 5710 -162
rect 5650 -352 5710 -292
rect 6106 -222 6166 -162
rect 6106 -352 6166 -292
rect 6562 -222 6622 -162
rect 6562 -352 6622 -292
rect 7020 -222 7080 -162
rect 7020 -352 7080 -292
rect 7476 -222 7536 -162
rect 7476 -352 7536 -292
rect 7932 -222 7992 -162
rect 7932 -352 7992 -292
rect 8406 -222 8466 -162
rect 8406 -352 8466 -292
rect 8862 -222 8922 -162
rect 8862 -352 8922 -292
rect 9320 -222 9380 -162
rect 9320 -352 9380 -292
rect 9776 -222 9836 -162
rect 9776 -352 9836 -292
rect 10232 -222 10292 -162
rect 10232 -352 10292 -292
rect 10690 -222 10750 -162
rect 10690 -352 10750 -292
rect 11146 -222 11206 -162
rect 11146 -352 11206 -292
rect 11602 -222 11662 -162
rect 11602 -352 11662 -292
rect 12060 -222 12120 -162
rect 12060 -352 12120 -292
rect 12516 -222 12576 -162
rect 12516 -352 12576 -292
rect 12972 -222 13032 -162
rect 12972 -352 13032 -292
rect 13430 -222 13490 -162
rect 13430 -352 13490 -292
rect 13886 -222 13946 -162
rect 13886 -352 13946 -292
rect 14342 -222 14402 -162
rect 14342 -352 14402 -292
rect 14800 -222 14860 -162
rect 14800 -352 14860 -292
rect 15256 -222 15316 -162
rect 15256 -352 15316 -292
rect 170 -724 230 -664
rect 170 -854 230 -794
rect 626 -724 686 -664
rect 626 -854 686 -794
rect 1082 -724 1142 -664
rect 1082 -854 1142 -794
rect 1540 -724 1600 -664
rect 1540 -854 1600 -794
rect 1996 -724 2056 -664
rect 1996 -854 2056 -794
rect 2452 -724 2512 -664
rect 2452 -854 2512 -794
rect 2910 -724 2970 -664
rect 2910 -854 2970 -794
rect 3366 -724 3426 -664
rect 3366 -854 3426 -794
rect 3822 -724 3882 -664
rect 3822 -854 3882 -794
rect 4280 -724 4340 -664
rect 4280 -854 4340 -794
rect 4736 -724 4796 -664
rect 4736 -854 4796 -794
rect 5192 -724 5252 -664
rect 5192 -854 5252 -794
rect 5650 -724 5710 -664
rect 5650 -854 5710 -794
rect 6106 -724 6166 -664
rect 6106 -854 6166 -794
rect 6562 -724 6622 -664
rect 6562 -854 6622 -794
rect 7020 -724 7080 -664
rect 7020 -854 7080 -794
rect 7476 -724 7536 -664
rect 7476 -854 7536 -794
rect 7932 -724 7992 -664
rect 7932 -854 7992 -794
rect 8406 -724 8466 -664
rect 8406 -854 8466 -794
rect 8862 -724 8922 -664
rect 8862 -854 8922 -794
rect 9320 -724 9380 -664
rect 9320 -854 9380 -794
rect 9776 -724 9836 -664
rect 9776 -854 9836 -794
rect 10232 -724 10292 -664
rect 10232 -854 10292 -794
rect 10690 -724 10750 -664
rect 10690 -854 10750 -794
rect 11146 -724 11206 -664
rect 11146 -854 11206 -794
rect 11602 -724 11662 -664
rect 11602 -854 11662 -794
rect 12060 -724 12120 -664
rect 12060 -854 12120 -794
rect 12516 -724 12576 -664
rect 12516 -854 12576 -794
rect 12972 -724 13032 -664
rect 12972 -854 13032 -794
rect 13430 -724 13490 -664
rect 13430 -854 13490 -794
rect 13886 -724 13946 -664
rect 13886 -854 13946 -794
rect 14342 -724 14402 -664
rect 14342 -854 14402 -794
rect 14800 -724 14860 -664
rect 14800 -854 14860 -794
rect 15256 -724 15316 -664
rect 15256 -854 15316 -794
rect 170 -1216 230 -1156
rect 170 -1346 230 -1286
rect 626 -1216 686 -1156
rect 626 -1346 686 -1286
rect 1082 -1216 1142 -1156
rect 1082 -1346 1142 -1286
rect 1540 -1216 1600 -1156
rect 1540 -1346 1600 -1286
rect 1996 -1216 2056 -1156
rect 1996 -1346 2056 -1286
rect 2452 -1216 2512 -1156
rect 2452 -1346 2512 -1286
rect 2910 -1216 2970 -1156
rect 2910 -1346 2970 -1286
rect 3366 -1216 3426 -1156
rect 3366 -1346 3426 -1286
rect 3822 -1216 3882 -1156
rect 3822 -1346 3882 -1286
rect 4280 -1216 4340 -1156
rect 4280 -1346 4340 -1286
rect 4736 -1216 4796 -1156
rect 4736 -1346 4796 -1286
rect 5192 -1216 5252 -1156
rect 5192 -1346 5252 -1286
rect 5650 -1216 5710 -1156
rect 5650 -1346 5710 -1286
rect 6106 -1216 6166 -1156
rect 6106 -1346 6166 -1286
rect 6562 -1216 6622 -1156
rect 6562 -1346 6622 -1286
rect 7020 -1216 7080 -1156
rect 7020 -1346 7080 -1286
rect 7476 -1216 7536 -1156
rect 7476 -1346 7536 -1286
rect 7932 -1216 7992 -1156
rect 7932 -1346 7992 -1286
rect 8406 -1216 8466 -1156
rect 8406 -1346 8466 -1286
rect 8862 -1216 8922 -1156
rect 8862 -1346 8922 -1286
rect 9320 -1216 9380 -1156
rect 9320 -1346 9380 -1286
rect 9776 -1216 9836 -1156
rect 9776 -1346 9836 -1286
rect 10232 -1216 10292 -1156
rect 10232 -1346 10292 -1286
rect 10690 -1216 10750 -1156
rect 10690 -1346 10750 -1286
rect 11146 -1216 11206 -1156
rect 11146 -1346 11206 -1286
rect 11602 -1216 11662 -1156
rect 11602 -1346 11662 -1286
rect 12060 -1216 12120 -1156
rect 12060 -1346 12120 -1286
rect 12516 -1216 12576 -1156
rect 12516 -1346 12576 -1286
rect 12972 -1216 13032 -1156
rect 12972 -1346 13032 -1286
rect 13430 -1216 13490 -1156
rect 13430 -1346 13490 -1286
rect 13886 -1216 13946 -1156
rect 13886 -1346 13946 -1286
rect 14342 -1216 14402 -1156
rect 14342 -1346 14402 -1286
rect 14800 -1216 14860 -1156
rect 14800 -1346 14860 -1286
rect 15256 -1216 15316 -1156
rect 15256 -1346 15316 -1286
rect 170 -1732 230 -1672
rect 170 -1862 230 -1802
rect 626 -1732 686 -1672
rect 626 -1862 686 -1802
rect 1082 -1732 1142 -1672
rect 1082 -1862 1142 -1802
rect 1540 -1732 1600 -1672
rect 1540 -1862 1600 -1802
rect 1996 -1732 2056 -1672
rect 1996 -1862 2056 -1802
rect 2452 -1732 2512 -1672
rect 2452 -1862 2512 -1802
rect 2910 -1732 2970 -1672
rect 2910 -1862 2970 -1802
rect 3366 -1732 3426 -1672
rect 3366 -1862 3426 -1802
rect 3822 -1732 3882 -1672
rect 3822 -1862 3882 -1802
rect 4280 -1732 4340 -1672
rect 4280 -1862 4340 -1802
rect 4736 -1732 4796 -1672
rect 4736 -1862 4796 -1802
rect 5192 -1732 5252 -1672
rect 5192 -1862 5252 -1802
rect 5650 -1732 5710 -1672
rect 5650 -1862 5710 -1802
rect 6106 -1732 6166 -1672
rect 6106 -1862 6166 -1802
rect 6562 -1732 6622 -1672
rect 6562 -1862 6622 -1802
rect 7020 -1732 7080 -1672
rect 7020 -1862 7080 -1802
rect 7476 -1732 7536 -1672
rect 7476 -1862 7536 -1802
rect 7932 -1732 7992 -1672
rect 7932 -1862 7992 -1802
rect 8406 -1732 8466 -1672
rect 8406 -1862 8466 -1802
rect 8862 -1732 8922 -1672
rect 8862 -1862 8922 -1802
rect 9320 -1732 9380 -1672
rect 9320 -1862 9380 -1802
rect 9776 -1732 9836 -1672
rect 9776 -1862 9836 -1802
rect 10232 -1732 10292 -1672
rect 10232 -1862 10292 -1802
rect 10690 -1732 10750 -1672
rect 10690 -1862 10750 -1802
rect 11146 -1732 11206 -1672
rect 11146 -1862 11206 -1802
rect 11602 -1732 11662 -1672
rect 11602 -1862 11662 -1802
rect 12060 -1732 12120 -1672
rect 12060 -1862 12120 -1802
rect 12516 -1732 12576 -1672
rect 12516 -1862 12576 -1802
rect 12972 -1732 13032 -1672
rect 12972 -1862 13032 -1802
rect 13430 -1732 13490 -1672
rect 13430 -1862 13490 -1802
rect 13886 -1732 13946 -1672
rect 13886 -1862 13946 -1802
rect 14342 -1732 14402 -1672
rect 14342 -1862 14402 -1802
rect 14800 -1732 14860 -1672
rect 14800 -1862 14860 -1802
rect 15256 -1732 15316 -1672
rect 15256 -1862 15316 -1802
rect 170 -2234 230 -2174
rect 170 -2364 230 -2304
rect 626 -2234 686 -2174
rect 626 -2364 686 -2304
rect 1082 -2234 1142 -2174
rect 1082 -2364 1142 -2304
rect 1540 -2234 1600 -2174
rect 1540 -2364 1600 -2304
rect 1996 -2234 2056 -2174
rect 1996 -2364 2056 -2304
rect 2452 -2234 2512 -2174
rect 2452 -2364 2512 -2304
rect 2910 -2234 2970 -2174
rect 2910 -2364 2970 -2304
rect 3366 -2234 3426 -2174
rect 3366 -2364 3426 -2304
rect 3822 -2234 3882 -2174
rect 3822 -2364 3882 -2304
rect 4280 -2234 4340 -2174
rect 4280 -2364 4340 -2304
rect 4736 -2234 4796 -2174
rect 4736 -2364 4796 -2304
rect 5192 -2234 5252 -2174
rect 5192 -2364 5252 -2304
rect 5650 -2234 5710 -2174
rect 5650 -2364 5710 -2304
rect 6106 -2234 6166 -2174
rect 6106 -2364 6166 -2304
rect 6562 -2234 6622 -2174
rect 6562 -2364 6622 -2304
rect 7020 -2234 7080 -2174
rect 7020 -2364 7080 -2304
rect 7476 -2234 7536 -2174
rect 7476 -2364 7536 -2304
rect 7932 -2234 7992 -2174
rect 7932 -2364 7992 -2304
rect 8406 -2234 8466 -2174
rect 8406 -2364 8466 -2304
rect 8862 -2234 8922 -2174
rect 8862 -2364 8922 -2304
rect 9320 -2234 9380 -2174
rect 9320 -2364 9380 -2304
rect 9776 -2234 9836 -2174
rect 9776 -2364 9836 -2304
rect 10232 -2234 10292 -2174
rect 10232 -2364 10292 -2304
rect 10690 -2234 10750 -2174
rect 10690 -2364 10750 -2304
rect 11146 -2234 11206 -2174
rect 11146 -2364 11206 -2304
rect 11602 -2234 11662 -2174
rect 11602 -2364 11662 -2304
rect 12060 -2234 12120 -2174
rect 12060 -2364 12120 -2304
rect 12516 -2234 12576 -2174
rect 12516 -2364 12576 -2304
rect 12972 -2234 13032 -2174
rect 12972 -2364 13032 -2304
rect 13430 -2234 13490 -2174
rect 13430 -2364 13490 -2304
rect 13886 -2234 13946 -2174
rect 13886 -2364 13946 -2304
rect 14342 -2234 14402 -2174
rect 14342 -2364 14402 -2304
rect 14800 -2234 14860 -2174
rect 14800 -2364 14860 -2304
rect 15256 -2234 15316 -2174
rect 15256 -2364 15316 -2304
rect 170 -2726 230 -2666
rect 170 -2856 230 -2796
rect 626 -2726 686 -2666
rect 626 -2856 686 -2796
rect 1082 -2726 1142 -2666
rect 1082 -2856 1142 -2796
rect 1540 -2726 1600 -2666
rect 1540 -2856 1600 -2796
rect 1996 -2726 2056 -2666
rect 1996 -2856 2056 -2796
rect 2452 -2726 2512 -2666
rect 2452 -2856 2512 -2796
rect 2910 -2726 2970 -2666
rect 2910 -2856 2970 -2796
rect 3366 -2726 3426 -2666
rect 3366 -2856 3426 -2796
rect 3822 -2726 3882 -2666
rect 3822 -2856 3882 -2796
rect 4280 -2726 4340 -2666
rect 4280 -2856 4340 -2796
rect 4736 -2726 4796 -2666
rect 4736 -2856 4796 -2796
rect 5192 -2726 5252 -2666
rect 5192 -2856 5252 -2796
rect 5650 -2726 5710 -2666
rect 5650 -2856 5710 -2796
rect 6106 -2726 6166 -2666
rect 6106 -2856 6166 -2796
rect 6562 -2726 6622 -2666
rect 6562 -2856 6622 -2796
rect 7020 -2726 7080 -2666
rect 7020 -2856 7080 -2796
rect 7476 -2726 7536 -2666
rect 7476 -2856 7536 -2796
rect 7932 -2726 7992 -2666
rect 7932 -2856 7992 -2796
rect 8406 -2726 8466 -2666
rect 8406 -2856 8466 -2796
rect 8862 -2726 8922 -2666
rect 8862 -2856 8922 -2796
rect 9320 -2726 9380 -2666
rect 9320 -2856 9380 -2796
rect 9776 -2726 9836 -2666
rect 9776 -2856 9836 -2796
rect 10232 -2726 10292 -2666
rect 10232 -2856 10292 -2796
rect 10690 -2726 10750 -2666
rect 10690 -2856 10750 -2796
rect 11146 -2726 11206 -2666
rect 11146 -2856 11206 -2796
rect 11602 -2726 11662 -2666
rect 11602 -2856 11662 -2796
rect 12060 -2726 12120 -2666
rect 12060 -2856 12120 -2796
rect 12516 -2726 12576 -2666
rect 12516 -2856 12576 -2796
rect 12972 -2726 13032 -2666
rect 12972 -2856 13032 -2796
rect 13430 -2726 13490 -2666
rect 13430 -2856 13490 -2796
rect 13886 -2726 13946 -2666
rect 13886 -2856 13946 -2796
rect 14342 -2726 14402 -2666
rect 14342 -2856 14402 -2796
rect 14800 -2726 14860 -2666
rect 14800 -2856 14860 -2796
rect 15256 -2726 15316 -2666
rect 15256 -2856 15316 -2796
rect 170 -3722 230 -3662
rect 170 -3852 230 -3792
rect 626 -3722 686 -3662
rect 626 -3852 686 -3792
rect 1082 -3722 1142 -3662
rect 1082 -3852 1142 -3792
rect 1540 -3722 1600 -3662
rect 1540 -3852 1600 -3792
rect 1996 -3722 2056 -3662
rect 1996 -3852 2056 -3792
rect 2452 -3722 2512 -3662
rect 2452 -3852 2512 -3792
rect 2910 -3722 2970 -3662
rect 2910 -3852 2970 -3792
rect 3366 -3722 3426 -3662
rect 3366 -3852 3426 -3792
rect 3822 -3722 3882 -3662
rect 3822 -3852 3882 -3792
rect 4280 -3722 4340 -3662
rect 4280 -3852 4340 -3792
rect 4736 -3722 4796 -3662
rect 4736 -3852 4796 -3792
rect 5192 -3722 5252 -3662
rect 5192 -3852 5252 -3792
rect 5650 -3722 5710 -3662
rect 5650 -3852 5710 -3792
rect 6106 -3722 6166 -3662
rect 6106 -3852 6166 -3792
rect 6562 -3722 6622 -3662
rect 6562 -3852 6622 -3792
rect 7020 -3722 7080 -3662
rect 7020 -3852 7080 -3792
rect 7476 -3722 7536 -3662
rect 7476 -3852 7536 -3792
rect 7932 -3722 7992 -3662
rect 7932 -3852 7992 -3792
rect 8406 -3722 8466 -3662
rect 8406 -3852 8466 -3792
rect 8862 -3722 8922 -3662
rect 8862 -3852 8922 -3792
rect 9320 -3722 9380 -3662
rect 9320 -3852 9380 -3792
rect 9776 -3722 9836 -3662
rect 9776 -3852 9836 -3792
rect 10232 -3722 10292 -3662
rect 10232 -3852 10292 -3792
rect 10690 -3722 10750 -3662
rect 10690 -3852 10750 -3792
rect 11146 -3722 11206 -3662
rect 11146 -3852 11206 -3792
rect 11602 -3722 11662 -3662
rect 11602 -3852 11662 -3792
rect 12060 -3722 12120 -3662
rect 12060 -3852 12120 -3792
rect 12516 -3722 12576 -3662
rect 12516 -3852 12576 -3792
rect 12972 -3722 13032 -3662
rect 12972 -3852 13032 -3792
rect 13430 -3722 13490 -3662
rect 13430 -3852 13490 -3792
rect 13886 -3722 13946 -3662
rect 13886 -3852 13946 -3792
rect 14342 -3722 14402 -3662
rect 14342 -3852 14402 -3792
rect 14800 -3722 14860 -3662
rect 14800 -3852 14860 -3792
rect 15256 -3722 15316 -3662
rect 15256 -3852 15316 -3792
rect 170 -4214 230 -4154
rect 170 -4344 230 -4284
rect 626 -4214 686 -4154
rect 626 -4344 686 -4284
rect 1082 -4214 1142 -4154
rect 1082 -4344 1142 -4284
rect 1540 -4214 1600 -4154
rect 1540 -4344 1600 -4284
rect 1996 -4214 2056 -4154
rect 1996 -4344 2056 -4284
rect 2452 -4214 2512 -4154
rect 2452 -4344 2512 -4284
rect 2910 -4214 2970 -4154
rect 2910 -4344 2970 -4284
rect 3366 -4214 3426 -4154
rect 3366 -4344 3426 -4284
rect 3822 -4214 3882 -4154
rect 3822 -4344 3882 -4284
rect 4280 -4214 4340 -4154
rect 4280 -4344 4340 -4284
rect 4736 -4214 4796 -4154
rect 4736 -4344 4796 -4284
rect 5192 -4214 5252 -4154
rect 5192 -4344 5252 -4284
rect 5650 -4214 5710 -4154
rect 5650 -4344 5710 -4284
rect 6106 -4214 6166 -4154
rect 6106 -4344 6166 -4284
rect 6562 -4214 6622 -4154
rect 6562 -4344 6622 -4284
rect 7020 -4214 7080 -4154
rect 7020 -4344 7080 -4284
rect 7476 -4214 7536 -4154
rect 7476 -4344 7536 -4284
rect 7932 -4214 7992 -4154
rect 7932 -4344 7992 -4284
rect 8406 -4214 8466 -4154
rect 8406 -4344 8466 -4284
rect 8862 -4214 8922 -4154
rect 8862 -4344 8922 -4284
rect 9320 -4214 9380 -4154
rect 9320 -4344 9380 -4284
rect 9776 -4214 9836 -4154
rect 9776 -4344 9836 -4284
rect 10232 -4214 10292 -4154
rect 10232 -4344 10292 -4284
rect 10690 -4214 10750 -4154
rect 10690 -4344 10750 -4284
rect 11146 -4214 11206 -4154
rect 11146 -4344 11206 -4284
rect 11602 -4214 11662 -4154
rect 11602 -4344 11662 -4284
rect 12060 -4214 12120 -4154
rect 12060 -4344 12120 -4284
rect 12516 -4214 12576 -4154
rect 12516 -4344 12576 -4284
rect 12972 -4214 13032 -4154
rect 12972 -4344 13032 -4284
rect 13430 -4214 13490 -4154
rect 13430 -4344 13490 -4284
rect 13886 -4214 13946 -4154
rect 13886 -4344 13946 -4284
rect 14342 -4214 14402 -4154
rect 14342 -4344 14402 -4284
rect 14800 -4214 14860 -4154
rect 14800 -4344 14860 -4284
rect 15256 -4214 15316 -4154
rect 15256 -4344 15316 -4284
rect 170 -4730 230 -4670
rect 170 -4860 230 -4800
rect 626 -4730 686 -4670
rect 626 -4860 686 -4800
rect 1082 -4730 1142 -4670
rect 1082 -4860 1142 -4800
rect 1540 -4730 1600 -4670
rect 1540 -4860 1600 -4800
rect 1996 -4730 2056 -4670
rect 1996 -4860 2056 -4800
rect 2452 -4730 2512 -4670
rect 2452 -4860 2512 -4800
rect 2910 -4730 2970 -4670
rect 2910 -4860 2970 -4800
rect 3366 -4730 3426 -4670
rect 3366 -4860 3426 -4800
rect 3822 -4730 3882 -4670
rect 3822 -4860 3882 -4800
rect 4280 -4730 4340 -4670
rect 4280 -4860 4340 -4800
rect 4736 -4730 4796 -4670
rect 4736 -4860 4796 -4800
rect 5192 -4730 5252 -4670
rect 5192 -4860 5252 -4800
rect 5650 -4730 5710 -4670
rect 5650 -4860 5710 -4800
rect 6106 -4730 6166 -4670
rect 6106 -4860 6166 -4800
rect 6562 -4730 6622 -4670
rect 6562 -4860 6622 -4800
rect 7020 -4730 7080 -4670
rect 7020 -4860 7080 -4800
rect 7476 -4730 7536 -4670
rect 7476 -4860 7536 -4800
rect 7932 -4730 7992 -4670
rect 7932 -4860 7992 -4800
rect 8406 -4730 8466 -4670
rect 8406 -4860 8466 -4800
rect 8862 -4730 8922 -4670
rect 8862 -4860 8922 -4800
rect 9320 -4730 9380 -4670
rect 9320 -4860 9380 -4800
rect 9776 -4730 9836 -4670
rect 9776 -4860 9836 -4800
rect 10232 -4730 10292 -4670
rect 10232 -4860 10292 -4800
rect 10690 -4730 10750 -4670
rect 10690 -4860 10750 -4800
rect 11146 -4730 11206 -4670
rect 11146 -4860 11206 -4800
rect 11602 -4730 11662 -4670
rect 11602 -4860 11662 -4800
rect 12060 -4730 12120 -4670
rect 12060 -4860 12120 -4800
rect 12516 -4730 12576 -4670
rect 12516 -4860 12576 -4800
rect 12972 -4730 13032 -4670
rect 12972 -4860 13032 -4800
rect 13430 -4730 13490 -4670
rect 13430 -4860 13490 -4800
rect 13886 -4730 13946 -4670
rect 13886 -4860 13946 -4800
rect 14342 -4730 14402 -4670
rect 14342 -4860 14402 -4800
rect 14800 -4730 14860 -4670
rect 14800 -4860 14860 -4800
rect 15256 -4730 15316 -4670
rect 15256 -4860 15316 -4800
rect 170 -5232 230 -5172
rect 170 -5362 230 -5302
rect 626 -5232 686 -5172
rect 626 -5362 686 -5302
rect 1082 -5232 1142 -5172
rect 1082 -5362 1142 -5302
rect 1540 -5232 1600 -5172
rect 1540 -5362 1600 -5302
rect 1996 -5232 2056 -5172
rect 1996 -5362 2056 -5302
rect 2452 -5232 2512 -5172
rect 2452 -5362 2512 -5302
rect 2910 -5232 2970 -5172
rect 2910 -5362 2970 -5302
rect 3366 -5232 3426 -5172
rect 3366 -5362 3426 -5302
rect 3822 -5232 3882 -5172
rect 3822 -5362 3882 -5302
rect 4280 -5232 4340 -5172
rect 4280 -5362 4340 -5302
rect 4736 -5232 4796 -5172
rect 4736 -5362 4796 -5302
rect 5192 -5232 5252 -5172
rect 5192 -5362 5252 -5302
rect 5650 -5232 5710 -5172
rect 5650 -5362 5710 -5302
rect 6106 -5232 6166 -5172
rect 6106 -5362 6166 -5302
rect 6562 -5232 6622 -5172
rect 6562 -5362 6622 -5302
rect 7020 -5232 7080 -5172
rect 7020 -5362 7080 -5302
rect 7476 -5232 7536 -5172
rect 7476 -5362 7536 -5302
rect 7932 -5232 7992 -5172
rect 7932 -5362 7992 -5302
rect 8406 -5232 8466 -5172
rect 8406 -5362 8466 -5302
rect 8862 -5232 8922 -5172
rect 8862 -5362 8922 -5302
rect 9320 -5232 9380 -5172
rect 9320 -5362 9380 -5302
rect 9776 -5232 9836 -5172
rect 9776 -5362 9836 -5302
rect 10232 -5232 10292 -5172
rect 10232 -5362 10292 -5302
rect 10690 -5232 10750 -5172
rect 10690 -5362 10750 -5302
rect 11146 -5232 11206 -5172
rect 11146 -5362 11206 -5302
rect 11602 -5232 11662 -5172
rect 11602 -5362 11662 -5302
rect 12060 -5232 12120 -5172
rect 12060 -5362 12120 -5302
rect 12516 -5232 12576 -5172
rect 12516 -5362 12576 -5302
rect 12972 -5232 13032 -5172
rect 12972 -5362 13032 -5302
rect 13430 -5232 13490 -5172
rect 13430 -5362 13490 -5302
rect 13886 -5232 13946 -5172
rect 13886 -5362 13946 -5302
rect 14342 -5232 14402 -5172
rect 14342 -5362 14402 -5302
rect 14800 -5232 14860 -5172
rect 14800 -5362 14860 -5302
rect 15256 -5232 15316 -5172
rect 15256 -5362 15316 -5302
rect 170 -5724 230 -5664
rect 170 -5854 230 -5794
rect 626 -5724 686 -5664
rect 626 -5854 686 -5794
rect 1082 -5724 1142 -5664
rect 1082 -5854 1142 -5794
rect 1540 -5724 1600 -5664
rect 1540 -5854 1600 -5794
rect 1996 -5724 2056 -5664
rect 1996 -5854 2056 -5794
rect 2452 -5724 2512 -5664
rect 2452 -5854 2512 -5794
rect 2910 -5724 2970 -5664
rect 2910 -5854 2970 -5794
rect 3366 -5724 3426 -5664
rect 3366 -5854 3426 -5794
rect 3822 -5724 3882 -5664
rect 3822 -5854 3882 -5794
rect 4280 -5724 4340 -5664
rect 4280 -5854 4340 -5794
rect 4736 -5724 4796 -5664
rect 4736 -5854 4796 -5794
rect 5192 -5724 5252 -5664
rect 5192 -5854 5252 -5794
rect 5650 -5724 5710 -5664
rect 5650 -5854 5710 -5794
rect 6106 -5724 6166 -5664
rect 6106 -5854 6166 -5794
rect 6562 -5724 6622 -5664
rect 6562 -5854 6622 -5794
rect 7020 -5724 7080 -5664
rect 7020 -5854 7080 -5794
rect 7476 -5724 7536 -5664
rect 7476 -5854 7536 -5794
rect 7932 -5724 7992 -5664
rect 7932 -5854 7992 -5794
rect 8406 -5724 8466 -5664
rect 8406 -5854 8466 -5794
rect 8862 -5724 8922 -5664
rect 8862 -5854 8922 -5794
rect 9320 -5724 9380 -5664
rect 9320 -5854 9380 -5794
rect 9776 -5724 9836 -5664
rect 9776 -5854 9836 -5794
rect 10232 -5724 10292 -5664
rect 10232 -5854 10292 -5794
rect 10690 -5724 10750 -5664
rect 10690 -5854 10750 -5794
rect 11146 -5724 11206 -5664
rect 11146 -5854 11206 -5794
rect 11602 -5724 11662 -5664
rect 11602 -5854 11662 -5794
rect 12060 -5724 12120 -5664
rect 12060 -5854 12120 -5794
rect 12516 -5724 12576 -5664
rect 12516 -5854 12576 -5794
rect 12972 -5724 13032 -5664
rect 12972 -5854 13032 -5794
rect 13430 -5724 13490 -5664
rect 13430 -5854 13490 -5794
rect 13886 -5724 13946 -5664
rect 13886 -5854 13946 -5794
rect 14342 -5724 14402 -5664
rect 14342 -5854 14402 -5794
rect 14800 -5724 14860 -5664
rect 14800 -5854 14860 -5794
rect 15256 -5724 15316 -5664
rect 15256 -5854 15316 -5794
rect 171 -6221 231 -6161
rect 171 -6351 231 -6291
rect 627 -6221 687 -6161
rect 627 -6351 687 -6291
rect 1083 -6221 1143 -6161
rect 1083 -6351 1143 -6291
rect 1541 -6221 1601 -6161
rect 1541 -6351 1601 -6291
rect 1997 -6221 2057 -6161
rect 1997 -6351 2057 -6291
rect 2453 -6221 2513 -6161
rect 2453 -6351 2513 -6291
rect 2911 -6221 2971 -6161
rect 2911 -6351 2971 -6291
rect 3367 -6221 3427 -6161
rect 3367 -6351 3427 -6291
rect 3823 -6221 3883 -6161
rect 3823 -6351 3883 -6291
rect 4281 -6221 4341 -6161
rect 4281 -6351 4341 -6291
rect 4737 -6221 4797 -6161
rect 4737 -6351 4797 -6291
rect 5193 -6221 5253 -6161
rect 5193 -6351 5253 -6291
rect 5651 -6221 5711 -6161
rect 5651 -6351 5711 -6291
rect 6107 -6221 6167 -6161
rect 6107 -6351 6167 -6291
rect 6563 -6221 6623 -6161
rect 6563 -6351 6623 -6291
rect 7021 -6221 7081 -6161
rect 7021 -6351 7081 -6291
rect 7477 -6221 7537 -6161
rect 7477 -6351 7537 -6291
rect 7933 -6221 7993 -6161
rect 7933 -6351 7993 -6291
rect 8407 -6221 8467 -6161
rect 8407 -6351 8467 -6291
rect 8863 -6221 8923 -6161
rect 8863 -6351 8923 -6291
rect 9321 -6221 9381 -6161
rect 9321 -6351 9381 -6291
rect 9777 -6221 9837 -6161
rect 9777 -6351 9837 -6291
rect 10233 -6221 10293 -6161
rect 10233 -6351 10293 -6291
rect 10691 -6221 10751 -6161
rect 10691 -6351 10751 -6291
rect 11147 -6221 11207 -6161
rect 11147 -6351 11207 -6291
rect 11603 -6221 11663 -6161
rect 11603 -6351 11663 -6291
rect 12061 -6221 12121 -6161
rect 12061 -6351 12121 -6291
rect 12517 -6221 12577 -6161
rect 12517 -6351 12577 -6291
rect 12973 -6221 13033 -6161
rect 12973 -6351 13033 -6291
rect 13431 -6221 13491 -6161
rect 13431 -6351 13491 -6291
rect 13887 -6221 13947 -6161
rect 13887 -6351 13947 -6291
rect 14343 -6221 14403 -6161
rect 14343 -6351 14403 -6291
rect 14801 -6221 14861 -6161
rect 14801 -6351 14861 -6291
rect 15257 -6221 15317 -6161
rect 15257 -6351 15317 -6291
rect 171 -6713 231 -6653
rect 171 -6843 231 -6783
rect 627 -6713 687 -6653
rect 627 -6843 687 -6783
rect 1083 -6713 1143 -6653
rect 1083 -6843 1143 -6783
rect 1541 -6713 1601 -6653
rect 1541 -6843 1601 -6783
rect 1997 -6713 2057 -6653
rect 1997 -6843 2057 -6783
rect 2453 -6713 2513 -6653
rect 2453 -6843 2513 -6783
rect 2911 -6713 2971 -6653
rect 2911 -6843 2971 -6783
rect 3367 -6713 3427 -6653
rect 3367 -6843 3427 -6783
rect 3823 -6713 3883 -6653
rect 3823 -6843 3883 -6783
rect 4281 -6713 4341 -6653
rect 4281 -6843 4341 -6783
rect 4737 -6713 4797 -6653
rect 4737 -6843 4797 -6783
rect 5193 -6713 5253 -6653
rect 5193 -6843 5253 -6783
rect 5651 -6713 5711 -6653
rect 5651 -6843 5711 -6783
rect 6107 -6713 6167 -6653
rect 6107 -6843 6167 -6783
rect 6563 -6713 6623 -6653
rect 6563 -6843 6623 -6783
rect 7021 -6713 7081 -6653
rect 7021 -6843 7081 -6783
rect 7477 -6713 7537 -6653
rect 7477 -6843 7537 -6783
rect 7933 -6713 7993 -6653
rect 7933 -6843 7993 -6783
rect 8407 -6713 8467 -6653
rect 8407 -6843 8467 -6783
rect 8863 -6713 8923 -6653
rect 8863 -6843 8923 -6783
rect 9321 -6713 9381 -6653
rect 9321 -6843 9381 -6783
rect 9777 -6713 9837 -6653
rect 9777 -6843 9837 -6783
rect 10233 -6713 10293 -6653
rect 10233 -6843 10293 -6783
rect 10691 -6713 10751 -6653
rect 10691 -6843 10751 -6783
rect 11147 -6713 11207 -6653
rect 11147 -6843 11207 -6783
rect 11603 -6713 11663 -6653
rect 11603 -6843 11663 -6783
rect 12061 -6713 12121 -6653
rect 12061 -6843 12121 -6783
rect 12517 -6713 12577 -6653
rect 12517 -6843 12577 -6783
rect 12973 -6713 13033 -6653
rect 12973 -6843 13033 -6783
rect 13431 -6713 13491 -6653
rect 13431 -6843 13491 -6783
rect 13887 -6713 13947 -6653
rect 13887 -6843 13947 -6783
rect 14343 -6713 14403 -6653
rect 14343 -6843 14403 -6783
rect 14801 -6713 14861 -6653
rect 14801 -6843 14861 -6783
rect 15257 -6713 15317 -6653
rect 15257 -6843 15317 -6783
rect 171 -7229 231 -7169
rect 171 -7359 231 -7299
rect 627 -7229 687 -7169
rect 627 -7359 687 -7299
rect 1083 -7229 1143 -7169
rect 1083 -7359 1143 -7299
rect 1541 -7229 1601 -7169
rect 1541 -7359 1601 -7299
rect 1997 -7229 2057 -7169
rect 1997 -7359 2057 -7299
rect 2453 -7229 2513 -7169
rect 2453 -7359 2513 -7299
rect 2911 -7229 2971 -7169
rect 2911 -7359 2971 -7299
rect 3367 -7229 3427 -7169
rect 3367 -7359 3427 -7299
rect 3823 -7229 3883 -7169
rect 3823 -7359 3883 -7299
rect 4281 -7229 4341 -7169
rect 4281 -7359 4341 -7299
rect 4737 -7229 4797 -7169
rect 4737 -7359 4797 -7299
rect 5193 -7229 5253 -7169
rect 5193 -7359 5253 -7299
rect 5651 -7229 5711 -7169
rect 5651 -7359 5711 -7299
rect 6107 -7229 6167 -7169
rect 6107 -7359 6167 -7299
rect 6563 -7229 6623 -7169
rect 6563 -7359 6623 -7299
rect 7021 -7229 7081 -7169
rect 7021 -7359 7081 -7299
rect 7477 -7229 7537 -7169
rect 7477 -7359 7537 -7299
rect 7933 -7229 7993 -7169
rect 7933 -7359 7993 -7299
rect 8407 -7229 8467 -7169
rect 8407 -7359 8467 -7299
rect 8863 -7229 8923 -7169
rect 8863 -7359 8923 -7299
rect 9321 -7229 9381 -7169
rect 9321 -7359 9381 -7299
rect 9777 -7229 9837 -7169
rect 9777 -7359 9837 -7299
rect 10233 -7229 10293 -7169
rect 10233 -7359 10293 -7299
rect 10691 -7229 10751 -7169
rect 10691 -7359 10751 -7299
rect 11147 -7229 11207 -7169
rect 11147 -7359 11207 -7299
rect 11603 -7229 11663 -7169
rect 11603 -7359 11663 -7299
rect 12061 -7229 12121 -7169
rect 12061 -7359 12121 -7299
rect 12517 -7229 12577 -7169
rect 12517 -7359 12577 -7299
rect 12973 -7229 13033 -7169
rect 12973 -7359 13033 -7299
rect 13431 -7229 13491 -7169
rect 13431 -7359 13491 -7299
rect 13887 -7229 13947 -7169
rect 13887 -7359 13947 -7299
rect 14343 -7229 14403 -7169
rect 14343 -7359 14403 -7299
rect 14801 -7229 14861 -7169
rect 14801 -7359 14861 -7299
rect 15257 -7229 15317 -7169
rect 15257 -7359 15317 -7299
rect 171 -7731 231 -7671
rect 171 -7861 231 -7801
rect 627 -7731 687 -7671
rect 627 -7861 687 -7801
rect 1083 -7731 1143 -7671
rect 1083 -7861 1143 -7801
rect 1541 -7731 1601 -7671
rect 1541 -7861 1601 -7801
rect 1997 -7731 2057 -7671
rect 1997 -7861 2057 -7801
rect 2453 -7731 2513 -7671
rect 2453 -7861 2513 -7801
rect 2911 -7731 2971 -7671
rect 2911 -7861 2971 -7801
rect 3367 -7731 3427 -7671
rect 3367 -7861 3427 -7801
rect 3823 -7731 3883 -7671
rect 3823 -7861 3883 -7801
rect 4281 -7731 4341 -7671
rect 4281 -7861 4341 -7801
rect 4737 -7731 4797 -7671
rect 4737 -7861 4797 -7801
rect 5193 -7731 5253 -7671
rect 5193 -7861 5253 -7801
rect 5651 -7731 5711 -7671
rect 5651 -7861 5711 -7801
rect 6107 -7731 6167 -7671
rect 6107 -7861 6167 -7801
rect 6563 -7731 6623 -7671
rect 6563 -7861 6623 -7801
rect 7021 -7731 7081 -7671
rect 7021 -7861 7081 -7801
rect 7477 -7731 7537 -7671
rect 7477 -7861 7537 -7801
rect 7933 -7731 7993 -7671
rect 7933 -7861 7993 -7801
rect 8407 -7731 8467 -7671
rect 8407 -7861 8467 -7801
rect 8863 -7731 8923 -7671
rect 8863 -7861 8923 -7801
rect 9321 -7731 9381 -7671
rect 9321 -7861 9381 -7801
rect 9777 -7731 9837 -7671
rect 9777 -7861 9837 -7801
rect 10233 -7731 10293 -7671
rect 10233 -7861 10293 -7801
rect 10691 -7731 10751 -7671
rect 10691 -7861 10751 -7801
rect 11147 -7731 11207 -7671
rect 11147 -7861 11207 -7801
rect 11603 -7731 11663 -7671
rect 11603 -7861 11663 -7801
rect 12061 -7731 12121 -7671
rect 12061 -7861 12121 -7801
rect 12517 -7731 12577 -7671
rect 12517 -7861 12577 -7801
rect 12973 -7731 13033 -7671
rect 12973 -7861 13033 -7801
rect 13431 -7731 13491 -7671
rect 13431 -7861 13491 -7801
rect 13887 -7731 13947 -7671
rect 13887 -7861 13947 -7801
rect 14343 -7731 14403 -7671
rect 14343 -7861 14403 -7801
rect 14801 -7731 14861 -7671
rect 14801 -7861 14861 -7801
rect 15257 -7731 15317 -7671
rect 15257 -7861 15317 -7801
rect 171 -8223 231 -8163
rect 171 -8353 231 -8293
rect 627 -8223 687 -8163
rect 627 -8353 687 -8293
rect 1083 -8223 1143 -8163
rect 1083 -8353 1143 -8293
rect 1541 -8223 1601 -8163
rect 1541 -8353 1601 -8293
rect 1997 -8223 2057 -8163
rect 1997 -8353 2057 -8293
rect 2453 -8223 2513 -8163
rect 2453 -8353 2513 -8293
rect 2911 -8223 2971 -8163
rect 2911 -8353 2971 -8293
rect 3367 -8223 3427 -8163
rect 3367 -8353 3427 -8293
rect 3823 -8223 3883 -8163
rect 3823 -8353 3883 -8293
rect 4281 -8223 4341 -8163
rect 4281 -8353 4341 -8293
rect 4737 -8223 4797 -8163
rect 4737 -8353 4797 -8293
rect 5193 -8223 5253 -8163
rect 5193 -8353 5253 -8293
rect 5651 -8223 5711 -8163
rect 5651 -8353 5711 -8293
rect 6107 -8223 6167 -8163
rect 6107 -8353 6167 -8293
rect 6563 -8223 6623 -8163
rect 6563 -8353 6623 -8293
rect 7021 -8223 7081 -8163
rect 7021 -8353 7081 -8293
rect 7477 -8223 7537 -8163
rect 7477 -8353 7537 -8293
rect 7933 -8223 7993 -8163
rect 7933 -8353 7993 -8293
rect 8407 -8223 8467 -8163
rect 8407 -8353 8467 -8293
rect 8863 -8223 8923 -8163
rect 8863 -8353 8923 -8293
rect 9321 -8223 9381 -8163
rect 9321 -8353 9381 -8293
rect 9777 -8223 9837 -8163
rect 9777 -8353 9837 -8293
rect 10233 -8223 10293 -8163
rect 10233 -8353 10293 -8293
rect 10691 -8223 10751 -8163
rect 10691 -8353 10751 -8293
rect 11147 -8223 11207 -8163
rect 11147 -8353 11207 -8293
rect 11603 -8223 11663 -8163
rect 11603 -8353 11663 -8293
rect 12061 -8223 12121 -8163
rect 12061 -8353 12121 -8293
rect 12517 -8223 12577 -8163
rect 12517 -8353 12577 -8293
rect 12973 -8223 13033 -8163
rect 12973 -8353 13033 -8293
rect 13431 -8223 13491 -8163
rect 13431 -8353 13491 -8293
rect 13887 -8223 13947 -8163
rect 13887 -8353 13947 -8293
rect 14343 -8223 14403 -8163
rect 14343 -8353 14403 -8293
rect 14801 -8223 14861 -8163
rect 14801 -8353 14861 -8293
rect 15257 -8223 15317 -8163
rect 15257 -8353 15317 -8293
rect 171 -8717 231 -8657
rect 171 -8847 231 -8787
rect 627 -8717 687 -8657
rect 627 -8847 687 -8787
rect 1083 -8717 1143 -8657
rect 1083 -8847 1143 -8787
rect 1541 -8717 1601 -8657
rect 1541 -8847 1601 -8787
rect 1997 -8717 2057 -8657
rect 1997 -8847 2057 -8787
rect 2453 -8717 2513 -8657
rect 2453 -8847 2513 -8787
rect 2911 -8717 2971 -8657
rect 2911 -8847 2971 -8787
rect 3367 -8717 3427 -8657
rect 3367 -8847 3427 -8787
rect 3823 -8717 3883 -8657
rect 3823 -8847 3883 -8787
rect 4281 -8717 4341 -8657
rect 4281 -8847 4341 -8787
rect 4737 -8717 4797 -8657
rect 4737 -8847 4797 -8787
rect 5193 -8717 5253 -8657
rect 5193 -8847 5253 -8787
rect 5651 -8717 5711 -8657
rect 5651 -8847 5711 -8787
rect 6107 -8717 6167 -8657
rect 6107 -8847 6167 -8787
rect 6563 -8717 6623 -8657
rect 6563 -8847 6623 -8787
rect 7021 -8717 7081 -8657
rect 7021 -8847 7081 -8787
rect 7477 -8717 7537 -8657
rect 7477 -8847 7537 -8787
rect 7933 -8717 7993 -8657
rect 7933 -8847 7993 -8787
rect 8407 -8717 8467 -8657
rect 8407 -8847 8467 -8787
rect 8863 -8717 8923 -8657
rect 8863 -8847 8923 -8787
rect 9321 -8717 9381 -8657
rect 9321 -8847 9381 -8787
rect 9777 -8717 9837 -8657
rect 9777 -8847 9837 -8787
rect 10233 -8717 10293 -8657
rect 10233 -8847 10293 -8787
rect 10691 -8717 10751 -8657
rect 10691 -8847 10751 -8787
rect 11147 -8717 11207 -8657
rect 11147 -8847 11207 -8787
rect 11603 -8717 11663 -8657
rect 11603 -8847 11663 -8787
rect 12061 -8717 12121 -8657
rect 12061 -8847 12121 -8787
rect 12517 -8717 12577 -8657
rect 12517 -8847 12577 -8787
rect 12973 -8717 13033 -8657
rect 12973 -8847 13033 -8787
rect 13431 -8717 13491 -8657
rect 13431 -8847 13491 -8787
rect 13887 -8717 13947 -8657
rect 13887 -8847 13947 -8787
rect 14343 -8717 14403 -8657
rect 14343 -8847 14403 -8787
rect 14801 -8717 14861 -8657
rect 14801 -8847 14861 -8787
rect 15257 -8717 15317 -8657
rect 15257 -8847 15317 -8787
rect 171 -9219 231 -9159
rect 171 -9349 231 -9289
rect 627 -9219 687 -9159
rect 627 -9349 687 -9289
rect 1083 -9219 1143 -9159
rect 1083 -9349 1143 -9289
rect 1541 -9219 1601 -9159
rect 1541 -9349 1601 -9289
rect 1997 -9219 2057 -9159
rect 1997 -9349 2057 -9289
rect 2453 -9219 2513 -9159
rect 2453 -9349 2513 -9289
rect 2911 -9219 2971 -9159
rect 2911 -9349 2971 -9289
rect 3367 -9219 3427 -9159
rect 3367 -9349 3427 -9289
rect 3823 -9219 3883 -9159
rect 3823 -9349 3883 -9289
rect 4281 -9219 4341 -9159
rect 4281 -9349 4341 -9289
rect 4737 -9219 4797 -9159
rect 4737 -9349 4797 -9289
rect 5193 -9219 5253 -9159
rect 5193 -9349 5253 -9289
rect 5651 -9219 5711 -9159
rect 5651 -9349 5711 -9289
rect 6107 -9219 6167 -9159
rect 6107 -9349 6167 -9289
rect 6563 -9219 6623 -9159
rect 6563 -9349 6623 -9289
rect 7021 -9219 7081 -9159
rect 7021 -9349 7081 -9289
rect 7477 -9219 7537 -9159
rect 7477 -9349 7537 -9289
rect 7933 -9219 7993 -9159
rect 7933 -9349 7993 -9289
rect 8407 -9219 8467 -9159
rect 8407 -9349 8467 -9289
rect 8863 -9219 8923 -9159
rect 8863 -9349 8923 -9289
rect 9321 -9219 9381 -9159
rect 9321 -9349 9381 -9289
rect 9777 -9219 9837 -9159
rect 9777 -9349 9837 -9289
rect 10233 -9219 10293 -9159
rect 10233 -9349 10293 -9289
rect 10691 -9219 10751 -9159
rect 10691 -9349 10751 -9289
rect 11147 -9219 11207 -9159
rect 11147 -9349 11207 -9289
rect 11603 -9219 11663 -9159
rect 11603 -9349 11663 -9289
rect 12061 -9219 12121 -9159
rect 12061 -9349 12121 -9289
rect 12517 -9219 12577 -9159
rect 12517 -9349 12577 -9289
rect 12973 -9219 13033 -9159
rect 12973 -9349 13033 -9289
rect 13431 -9219 13491 -9159
rect 13431 -9349 13491 -9289
rect 13887 -9219 13947 -9159
rect 13887 -9349 13947 -9289
rect 14343 -9219 14403 -9159
rect 14343 -9349 14403 -9289
rect 14801 -9219 14861 -9159
rect 14801 -9349 14861 -9289
rect 15257 -9219 15317 -9159
rect 15257 -9349 15317 -9289
rect 171 -9711 231 -9651
rect 171 -9841 231 -9781
rect 627 -9711 687 -9651
rect 627 -9841 687 -9781
rect 1083 -9711 1143 -9651
rect 1083 -9841 1143 -9781
rect 1541 -9711 1601 -9651
rect 1541 -9841 1601 -9781
rect 1997 -9711 2057 -9651
rect 1997 -9841 2057 -9781
rect 2453 -9711 2513 -9651
rect 2453 -9841 2513 -9781
rect 2911 -9711 2971 -9651
rect 2911 -9841 2971 -9781
rect 3367 -9711 3427 -9651
rect 3367 -9841 3427 -9781
rect 3823 -9711 3883 -9651
rect 3823 -9841 3883 -9781
rect 4281 -9711 4341 -9651
rect 4281 -9841 4341 -9781
rect 4737 -9711 4797 -9651
rect 4737 -9841 4797 -9781
rect 5193 -9711 5253 -9651
rect 5193 -9841 5253 -9781
rect 5651 -9711 5711 -9651
rect 5651 -9841 5711 -9781
rect 6107 -9711 6167 -9651
rect 6107 -9841 6167 -9781
rect 6563 -9711 6623 -9651
rect 6563 -9841 6623 -9781
rect 7021 -9711 7081 -9651
rect 7021 -9841 7081 -9781
rect 7477 -9711 7537 -9651
rect 7477 -9841 7537 -9781
rect 7933 -9711 7993 -9651
rect 7933 -9841 7993 -9781
rect 8407 -9711 8467 -9651
rect 8407 -9841 8467 -9781
rect 8863 -9711 8923 -9651
rect 8863 -9841 8923 -9781
rect 9321 -9711 9381 -9651
rect 9321 -9841 9381 -9781
rect 9777 -9711 9837 -9651
rect 9777 -9841 9837 -9781
rect 10233 -9711 10293 -9651
rect 10233 -9841 10293 -9781
rect 10691 -9711 10751 -9651
rect 10691 -9841 10751 -9781
rect 11147 -9711 11207 -9651
rect 11147 -9841 11207 -9781
rect 11603 -9711 11663 -9651
rect 11603 -9841 11663 -9781
rect 12061 -9711 12121 -9651
rect 12061 -9841 12121 -9781
rect 12517 -9711 12577 -9651
rect 12517 -9841 12577 -9781
rect 12973 -9711 13033 -9651
rect 12973 -9841 13033 -9781
rect 13431 -9711 13491 -9651
rect 13431 -9841 13491 -9781
rect 13887 -9711 13947 -9651
rect 13887 -9841 13947 -9781
rect 14343 -9711 14403 -9651
rect 14343 -9841 14403 -9781
rect 14801 -9711 14861 -9651
rect 14801 -9841 14861 -9781
rect 15257 -9711 15317 -9651
rect 15257 -9841 15317 -9781
rect 171 -10227 231 -10167
rect 171 -10357 231 -10297
rect 627 -10227 687 -10167
rect 627 -10357 687 -10297
rect 1083 -10227 1143 -10167
rect 1083 -10357 1143 -10297
rect 1541 -10227 1601 -10167
rect 1541 -10357 1601 -10297
rect 1997 -10227 2057 -10167
rect 1997 -10357 2057 -10297
rect 2453 -10227 2513 -10167
rect 2453 -10357 2513 -10297
rect 2911 -10227 2971 -10167
rect 2911 -10357 2971 -10297
rect 3367 -10227 3427 -10167
rect 3367 -10357 3427 -10297
rect 3823 -10227 3883 -10167
rect 3823 -10357 3883 -10297
rect 4281 -10227 4341 -10167
rect 4281 -10357 4341 -10297
rect 4737 -10227 4797 -10167
rect 4737 -10357 4797 -10297
rect 5193 -10227 5253 -10167
rect 5193 -10357 5253 -10297
rect 5651 -10227 5711 -10167
rect 5651 -10357 5711 -10297
rect 6107 -10227 6167 -10167
rect 6107 -10357 6167 -10297
rect 6563 -10227 6623 -10167
rect 6563 -10357 6623 -10297
rect 7021 -10227 7081 -10167
rect 7021 -10357 7081 -10297
rect 7477 -10227 7537 -10167
rect 7477 -10357 7537 -10297
rect 7933 -10227 7993 -10167
rect 7933 -10357 7993 -10297
rect 8407 -10227 8467 -10167
rect 8407 -10357 8467 -10297
rect 8863 -10227 8923 -10167
rect 8863 -10357 8923 -10297
rect 9321 -10227 9381 -10167
rect 9321 -10357 9381 -10297
rect 9777 -10227 9837 -10167
rect 9777 -10357 9837 -10297
rect 10233 -10227 10293 -10167
rect 10233 -10357 10293 -10297
rect 10691 -10227 10751 -10167
rect 10691 -10357 10751 -10297
rect 11147 -10227 11207 -10167
rect 11147 -10357 11207 -10297
rect 11603 -10227 11663 -10167
rect 11603 -10357 11663 -10297
rect 12061 -10227 12121 -10167
rect 12061 -10357 12121 -10297
rect 12517 -10227 12577 -10167
rect 12517 -10357 12577 -10297
rect 12973 -10227 13033 -10167
rect 12973 -10357 13033 -10297
rect 13431 -10227 13491 -10167
rect 13431 -10357 13491 -10297
rect 13887 -10227 13947 -10167
rect 13887 -10357 13947 -10297
rect 14343 -10227 14403 -10167
rect 14343 -10357 14403 -10297
rect 14801 -10227 14861 -10167
rect 14801 -10357 14861 -10297
rect 15257 -10227 15317 -10167
rect 15257 -10357 15317 -10297
rect 171 -10729 231 -10669
rect 171 -10859 231 -10799
rect 627 -10729 687 -10669
rect 627 -10859 687 -10799
rect 1083 -10729 1143 -10669
rect 1083 -10859 1143 -10799
rect 1541 -10729 1601 -10669
rect 1541 -10859 1601 -10799
rect 1997 -10729 2057 -10669
rect 1997 -10859 2057 -10799
rect 2453 -10729 2513 -10669
rect 2453 -10859 2513 -10799
rect 2911 -10729 2971 -10669
rect 2911 -10859 2971 -10799
rect 3367 -10729 3427 -10669
rect 3367 -10859 3427 -10799
rect 3823 -10729 3883 -10669
rect 3823 -10859 3883 -10799
rect 4281 -10729 4341 -10669
rect 4281 -10859 4341 -10799
rect 4737 -10729 4797 -10669
rect 4737 -10859 4797 -10799
rect 5193 -10729 5253 -10669
rect 5193 -10859 5253 -10799
rect 5651 -10729 5711 -10669
rect 5651 -10859 5711 -10799
rect 6107 -10729 6167 -10669
rect 6107 -10859 6167 -10799
rect 6563 -10729 6623 -10669
rect 6563 -10859 6623 -10799
rect 7021 -10729 7081 -10669
rect 7021 -10859 7081 -10799
rect 7477 -10729 7537 -10669
rect 7477 -10859 7537 -10799
rect 7933 -10729 7993 -10669
rect 7933 -10859 7993 -10799
rect 8407 -10729 8467 -10669
rect 8407 -10859 8467 -10799
rect 8863 -10729 8923 -10669
rect 8863 -10859 8923 -10799
rect 9321 -10729 9381 -10669
rect 9321 -10859 9381 -10799
rect 9777 -10729 9837 -10669
rect 9777 -10859 9837 -10799
rect 10233 -10729 10293 -10669
rect 10233 -10859 10293 -10799
rect 10691 -10729 10751 -10669
rect 10691 -10859 10751 -10799
rect 11147 -10729 11207 -10669
rect 11147 -10859 11207 -10799
rect 11603 -10729 11663 -10669
rect 11603 -10859 11663 -10799
rect 12061 -10729 12121 -10669
rect 12061 -10859 12121 -10799
rect 12517 -10729 12577 -10669
rect 12517 -10859 12577 -10799
rect 12973 -10729 13033 -10669
rect 12973 -10859 13033 -10799
rect 13431 -10729 13491 -10669
rect 13431 -10859 13491 -10799
rect 13887 -10729 13947 -10669
rect 13887 -10859 13947 -10799
rect 14343 -10729 14403 -10669
rect 14343 -10859 14403 -10799
rect 14801 -10729 14861 -10669
rect 14801 -10859 14861 -10799
rect 15257 -10729 15317 -10669
rect 15257 -10859 15317 -10799
rect 171 -11221 231 -11161
rect 171 -11351 231 -11291
rect 627 -11221 687 -11161
rect 627 -11351 687 -11291
rect 1083 -11221 1143 -11161
rect 1083 -11351 1143 -11291
rect 1541 -11221 1601 -11161
rect 1541 -11351 1601 -11291
rect 1997 -11221 2057 -11161
rect 1997 -11351 2057 -11291
rect 2453 -11221 2513 -11161
rect 2453 -11351 2513 -11291
rect 2911 -11221 2971 -11161
rect 2911 -11351 2971 -11291
rect 3367 -11221 3427 -11161
rect 3367 -11351 3427 -11291
rect 3823 -11221 3883 -11161
rect 3823 -11351 3883 -11291
rect 4281 -11221 4341 -11161
rect 4281 -11351 4341 -11291
rect 4737 -11221 4797 -11161
rect 4737 -11351 4797 -11291
rect 5193 -11221 5253 -11161
rect 5193 -11351 5253 -11291
rect 5651 -11221 5711 -11161
rect 5651 -11351 5711 -11291
rect 6107 -11221 6167 -11161
rect 6107 -11351 6167 -11291
rect 6563 -11221 6623 -11161
rect 6563 -11351 6623 -11291
rect 7021 -11221 7081 -11161
rect 7021 -11351 7081 -11291
rect 7477 -11221 7537 -11161
rect 7477 -11351 7537 -11291
rect 7933 -11221 7993 -11161
rect 7933 -11351 7993 -11291
rect 8407 -11221 8467 -11161
rect 8407 -11351 8467 -11291
rect 8863 -11221 8923 -11161
rect 8863 -11351 8923 -11291
rect 9321 -11221 9381 -11161
rect 9321 -11351 9381 -11291
rect 9777 -11221 9837 -11161
rect 9777 -11351 9837 -11291
rect 10233 -11221 10293 -11161
rect 10233 -11351 10293 -11291
rect 10691 -11221 10751 -11161
rect 10691 -11351 10751 -11291
rect 11147 -11221 11207 -11161
rect 11147 -11351 11207 -11291
rect 11603 -11221 11663 -11161
rect 11603 -11351 11663 -11291
rect 12061 -11221 12121 -11161
rect 12061 -11351 12121 -11291
rect 12517 -11221 12577 -11161
rect 12517 -11351 12577 -11291
rect 12973 -11221 13033 -11161
rect 12973 -11351 13033 -11291
rect 13431 -11221 13491 -11161
rect 13431 -11351 13491 -11291
rect 13887 -11221 13947 -11161
rect 13887 -11351 13947 -11291
rect 14343 -11221 14403 -11161
rect 14343 -11351 14403 -11291
rect 14801 -11221 14861 -11161
rect 14801 -11351 14861 -11291
rect 15257 -11221 15317 -11161
rect 15257 -11351 15317 -11291
rect 170 -11714 230 -11654
rect 170 -11844 230 -11784
rect 626 -11714 686 -11654
rect 626 -11844 686 -11784
rect 1082 -11714 1142 -11654
rect 1082 -11844 1142 -11784
rect 1540 -11714 1600 -11654
rect 1540 -11844 1600 -11784
rect 1996 -11714 2056 -11654
rect 1996 -11844 2056 -11784
rect 2452 -11714 2512 -11654
rect 2452 -11844 2512 -11784
rect 2910 -11714 2970 -11654
rect 2910 -11844 2970 -11784
rect 3366 -11714 3426 -11654
rect 3366 -11844 3426 -11784
rect 3822 -11714 3882 -11654
rect 3822 -11844 3882 -11784
rect 4280 -11714 4340 -11654
rect 4280 -11844 4340 -11784
rect 4736 -11714 4796 -11654
rect 4736 -11844 4796 -11784
rect 5192 -11714 5252 -11654
rect 5192 -11844 5252 -11784
rect 5650 -11714 5710 -11654
rect 5650 -11844 5710 -11784
rect 6106 -11714 6166 -11654
rect 6106 -11844 6166 -11784
rect 6562 -11714 6622 -11654
rect 6562 -11844 6622 -11784
rect 7020 -11714 7080 -11654
rect 7020 -11844 7080 -11784
rect 7476 -11714 7536 -11654
rect 7476 -11844 7536 -11784
rect 7932 -11714 7992 -11654
rect 7932 -11844 7992 -11784
rect 8406 -11714 8466 -11654
rect 8406 -11844 8466 -11784
rect 8862 -11714 8922 -11654
rect 8862 -11844 8922 -11784
rect 9320 -11714 9380 -11654
rect 9320 -11844 9380 -11784
rect 9776 -11714 9836 -11654
rect 9776 -11844 9836 -11784
rect 10232 -11714 10292 -11654
rect 10232 -11844 10292 -11784
rect 10690 -11714 10750 -11654
rect 10690 -11844 10750 -11784
rect 11146 -11714 11206 -11654
rect 11146 -11844 11206 -11784
rect 11602 -11714 11662 -11654
rect 11602 -11844 11662 -11784
rect 12060 -11714 12120 -11654
rect 12060 -11844 12120 -11784
rect 12516 -11714 12576 -11654
rect 12516 -11844 12576 -11784
rect 12972 -11714 13032 -11654
rect 12972 -11844 13032 -11784
rect 13430 -11714 13490 -11654
rect 13430 -11844 13490 -11784
rect 13886 -11714 13946 -11654
rect 13886 -11844 13946 -11784
rect 14342 -11714 14402 -11654
rect 14342 -11844 14402 -11784
rect 14800 -11714 14860 -11654
rect 14800 -11844 14860 -11784
rect 15256 -11714 15316 -11654
rect 15256 -11844 15316 -11784
rect 170 -12206 230 -12146
rect 170 -12336 230 -12276
rect 626 -12206 686 -12146
rect 626 -12336 686 -12276
rect 1082 -12206 1142 -12146
rect 1082 -12336 1142 -12276
rect 1540 -12206 1600 -12146
rect 1540 -12336 1600 -12276
rect 1996 -12206 2056 -12146
rect 1996 -12336 2056 -12276
rect 2452 -12206 2512 -12146
rect 2452 -12336 2512 -12276
rect 2910 -12206 2970 -12146
rect 2910 -12336 2970 -12276
rect 3366 -12206 3426 -12146
rect 3366 -12336 3426 -12276
rect 3822 -12206 3882 -12146
rect 3822 -12336 3882 -12276
rect 4280 -12206 4340 -12146
rect 4280 -12336 4340 -12276
rect 4736 -12206 4796 -12146
rect 4736 -12336 4796 -12276
rect 5192 -12206 5252 -12146
rect 5192 -12336 5252 -12276
rect 5650 -12206 5710 -12146
rect 5650 -12336 5710 -12276
rect 6106 -12206 6166 -12146
rect 6106 -12336 6166 -12276
rect 6562 -12206 6622 -12146
rect 6562 -12336 6622 -12276
rect 7020 -12206 7080 -12146
rect 7020 -12336 7080 -12276
rect 7476 -12206 7536 -12146
rect 7476 -12336 7536 -12276
rect 7932 -12206 7992 -12146
rect 7932 -12336 7992 -12276
rect 8406 -12206 8466 -12146
rect 8406 -12336 8466 -12276
rect 8862 -12206 8922 -12146
rect 8862 -12336 8922 -12276
rect 9320 -12206 9380 -12146
rect 9320 -12336 9380 -12276
rect 9776 -12206 9836 -12146
rect 9776 -12336 9836 -12276
rect 10232 -12206 10292 -12146
rect 10232 -12336 10292 -12276
rect 10690 -12206 10750 -12146
rect 10690 -12336 10750 -12276
rect 11146 -12206 11206 -12146
rect 11146 -12336 11206 -12276
rect 11602 -12206 11662 -12146
rect 11602 -12336 11662 -12276
rect 12060 -12206 12120 -12146
rect 12060 -12336 12120 -12276
rect 12516 -12206 12576 -12146
rect 12516 -12336 12576 -12276
rect 12972 -12206 13032 -12146
rect 12972 -12336 13032 -12276
rect 13430 -12206 13490 -12146
rect 13430 -12336 13490 -12276
rect 13886 -12206 13946 -12146
rect 13886 -12336 13946 -12276
rect 14342 -12206 14402 -12146
rect 14342 -12336 14402 -12276
rect 14800 -12206 14860 -12146
rect 14800 -12336 14860 -12276
rect 15256 -12206 15316 -12146
rect 15256 -12336 15316 -12276
rect 170 -12722 230 -12662
rect 170 -12852 230 -12792
rect 626 -12722 686 -12662
rect 626 -12852 686 -12792
rect 1082 -12722 1142 -12662
rect 1082 -12852 1142 -12792
rect 1540 -12722 1600 -12662
rect 1540 -12852 1600 -12792
rect 1996 -12722 2056 -12662
rect 1996 -12852 2056 -12792
rect 2452 -12722 2512 -12662
rect 2452 -12852 2512 -12792
rect 2910 -12722 2970 -12662
rect 2910 -12852 2970 -12792
rect 3366 -12722 3426 -12662
rect 3366 -12852 3426 -12792
rect 3822 -12722 3882 -12662
rect 3822 -12852 3882 -12792
rect 4280 -12722 4340 -12662
rect 4280 -12852 4340 -12792
rect 4736 -12722 4796 -12662
rect 4736 -12852 4796 -12792
rect 5192 -12722 5252 -12662
rect 5192 -12852 5252 -12792
rect 5650 -12722 5710 -12662
rect 5650 -12852 5710 -12792
rect 6106 -12722 6166 -12662
rect 6106 -12852 6166 -12792
rect 6562 -12722 6622 -12662
rect 6562 -12852 6622 -12792
rect 7020 -12722 7080 -12662
rect 7020 -12852 7080 -12792
rect 7476 -12722 7536 -12662
rect 7476 -12852 7536 -12792
rect 7932 -12722 7992 -12662
rect 7932 -12852 7992 -12792
rect 8406 -12722 8466 -12662
rect 8406 -12852 8466 -12792
rect 8862 -12722 8922 -12662
rect 8862 -12852 8922 -12792
rect 9320 -12722 9380 -12662
rect 9320 -12852 9380 -12792
rect 9776 -12722 9836 -12662
rect 9776 -12852 9836 -12792
rect 10232 -12722 10292 -12662
rect 10232 -12852 10292 -12792
rect 10690 -12722 10750 -12662
rect 10690 -12852 10750 -12792
rect 11146 -12722 11206 -12662
rect 11146 -12852 11206 -12792
rect 11602 -12722 11662 -12662
rect 11602 -12852 11662 -12792
rect 12060 -12722 12120 -12662
rect 12060 -12852 12120 -12792
rect 12516 -12722 12576 -12662
rect 12516 -12852 12576 -12792
rect 12972 -12722 13032 -12662
rect 12972 -12852 13032 -12792
rect 13430 -12722 13490 -12662
rect 13430 -12852 13490 -12792
rect 13886 -12722 13946 -12662
rect 13886 -12852 13946 -12792
rect 14342 -12722 14402 -12662
rect 14342 -12852 14402 -12792
rect 14800 -12722 14860 -12662
rect 14800 -12852 14860 -12792
rect 15256 -12722 15316 -12662
rect 15256 -12852 15316 -12792
rect 170 -13224 230 -13164
rect 170 -13354 230 -13294
rect 626 -13224 686 -13164
rect 626 -13354 686 -13294
rect 1082 -13224 1142 -13164
rect 1082 -13354 1142 -13294
rect 1540 -13224 1600 -13164
rect 1540 -13354 1600 -13294
rect 1996 -13224 2056 -13164
rect 1996 -13354 2056 -13294
rect 2452 -13224 2512 -13164
rect 2452 -13354 2512 -13294
rect 2910 -13224 2970 -13164
rect 2910 -13354 2970 -13294
rect 3366 -13224 3426 -13164
rect 3366 -13354 3426 -13294
rect 3822 -13224 3882 -13164
rect 3822 -13354 3882 -13294
rect 4280 -13224 4340 -13164
rect 4280 -13354 4340 -13294
rect 4736 -13224 4796 -13164
rect 4736 -13354 4796 -13294
rect 5192 -13224 5252 -13164
rect 5192 -13354 5252 -13294
rect 5650 -13224 5710 -13164
rect 5650 -13354 5710 -13294
rect 6106 -13224 6166 -13164
rect 6106 -13354 6166 -13294
rect 6562 -13224 6622 -13164
rect 6562 -13354 6622 -13294
rect 7020 -13224 7080 -13164
rect 7020 -13354 7080 -13294
rect 7476 -13224 7536 -13164
rect 7476 -13354 7536 -13294
rect 7932 -13224 7992 -13164
rect 7932 -13354 7992 -13294
rect 8406 -13224 8466 -13164
rect 8406 -13354 8466 -13294
rect 8862 -13224 8922 -13164
rect 8862 -13354 8922 -13294
rect 9320 -13224 9380 -13164
rect 9320 -13354 9380 -13294
rect 9776 -13224 9836 -13164
rect 9776 -13354 9836 -13294
rect 10232 -13224 10292 -13164
rect 10232 -13354 10292 -13294
rect 10690 -13224 10750 -13164
rect 10690 -13354 10750 -13294
rect 11146 -13224 11206 -13164
rect 11146 -13354 11206 -13294
rect 11602 -13224 11662 -13164
rect 11602 -13354 11662 -13294
rect 12060 -13224 12120 -13164
rect 12060 -13354 12120 -13294
rect 12516 -13224 12576 -13164
rect 12516 -13354 12576 -13294
rect 12972 -13224 13032 -13164
rect 12972 -13354 13032 -13294
rect 13430 -13224 13490 -13164
rect 13430 -13354 13490 -13294
rect 13886 -13224 13946 -13164
rect 13886 -13354 13946 -13294
rect 14342 -13224 14402 -13164
rect 14342 -13354 14402 -13294
rect 14800 -13224 14860 -13164
rect 14800 -13354 14860 -13294
rect 15256 -13224 15316 -13164
rect 15256 -13354 15316 -13294
rect 170 -13716 230 -13656
rect 170 -13846 230 -13786
rect 626 -13716 686 -13656
rect 626 -13846 686 -13786
rect 1082 -13716 1142 -13656
rect 1082 -13846 1142 -13786
rect 1540 -13716 1600 -13656
rect 1540 -13846 1600 -13786
rect 1996 -13716 2056 -13656
rect 1996 -13846 2056 -13786
rect 2452 -13716 2512 -13656
rect 2452 -13846 2512 -13786
rect 2910 -13716 2970 -13656
rect 2910 -13846 2970 -13786
rect 3366 -13716 3426 -13656
rect 3366 -13846 3426 -13786
rect 3822 -13716 3882 -13656
rect 3822 -13846 3882 -13786
rect 4280 -13716 4340 -13656
rect 4280 -13846 4340 -13786
rect 4736 -13716 4796 -13656
rect 4736 -13846 4796 -13786
rect 5192 -13716 5252 -13656
rect 5192 -13846 5252 -13786
rect 5650 -13716 5710 -13656
rect 5650 -13846 5710 -13786
rect 6106 -13716 6166 -13656
rect 6106 -13846 6166 -13786
rect 6562 -13716 6622 -13656
rect 6562 -13846 6622 -13786
rect 7020 -13716 7080 -13656
rect 7020 -13846 7080 -13786
rect 7476 -13716 7536 -13656
rect 7476 -13846 7536 -13786
rect 7932 -13716 7992 -13656
rect 7932 -13846 7992 -13786
rect 8406 -13716 8466 -13656
rect 8406 -13846 8466 -13786
rect 8862 -13716 8922 -13656
rect 8862 -13846 8922 -13786
rect 9320 -13716 9380 -13656
rect 9320 -13846 9380 -13786
rect 9776 -13716 9836 -13656
rect 9776 -13846 9836 -13786
rect 10232 -13716 10292 -13656
rect 10232 -13846 10292 -13786
rect 10690 -13716 10750 -13656
rect 10690 -13846 10750 -13786
rect 11146 -13716 11206 -13656
rect 11146 -13846 11206 -13786
rect 11602 -13716 11662 -13656
rect 11602 -13846 11662 -13786
rect 12060 -13716 12120 -13656
rect 12060 -13846 12120 -13786
rect 12516 -13716 12576 -13656
rect 12516 -13846 12576 -13786
rect 12972 -13716 13032 -13656
rect 12972 -13846 13032 -13786
rect 13430 -13716 13490 -13656
rect 13430 -13846 13490 -13786
rect 13886 -13716 13946 -13656
rect 13886 -13846 13946 -13786
rect 14342 -13716 14402 -13656
rect 14342 -13846 14402 -13786
rect 14800 -13716 14860 -13656
rect 14800 -13846 14860 -13786
rect 15256 -13716 15316 -13656
rect 15256 -13846 15316 -13786
rect 170 -14210 230 -14150
rect 170 -14340 230 -14280
rect 626 -14210 686 -14150
rect 626 -14340 686 -14280
rect 1082 -14210 1142 -14150
rect 1082 -14340 1142 -14280
rect 1540 -14210 1600 -14150
rect 1540 -14340 1600 -14280
rect 1996 -14210 2056 -14150
rect 1996 -14340 2056 -14280
rect 2452 -14210 2512 -14150
rect 2452 -14340 2512 -14280
rect 2910 -14210 2970 -14150
rect 2910 -14340 2970 -14280
rect 3366 -14210 3426 -14150
rect 3366 -14340 3426 -14280
rect 3822 -14210 3882 -14150
rect 3822 -14340 3882 -14280
rect 4280 -14210 4340 -14150
rect 4280 -14340 4340 -14280
rect 4736 -14210 4796 -14150
rect 4736 -14340 4796 -14280
rect 5192 -14210 5252 -14150
rect 5192 -14340 5252 -14280
rect 5650 -14210 5710 -14150
rect 5650 -14340 5710 -14280
rect 6106 -14210 6166 -14150
rect 6106 -14340 6166 -14280
rect 6562 -14210 6622 -14150
rect 6562 -14340 6622 -14280
rect 7020 -14210 7080 -14150
rect 7020 -14340 7080 -14280
rect 7476 -14210 7536 -14150
rect 7476 -14340 7536 -14280
rect 7932 -14210 7992 -14150
rect 7932 -14340 7992 -14280
rect 8406 -14210 8466 -14150
rect 8406 -14340 8466 -14280
rect 8862 -14210 8922 -14150
rect 8862 -14340 8922 -14280
rect 9320 -14210 9380 -14150
rect 9320 -14340 9380 -14280
rect 9776 -14210 9836 -14150
rect 9776 -14340 9836 -14280
rect 10232 -14210 10292 -14150
rect 10232 -14340 10292 -14280
rect 10690 -14210 10750 -14150
rect 10690 -14340 10750 -14280
rect 11146 -14210 11206 -14150
rect 11146 -14340 11206 -14280
rect 11602 -14210 11662 -14150
rect 11602 -14340 11662 -14280
rect 12060 -14210 12120 -14150
rect 12060 -14340 12120 -14280
rect 12516 -14210 12576 -14150
rect 12516 -14340 12576 -14280
rect 12972 -14210 13032 -14150
rect 12972 -14340 13032 -14280
rect 13430 -14210 13490 -14150
rect 13430 -14340 13490 -14280
rect 13886 -14210 13946 -14150
rect 13886 -14340 13946 -14280
rect 14342 -14210 14402 -14150
rect 14342 -14340 14402 -14280
rect 14800 -14210 14860 -14150
rect 14800 -14340 14860 -14280
rect 15256 -14210 15316 -14150
rect 15256 -14340 15316 -14280
rect 170 -14712 230 -14652
rect 170 -14842 230 -14782
rect 626 -14712 686 -14652
rect 626 -14842 686 -14782
rect 1082 -14712 1142 -14652
rect 1082 -14842 1142 -14782
rect 1540 -14712 1600 -14652
rect 1540 -14842 1600 -14782
rect 1996 -14712 2056 -14652
rect 1996 -14842 2056 -14782
rect 2452 -14712 2512 -14652
rect 2452 -14842 2512 -14782
rect 2910 -14712 2970 -14652
rect 2910 -14842 2970 -14782
rect 3366 -14712 3426 -14652
rect 3366 -14842 3426 -14782
rect 3822 -14712 3882 -14652
rect 3822 -14842 3882 -14782
rect 4280 -14712 4340 -14652
rect 4280 -14842 4340 -14782
rect 4736 -14712 4796 -14652
rect 4736 -14842 4796 -14782
rect 5192 -14712 5252 -14652
rect 5192 -14842 5252 -14782
rect 5650 -14712 5710 -14652
rect 5650 -14842 5710 -14782
rect 6106 -14712 6166 -14652
rect 6106 -14842 6166 -14782
rect 6562 -14712 6622 -14652
rect 6562 -14842 6622 -14782
rect 7020 -14712 7080 -14652
rect 7020 -14842 7080 -14782
rect 7476 -14712 7536 -14652
rect 7476 -14842 7536 -14782
rect 7932 -14712 7992 -14652
rect 7932 -14842 7992 -14782
rect 8406 -14712 8466 -14652
rect 8406 -14842 8466 -14782
rect 8862 -14712 8922 -14652
rect 8862 -14842 8922 -14782
rect 9320 -14712 9380 -14652
rect 9320 -14842 9380 -14782
rect 9776 -14712 9836 -14652
rect 9776 -14842 9836 -14782
rect 10232 -14712 10292 -14652
rect 10232 -14842 10292 -14782
rect 10690 -14712 10750 -14652
rect 10690 -14842 10750 -14782
rect 11146 -14712 11206 -14652
rect 11146 -14842 11206 -14782
rect 11602 -14712 11662 -14652
rect 11602 -14842 11662 -14782
rect 12060 -14712 12120 -14652
rect 12060 -14842 12120 -14782
rect 12516 -14712 12576 -14652
rect 12516 -14842 12576 -14782
rect 12972 -14712 13032 -14652
rect 12972 -14842 13032 -14782
rect 13430 -14712 13490 -14652
rect 13430 -14842 13490 -14782
rect 13886 -14712 13946 -14652
rect 13886 -14842 13946 -14782
rect 14342 -14712 14402 -14652
rect 14342 -14842 14402 -14782
rect 14800 -14712 14860 -14652
rect 14800 -14842 14860 -14782
rect 15256 -14712 15316 -14652
rect 15256 -14842 15316 -14782
rect 170 -15204 230 -15144
rect 170 -15334 230 -15274
rect 626 -15204 686 -15144
rect 626 -15334 686 -15274
rect 1082 -15204 1142 -15144
rect 1082 -15334 1142 -15274
rect 1540 -15204 1600 -15144
rect 1540 -15334 1600 -15274
rect 1996 -15204 2056 -15144
rect 1996 -15334 2056 -15274
rect 2452 -15204 2512 -15144
rect 2452 -15334 2512 -15274
rect 2910 -15204 2970 -15144
rect 2910 -15334 2970 -15274
rect 3366 -15204 3426 -15144
rect 3366 -15334 3426 -15274
rect 3822 -15204 3882 -15144
rect 3822 -15334 3882 -15274
rect 4280 -15204 4340 -15144
rect 4280 -15334 4340 -15274
rect 4736 -15204 4796 -15144
rect 4736 -15334 4796 -15274
rect 5192 -15204 5252 -15144
rect 5192 -15334 5252 -15274
rect 5650 -15204 5710 -15144
rect 5650 -15334 5710 -15274
rect 6106 -15204 6166 -15144
rect 6106 -15334 6166 -15274
rect 6562 -15204 6622 -15144
rect 6562 -15334 6622 -15274
rect 7020 -15204 7080 -15144
rect 7020 -15334 7080 -15274
rect 7476 -15204 7536 -15144
rect 7476 -15334 7536 -15274
rect 7932 -15204 7992 -15144
rect 7932 -15334 7992 -15274
rect 8406 -15204 8466 -15144
rect 8406 -15334 8466 -15274
rect 8862 -15204 8922 -15144
rect 8862 -15334 8922 -15274
rect 9320 -15204 9380 -15144
rect 9320 -15334 9380 -15274
rect 9776 -15204 9836 -15144
rect 9776 -15334 9836 -15274
rect 10232 -15204 10292 -15144
rect 10232 -15334 10292 -15274
rect 10690 -15204 10750 -15144
rect 10690 -15334 10750 -15274
rect 11146 -15204 11206 -15144
rect 11146 -15334 11206 -15274
rect 11602 -15204 11662 -15144
rect 11602 -15334 11662 -15274
rect 12060 -15204 12120 -15144
rect 12060 -15334 12120 -15274
rect 12516 -15204 12576 -15144
rect 12516 -15334 12576 -15274
rect 12972 -15204 13032 -15144
rect 12972 -15334 13032 -15274
rect 13430 -15204 13490 -15144
rect 13430 -15334 13490 -15274
rect 13886 -15204 13946 -15144
rect 13886 -15334 13946 -15274
rect 14342 -15204 14402 -15144
rect 14342 -15334 14402 -15274
rect 14800 -15204 14860 -15144
rect 14800 -15334 14860 -15274
rect 15256 -15204 15316 -15144
rect 15256 -15334 15316 -15274
rect 170 -15720 230 -15660
rect 170 -15850 230 -15790
rect 626 -15720 686 -15660
rect 626 -15850 686 -15790
rect 1082 -15720 1142 -15660
rect 1082 -15850 1142 -15790
rect 1540 -15720 1600 -15660
rect 1540 -15850 1600 -15790
rect 1996 -15720 2056 -15660
rect 1996 -15850 2056 -15790
rect 2452 -15720 2512 -15660
rect 2452 -15850 2512 -15790
rect 2910 -15720 2970 -15660
rect 2910 -15850 2970 -15790
rect 3366 -15720 3426 -15660
rect 3366 -15850 3426 -15790
rect 3822 -15720 3882 -15660
rect 3822 -15850 3882 -15790
rect 4280 -15720 4340 -15660
rect 4280 -15850 4340 -15790
rect 4736 -15720 4796 -15660
rect 4736 -15850 4796 -15790
rect 5192 -15720 5252 -15660
rect 5192 -15850 5252 -15790
rect 5650 -15720 5710 -15660
rect 5650 -15850 5710 -15790
rect 6106 -15720 6166 -15660
rect 6106 -15850 6166 -15790
rect 6562 -15720 6622 -15660
rect 6562 -15850 6622 -15790
rect 7020 -15720 7080 -15660
rect 7020 -15850 7080 -15790
rect 7476 -15720 7536 -15660
rect 7476 -15850 7536 -15790
rect 7932 -15720 7992 -15660
rect 7932 -15850 7992 -15790
rect 8406 -15720 8466 -15660
rect 8406 -15850 8466 -15790
rect 8862 -15720 8922 -15660
rect 8862 -15850 8922 -15790
rect 9320 -15720 9380 -15660
rect 9320 -15850 9380 -15790
rect 9776 -15720 9836 -15660
rect 9776 -15850 9836 -15790
rect 10232 -15720 10292 -15660
rect 10232 -15850 10292 -15790
rect 10690 -15720 10750 -15660
rect 10690 -15850 10750 -15790
rect 11146 -15720 11206 -15660
rect 11146 -15850 11206 -15790
rect 11602 -15720 11662 -15660
rect 11602 -15850 11662 -15790
rect 12060 -15720 12120 -15660
rect 12060 -15850 12120 -15790
rect 12516 -15720 12576 -15660
rect 12516 -15850 12576 -15790
rect 12972 -15720 13032 -15660
rect 12972 -15850 13032 -15790
rect 13430 -15720 13490 -15660
rect 13430 -15850 13490 -15790
rect 13886 -15720 13946 -15660
rect 13886 -15850 13946 -15790
rect 14342 -15720 14402 -15660
rect 14342 -15850 14402 -15790
rect 14800 -15720 14860 -15660
rect 14800 -15850 14860 -15790
rect 15256 -15720 15316 -15660
rect 15256 -15850 15316 -15790
rect 170 -16222 230 -16162
rect 170 -16352 230 -16292
rect 626 -16222 686 -16162
rect 626 -16352 686 -16292
rect 1082 -16222 1142 -16162
rect 1082 -16352 1142 -16292
rect 1540 -16222 1600 -16162
rect 1540 -16352 1600 -16292
rect 1996 -16222 2056 -16162
rect 1996 -16352 2056 -16292
rect 2452 -16222 2512 -16162
rect 2452 -16352 2512 -16292
rect 2910 -16222 2970 -16162
rect 2910 -16352 2970 -16292
rect 3366 -16222 3426 -16162
rect 3366 -16352 3426 -16292
rect 3822 -16222 3882 -16162
rect 3822 -16352 3882 -16292
rect 4280 -16222 4340 -16162
rect 4280 -16352 4340 -16292
rect 4736 -16222 4796 -16162
rect 4736 -16352 4796 -16292
rect 5192 -16222 5252 -16162
rect 5192 -16352 5252 -16292
rect 5650 -16222 5710 -16162
rect 5650 -16352 5710 -16292
rect 6106 -16222 6166 -16162
rect 6106 -16352 6166 -16292
rect 6562 -16222 6622 -16162
rect 6562 -16352 6622 -16292
rect 7020 -16222 7080 -16162
rect 7020 -16352 7080 -16292
rect 7476 -16222 7536 -16162
rect 7476 -16352 7536 -16292
rect 7932 -16222 7992 -16162
rect 7932 -16352 7992 -16292
rect 8406 -16222 8466 -16162
rect 8406 -16352 8466 -16292
rect 8862 -16222 8922 -16162
rect 8862 -16352 8922 -16292
rect 9320 -16222 9380 -16162
rect 9320 -16352 9380 -16292
rect 9776 -16222 9836 -16162
rect 9776 -16352 9836 -16292
rect 10232 -16222 10292 -16162
rect 10232 -16352 10292 -16292
rect 10690 -16222 10750 -16162
rect 10690 -16352 10750 -16292
rect 11146 -16222 11206 -16162
rect 11146 -16352 11206 -16292
rect 11602 -16222 11662 -16162
rect 11602 -16352 11662 -16292
rect 12060 -16222 12120 -16162
rect 12060 -16352 12120 -16292
rect 12516 -16222 12576 -16162
rect 12516 -16352 12576 -16292
rect 12972 -16222 13032 -16162
rect 12972 -16352 13032 -16292
rect 13430 -16222 13490 -16162
rect 13430 -16352 13490 -16292
rect 13886 -16222 13946 -16162
rect 13886 -16352 13946 -16292
rect 14342 -16222 14402 -16162
rect 14342 -16352 14402 -16292
rect 14800 -16222 14860 -16162
rect 14800 -16352 14860 -16292
rect 15256 -16222 15316 -16162
rect 15256 -16352 15316 -16292
rect 170 -16714 230 -16654
rect 170 -16844 230 -16784
rect 626 -16714 686 -16654
rect 626 -16844 686 -16784
rect 1082 -16714 1142 -16654
rect 1082 -16844 1142 -16784
rect 1540 -16714 1600 -16654
rect 1540 -16844 1600 -16784
rect 1996 -16714 2056 -16654
rect 1996 -16844 2056 -16784
rect 2452 -16714 2512 -16654
rect 2452 -16844 2512 -16784
rect 2910 -16714 2970 -16654
rect 2910 -16844 2970 -16784
rect 3366 -16714 3426 -16654
rect 3366 -16844 3426 -16784
rect 3822 -16714 3882 -16654
rect 3822 -16844 3882 -16784
rect 4280 -16714 4340 -16654
rect 4280 -16844 4340 -16784
rect 4736 -16714 4796 -16654
rect 4736 -16844 4796 -16784
rect 5192 -16714 5252 -16654
rect 5192 -16844 5252 -16784
rect 5650 -16714 5710 -16654
rect 5650 -16844 5710 -16784
rect 6106 -16714 6166 -16654
rect 6106 -16844 6166 -16784
rect 6562 -16714 6622 -16654
rect 6562 -16844 6622 -16784
rect 7020 -16714 7080 -16654
rect 7020 -16844 7080 -16784
rect 7476 -16714 7536 -16654
rect 7476 -16844 7536 -16784
rect 7932 -16714 7992 -16654
rect 7932 -16844 7992 -16784
rect 8406 -16714 8466 -16654
rect 8406 -16844 8466 -16784
rect 8862 -16714 8922 -16654
rect 8862 -16844 8922 -16784
rect 9320 -16714 9380 -16654
rect 9320 -16844 9380 -16784
rect 9776 -16714 9836 -16654
rect 9776 -16844 9836 -16784
rect 10232 -16714 10292 -16654
rect 10232 -16844 10292 -16784
rect 10690 -16714 10750 -16654
rect 10690 -16844 10750 -16784
rect 11146 -16714 11206 -16654
rect 11146 -16844 11206 -16784
rect 11602 -16714 11662 -16654
rect 11602 -16844 11662 -16784
rect 12060 -16714 12120 -16654
rect 12060 -16844 12120 -16784
rect 12516 -16714 12576 -16654
rect 12516 -16844 12576 -16784
rect 12972 -16714 13032 -16654
rect 12972 -16844 13032 -16784
rect 13430 -16714 13490 -16654
rect 13430 -16844 13490 -16784
rect 13886 -16714 13946 -16654
rect 13886 -16844 13946 -16784
rect 14342 -16714 14402 -16654
rect 14342 -16844 14402 -16784
rect 14800 -16714 14860 -16654
rect 14800 -16844 14860 -16784
rect 15256 -16714 15316 -16654
rect 15256 -16844 15316 -16784
rect 171 -17211 231 -17151
rect 171 -17341 231 -17281
rect 627 -17211 687 -17151
rect 627 -17341 687 -17281
rect 1083 -17211 1143 -17151
rect 1083 -17341 1143 -17281
rect 1541 -17211 1601 -17151
rect 1541 -17341 1601 -17281
rect 1997 -17211 2057 -17151
rect 1997 -17341 2057 -17281
rect 2453 -17211 2513 -17151
rect 2453 -17341 2513 -17281
rect 2911 -17211 2971 -17151
rect 2911 -17341 2971 -17281
rect 3367 -17211 3427 -17151
rect 3367 -17341 3427 -17281
rect 3823 -17211 3883 -17151
rect 3823 -17341 3883 -17281
rect 4281 -17211 4341 -17151
rect 4281 -17341 4341 -17281
rect 4737 -17211 4797 -17151
rect 4737 -17341 4797 -17281
rect 5193 -17211 5253 -17151
rect 5193 -17341 5253 -17281
rect 5651 -17211 5711 -17151
rect 5651 -17341 5711 -17281
rect 6107 -17211 6167 -17151
rect 6107 -17341 6167 -17281
rect 6563 -17211 6623 -17151
rect 6563 -17341 6623 -17281
rect 7021 -17211 7081 -17151
rect 7021 -17341 7081 -17281
rect 7477 -17211 7537 -17151
rect 7477 -17341 7537 -17281
rect 7933 -17211 7993 -17151
rect 7933 -17341 7993 -17281
rect 8407 -17211 8467 -17151
rect 8407 -17341 8467 -17281
rect 8863 -17211 8923 -17151
rect 8863 -17341 8923 -17281
rect 9321 -17211 9381 -17151
rect 9321 -17341 9381 -17281
rect 9777 -17211 9837 -17151
rect 9777 -17341 9837 -17281
rect 10233 -17211 10293 -17151
rect 10233 -17341 10293 -17281
rect 10691 -17211 10751 -17151
rect 10691 -17341 10751 -17281
rect 11147 -17211 11207 -17151
rect 11147 -17341 11207 -17281
rect 11603 -17211 11663 -17151
rect 11603 -17341 11663 -17281
rect 12061 -17211 12121 -17151
rect 12061 -17341 12121 -17281
rect 12517 -17211 12577 -17151
rect 12517 -17341 12577 -17281
rect 12973 -17211 13033 -17151
rect 12973 -17341 13033 -17281
rect 13431 -17211 13491 -17151
rect 13431 -17341 13491 -17281
rect 13887 -17211 13947 -17151
rect 13887 -17341 13947 -17281
rect 14343 -17211 14403 -17151
rect 14343 -17341 14403 -17281
rect 14801 -17211 14861 -17151
rect 14801 -17341 14861 -17281
rect 15257 -17211 15317 -17151
rect 15257 -17341 15317 -17281
rect 171 -17703 231 -17643
rect 171 -17833 231 -17773
rect 627 -17703 687 -17643
rect 627 -17833 687 -17773
rect 1083 -17703 1143 -17643
rect 1083 -17833 1143 -17773
rect 1541 -17703 1601 -17643
rect 1541 -17833 1601 -17773
rect 1997 -17703 2057 -17643
rect 1997 -17833 2057 -17773
rect 2453 -17703 2513 -17643
rect 2453 -17833 2513 -17773
rect 2911 -17703 2971 -17643
rect 2911 -17833 2971 -17773
rect 3367 -17703 3427 -17643
rect 3367 -17833 3427 -17773
rect 3823 -17703 3883 -17643
rect 3823 -17833 3883 -17773
rect 4281 -17703 4341 -17643
rect 4281 -17833 4341 -17773
rect 4737 -17703 4797 -17643
rect 4737 -17833 4797 -17773
rect 5193 -17703 5253 -17643
rect 5193 -17833 5253 -17773
rect 5651 -17703 5711 -17643
rect 5651 -17833 5711 -17773
rect 6107 -17703 6167 -17643
rect 6107 -17833 6167 -17773
rect 6563 -17703 6623 -17643
rect 6563 -17833 6623 -17773
rect 7021 -17703 7081 -17643
rect 7021 -17833 7081 -17773
rect 7477 -17703 7537 -17643
rect 7477 -17833 7537 -17773
rect 7933 -17703 7993 -17643
rect 7933 -17833 7993 -17773
rect 8407 -17703 8467 -17643
rect 8407 -17833 8467 -17773
rect 8863 -17703 8923 -17643
rect 8863 -17833 8923 -17773
rect 9321 -17703 9381 -17643
rect 9321 -17833 9381 -17773
rect 9777 -17703 9837 -17643
rect 9777 -17833 9837 -17773
rect 10233 -17703 10293 -17643
rect 10233 -17833 10293 -17773
rect 10691 -17703 10751 -17643
rect 10691 -17833 10751 -17773
rect 11147 -17703 11207 -17643
rect 11147 -17833 11207 -17773
rect 11603 -17703 11663 -17643
rect 11603 -17833 11663 -17773
rect 12061 -17703 12121 -17643
rect 12061 -17833 12121 -17773
rect 12517 -17703 12577 -17643
rect 12517 -17833 12577 -17773
rect 12973 -17703 13033 -17643
rect 12973 -17833 13033 -17773
rect 13431 -17703 13491 -17643
rect 13431 -17833 13491 -17773
rect 13887 -17703 13947 -17643
rect 13887 -17833 13947 -17773
rect 14343 -17703 14403 -17643
rect 14343 -17833 14403 -17773
rect 14801 -17703 14861 -17643
rect 14801 -17833 14861 -17773
rect 15257 -17703 15317 -17643
rect 15257 -17833 15317 -17773
rect 171 -18219 231 -18159
rect 171 -18349 231 -18289
rect 627 -18219 687 -18159
rect 627 -18349 687 -18289
rect 1083 -18219 1143 -18159
rect 1083 -18349 1143 -18289
rect 1541 -18219 1601 -18159
rect 1541 -18349 1601 -18289
rect 1997 -18219 2057 -18159
rect 1997 -18349 2057 -18289
rect 2453 -18219 2513 -18159
rect 2453 -18349 2513 -18289
rect 2911 -18219 2971 -18159
rect 2911 -18349 2971 -18289
rect 3367 -18219 3427 -18159
rect 3367 -18349 3427 -18289
rect 3823 -18219 3883 -18159
rect 3823 -18349 3883 -18289
rect 4281 -18219 4341 -18159
rect 4281 -18349 4341 -18289
rect 4737 -18219 4797 -18159
rect 4737 -18349 4797 -18289
rect 5193 -18219 5253 -18159
rect 5193 -18349 5253 -18289
rect 5651 -18219 5711 -18159
rect 5651 -18349 5711 -18289
rect 6107 -18219 6167 -18159
rect 6107 -18349 6167 -18289
rect 6563 -18219 6623 -18159
rect 6563 -18349 6623 -18289
rect 7021 -18219 7081 -18159
rect 7021 -18349 7081 -18289
rect 7477 -18219 7537 -18159
rect 7477 -18349 7537 -18289
rect 7933 -18219 7993 -18159
rect 7933 -18349 7993 -18289
rect 8407 -18219 8467 -18159
rect 8407 -18349 8467 -18289
rect 8863 -18219 8923 -18159
rect 8863 -18349 8923 -18289
rect 9321 -18219 9381 -18159
rect 9321 -18349 9381 -18289
rect 9777 -18219 9837 -18159
rect 9777 -18349 9837 -18289
rect 10233 -18219 10293 -18159
rect 10233 -18349 10293 -18289
rect 10691 -18219 10751 -18159
rect 10691 -18349 10751 -18289
rect 11147 -18219 11207 -18159
rect 11147 -18349 11207 -18289
rect 11603 -18219 11663 -18159
rect 11603 -18349 11663 -18289
rect 12061 -18219 12121 -18159
rect 12061 -18349 12121 -18289
rect 12517 -18219 12577 -18159
rect 12517 -18349 12577 -18289
rect 12973 -18219 13033 -18159
rect 12973 -18349 13033 -18289
rect 13431 -18219 13491 -18159
rect 13431 -18349 13491 -18289
rect 13887 -18219 13947 -18159
rect 13887 -18349 13947 -18289
rect 14343 -18219 14403 -18159
rect 14343 -18349 14403 -18289
rect 14801 -18219 14861 -18159
rect 14801 -18349 14861 -18289
rect 15257 -18219 15317 -18159
rect 15257 -18349 15317 -18289
rect 171 -18721 231 -18661
rect 171 -18851 231 -18791
rect 627 -18721 687 -18661
rect 627 -18851 687 -18791
rect 1083 -18721 1143 -18661
rect 1083 -18851 1143 -18791
rect 1541 -18721 1601 -18661
rect 1541 -18851 1601 -18791
rect 1997 -18721 2057 -18661
rect 1997 -18851 2057 -18791
rect 2453 -18721 2513 -18661
rect 2453 -18851 2513 -18791
rect 2911 -18721 2971 -18661
rect 2911 -18851 2971 -18791
rect 3367 -18721 3427 -18661
rect 3367 -18851 3427 -18791
rect 3823 -18721 3883 -18661
rect 3823 -18851 3883 -18791
rect 4281 -18721 4341 -18661
rect 4281 -18851 4341 -18791
rect 4737 -18721 4797 -18661
rect 4737 -18851 4797 -18791
rect 5193 -18721 5253 -18661
rect 5193 -18851 5253 -18791
rect 5651 -18721 5711 -18661
rect 5651 -18851 5711 -18791
rect 6107 -18721 6167 -18661
rect 6107 -18851 6167 -18791
rect 6563 -18721 6623 -18661
rect 6563 -18851 6623 -18791
rect 7021 -18721 7081 -18661
rect 7021 -18851 7081 -18791
rect 7477 -18721 7537 -18661
rect 7477 -18851 7537 -18791
rect 7933 -18721 7993 -18661
rect 7933 -18851 7993 -18791
rect 8407 -18721 8467 -18661
rect 8407 -18851 8467 -18791
rect 8863 -18721 8923 -18661
rect 8863 -18851 8923 -18791
rect 9321 -18721 9381 -18661
rect 9321 -18851 9381 -18791
rect 9777 -18721 9837 -18661
rect 9777 -18851 9837 -18791
rect 10233 -18721 10293 -18661
rect 10233 -18851 10293 -18791
rect 10691 -18721 10751 -18661
rect 10691 -18851 10751 -18791
rect 11147 -18721 11207 -18661
rect 11147 -18851 11207 -18791
rect 11603 -18721 11663 -18661
rect 11603 -18851 11663 -18791
rect 12061 -18721 12121 -18661
rect 12061 -18851 12121 -18791
rect 12517 -18721 12577 -18661
rect 12517 -18851 12577 -18791
rect 12973 -18721 13033 -18661
rect 12973 -18851 13033 -18791
rect 13431 -18721 13491 -18661
rect 13431 -18851 13491 -18791
rect 13887 -18721 13947 -18661
rect 13887 -18851 13947 -18791
rect 14343 -18721 14403 -18661
rect 14343 -18851 14403 -18791
rect 14801 -18721 14861 -18661
rect 14801 -18851 14861 -18791
rect 15257 -18721 15317 -18661
rect 15257 -18851 15317 -18791
rect 171 -19213 231 -19153
rect 171 -19343 231 -19283
rect 627 -19213 687 -19153
rect 627 -19343 687 -19283
rect 1083 -19213 1143 -19153
rect 1083 -19343 1143 -19283
rect 1541 -19213 1601 -19153
rect 1541 -19343 1601 -19283
rect 1997 -19213 2057 -19153
rect 1997 -19343 2057 -19283
rect 2453 -19213 2513 -19153
rect 2453 -19343 2513 -19283
rect 2911 -19213 2971 -19153
rect 2911 -19343 2971 -19283
rect 3367 -19213 3427 -19153
rect 3367 -19343 3427 -19283
rect 3823 -19213 3883 -19153
rect 3823 -19343 3883 -19283
rect 4281 -19213 4341 -19153
rect 4281 -19343 4341 -19283
rect 4737 -19213 4797 -19153
rect 4737 -19343 4797 -19283
rect 5193 -19213 5253 -19153
rect 5193 -19343 5253 -19283
rect 5651 -19213 5711 -19153
rect 5651 -19343 5711 -19283
rect 6107 -19213 6167 -19153
rect 6107 -19343 6167 -19283
rect 6563 -19213 6623 -19153
rect 6563 -19343 6623 -19283
rect 7021 -19213 7081 -19153
rect 7021 -19343 7081 -19283
rect 7477 -19213 7537 -19153
rect 7477 -19343 7537 -19283
rect 7933 -19213 7993 -19153
rect 7933 -19343 7993 -19283
rect 8407 -19213 8467 -19153
rect 8407 -19343 8467 -19283
rect 8863 -19213 8923 -19153
rect 8863 -19343 8923 -19283
rect 9321 -19213 9381 -19153
rect 9321 -19343 9381 -19283
rect 9777 -19213 9837 -19153
rect 9777 -19343 9837 -19283
rect 10233 -19213 10293 -19153
rect 10233 -19343 10293 -19283
rect 10691 -19213 10751 -19153
rect 10691 -19343 10751 -19283
rect 11147 -19213 11207 -19153
rect 11147 -19343 11207 -19283
rect 11603 -19213 11663 -19153
rect 11603 -19343 11663 -19283
rect 12061 -19213 12121 -19153
rect 12061 -19343 12121 -19283
rect 12517 -19213 12577 -19153
rect 12517 -19343 12577 -19283
rect 12973 -19213 13033 -19153
rect 12973 -19343 13033 -19283
rect 13431 -19213 13491 -19153
rect 13431 -19343 13491 -19283
rect 13887 -19213 13947 -19153
rect 13887 -19343 13947 -19283
rect 14343 -19213 14403 -19153
rect 14343 -19343 14403 -19283
rect 14801 -19213 14861 -19153
rect 14801 -19343 14861 -19283
rect 15257 -19213 15317 -19153
rect 15257 -19343 15317 -19283
rect 171 -19707 231 -19647
rect 171 -19837 231 -19777
rect 627 -19707 687 -19647
rect 627 -19837 687 -19777
rect 1083 -19707 1143 -19647
rect 1083 -19837 1143 -19777
rect 1541 -19707 1601 -19647
rect 1541 -19837 1601 -19777
rect 1997 -19707 2057 -19647
rect 1997 -19837 2057 -19777
rect 2453 -19707 2513 -19647
rect 2453 -19837 2513 -19777
rect 2911 -19707 2971 -19647
rect 2911 -19837 2971 -19777
rect 3367 -19707 3427 -19647
rect 3367 -19837 3427 -19777
rect 3823 -19707 3883 -19647
rect 3823 -19837 3883 -19777
rect 4281 -19707 4341 -19647
rect 4281 -19837 4341 -19777
rect 4737 -19707 4797 -19647
rect 4737 -19837 4797 -19777
rect 5193 -19707 5253 -19647
rect 5193 -19837 5253 -19777
rect 5651 -19707 5711 -19647
rect 5651 -19837 5711 -19777
rect 6107 -19707 6167 -19647
rect 6107 -19837 6167 -19777
rect 6563 -19707 6623 -19647
rect 6563 -19837 6623 -19777
rect 7021 -19707 7081 -19647
rect 7021 -19837 7081 -19777
rect 7477 -19707 7537 -19647
rect 7477 -19837 7537 -19777
rect 7933 -19707 7993 -19647
rect 7933 -19837 7993 -19777
rect 8407 -19707 8467 -19647
rect 8407 -19837 8467 -19777
rect 8863 -19707 8923 -19647
rect 8863 -19837 8923 -19777
rect 9321 -19707 9381 -19647
rect 9321 -19837 9381 -19777
rect 9777 -19707 9837 -19647
rect 9777 -19837 9837 -19777
rect 10233 -19707 10293 -19647
rect 10233 -19837 10293 -19777
rect 10691 -19707 10751 -19647
rect 10691 -19837 10751 -19777
rect 11147 -19707 11207 -19647
rect 11147 -19837 11207 -19777
rect 11603 -19707 11663 -19647
rect 11603 -19837 11663 -19777
rect 12061 -19707 12121 -19647
rect 12061 -19837 12121 -19777
rect 12517 -19707 12577 -19647
rect 12517 -19837 12577 -19777
rect 12973 -19707 13033 -19647
rect 12973 -19837 13033 -19777
rect 13431 -19707 13491 -19647
rect 13431 -19837 13491 -19777
rect 13887 -19707 13947 -19647
rect 13887 -19837 13947 -19777
rect 14343 -19707 14403 -19647
rect 14343 -19837 14403 -19777
rect 14801 -19707 14861 -19647
rect 14801 -19837 14861 -19777
rect 15257 -19707 15317 -19647
rect 15257 -19837 15317 -19777
rect 171 -20209 231 -20149
rect 171 -20339 231 -20279
rect 627 -20209 687 -20149
rect 627 -20339 687 -20279
rect 1083 -20209 1143 -20149
rect 1083 -20339 1143 -20279
rect 1541 -20209 1601 -20149
rect 1541 -20339 1601 -20279
rect 1997 -20209 2057 -20149
rect 1997 -20339 2057 -20279
rect 2453 -20209 2513 -20149
rect 2453 -20339 2513 -20279
rect 2911 -20209 2971 -20149
rect 2911 -20339 2971 -20279
rect 3367 -20209 3427 -20149
rect 3367 -20339 3427 -20279
rect 3823 -20209 3883 -20149
rect 3823 -20339 3883 -20279
rect 4281 -20209 4341 -20149
rect 4281 -20339 4341 -20279
rect 4737 -20209 4797 -20149
rect 4737 -20339 4797 -20279
rect 5193 -20209 5253 -20149
rect 5193 -20339 5253 -20279
rect 5651 -20209 5711 -20149
rect 5651 -20339 5711 -20279
rect 6107 -20209 6167 -20149
rect 6107 -20339 6167 -20279
rect 6563 -20209 6623 -20149
rect 6563 -20339 6623 -20279
rect 7021 -20209 7081 -20149
rect 7021 -20339 7081 -20279
rect 7477 -20209 7537 -20149
rect 7477 -20339 7537 -20279
rect 7933 -20209 7993 -20149
rect 7933 -20339 7993 -20279
rect 8407 -20209 8467 -20149
rect 8407 -20339 8467 -20279
rect 8863 -20209 8923 -20149
rect 8863 -20339 8923 -20279
rect 9321 -20209 9381 -20149
rect 9321 -20339 9381 -20279
rect 9777 -20209 9837 -20149
rect 9777 -20339 9837 -20279
rect 10233 -20209 10293 -20149
rect 10233 -20339 10293 -20279
rect 10691 -20209 10751 -20149
rect 10691 -20339 10751 -20279
rect 11147 -20209 11207 -20149
rect 11147 -20339 11207 -20279
rect 11603 -20209 11663 -20149
rect 11603 -20339 11663 -20279
rect 12061 -20209 12121 -20149
rect 12061 -20339 12121 -20279
rect 12517 -20209 12577 -20149
rect 12517 -20339 12577 -20279
rect 12973 -20209 13033 -20149
rect 12973 -20339 13033 -20279
rect 13431 -20209 13491 -20149
rect 13431 -20339 13491 -20279
rect 13887 -20209 13947 -20149
rect 13887 -20339 13947 -20279
rect 14343 -20209 14403 -20149
rect 14343 -20339 14403 -20279
rect 14801 -20209 14861 -20149
rect 14801 -20339 14861 -20279
rect 15257 -20209 15317 -20149
rect 15257 -20339 15317 -20279
rect 171 -20701 231 -20641
rect 171 -20831 231 -20771
rect 627 -20701 687 -20641
rect 627 -20831 687 -20771
rect 1083 -20701 1143 -20641
rect 1083 -20831 1143 -20771
rect 1541 -20701 1601 -20641
rect 1541 -20831 1601 -20771
rect 1997 -20701 2057 -20641
rect 1997 -20831 2057 -20771
rect 2453 -20701 2513 -20641
rect 2453 -20831 2513 -20771
rect 2911 -20701 2971 -20641
rect 2911 -20831 2971 -20771
rect 3367 -20701 3427 -20641
rect 3367 -20831 3427 -20771
rect 3823 -20701 3883 -20641
rect 3823 -20831 3883 -20771
rect 4281 -20701 4341 -20641
rect 4281 -20831 4341 -20771
rect 4737 -20701 4797 -20641
rect 4737 -20831 4797 -20771
rect 5193 -20701 5253 -20641
rect 5193 -20831 5253 -20771
rect 5651 -20701 5711 -20641
rect 5651 -20831 5711 -20771
rect 6107 -20701 6167 -20641
rect 6107 -20831 6167 -20771
rect 6563 -20701 6623 -20641
rect 6563 -20831 6623 -20771
rect 7021 -20701 7081 -20641
rect 7021 -20831 7081 -20771
rect 7477 -20701 7537 -20641
rect 7477 -20831 7537 -20771
rect 7933 -20701 7993 -20641
rect 7933 -20831 7993 -20771
rect 8407 -20701 8467 -20641
rect 8407 -20831 8467 -20771
rect 8863 -20701 8923 -20641
rect 8863 -20831 8923 -20771
rect 9321 -20701 9381 -20641
rect 9321 -20831 9381 -20771
rect 9777 -20701 9837 -20641
rect 9777 -20831 9837 -20771
rect 10233 -20701 10293 -20641
rect 10233 -20831 10293 -20771
rect 10691 -20701 10751 -20641
rect 10691 -20831 10751 -20771
rect 11147 -20701 11207 -20641
rect 11147 -20831 11207 -20771
rect 11603 -20701 11663 -20641
rect 11603 -20831 11663 -20771
rect 12061 -20701 12121 -20641
rect 12061 -20831 12121 -20771
rect 12517 -20701 12577 -20641
rect 12517 -20831 12577 -20771
rect 12973 -20701 13033 -20641
rect 12973 -20831 13033 -20771
rect 13431 -20701 13491 -20641
rect 13431 -20831 13491 -20771
rect 13887 -20701 13947 -20641
rect 13887 -20831 13947 -20771
rect 14343 -20701 14403 -20641
rect 14343 -20831 14403 -20771
rect 14801 -20701 14861 -20641
rect 14801 -20831 14861 -20771
rect 15257 -20701 15317 -20641
rect 15257 -20831 15317 -20771
rect 171 -21217 231 -21157
rect 171 -21347 231 -21287
rect 627 -21217 687 -21157
rect 627 -21347 687 -21287
rect 1083 -21217 1143 -21157
rect 1083 -21347 1143 -21287
rect 1541 -21217 1601 -21157
rect 1541 -21347 1601 -21287
rect 1997 -21217 2057 -21157
rect 1997 -21347 2057 -21287
rect 2453 -21217 2513 -21157
rect 2453 -21347 2513 -21287
rect 2911 -21217 2971 -21157
rect 2911 -21347 2971 -21287
rect 3367 -21217 3427 -21157
rect 3367 -21347 3427 -21287
rect 3823 -21217 3883 -21157
rect 3823 -21347 3883 -21287
rect 4281 -21217 4341 -21157
rect 4281 -21347 4341 -21287
rect 4737 -21217 4797 -21157
rect 4737 -21347 4797 -21287
rect 5193 -21217 5253 -21157
rect 5193 -21347 5253 -21287
rect 5651 -21217 5711 -21157
rect 5651 -21347 5711 -21287
rect 6107 -21217 6167 -21157
rect 6107 -21347 6167 -21287
rect 6563 -21217 6623 -21157
rect 6563 -21347 6623 -21287
rect 7021 -21217 7081 -21157
rect 7021 -21347 7081 -21287
rect 7477 -21217 7537 -21157
rect 7477 -21347 7537 -21287
rect 7933 -21217 7993 -21157
rect 7933 -21347 7993 -21287
rect 8407 -21217 8467 -21157
rect 8407 -21347 8467 -21287
rect 8863 -21217 8923 -21157
rect 8863 -21347 8923 -21287
rect 9321 -21217 9381 -21157
rect 9321 -21347 9381 -21287
rect 9777 -21217 9837 -21157
rect 9777 -21347 9837 -21287
rect 10233 -21217 10293 -21157
rect 10233 -21347 10293 -21287
rect 10691 -21217 10751 -21157
rect 10691 -21347 10751 -21287
rect 11147 -21217 11207 -21157
rect 11147 -21347 11207 -21287
rect 11603 -21217 11663 -21157
rect 11603 -21347 11663 -21287
rect 12061 -21217 12121 -21157
rect 12061 -21347 12121 -21287
rect 12517 -21217 12577 -21157
rect 12517 -21347 12577 -21287
rect 12973 -21217 13033 -21157
rect 12973 -21347 13033 -21287
rect 13431 -21217 13491 -21157
rect 13431 -21347 13491 -21287
rect 13887 -21217 13947 -21157
rect 13887 -21347 13947 -21287
rect 14343 -21217 14403 -21157
rect 14343 -21347 14403 -21287
rect 14801 -21217 14861 -21157
rect 14801 -21347 14861 -21287
rect 15257 -21217 15317 -21157
rect 15257 -21347 15317 -21287
rect 171 -21719 231 -21659
rect 171 -21849 231 -21789
rect 627 -21719 687 -21659
rect 627 -21849 687 -21789
rect 1083 -21719 1143 -21659
rect 1083 -21849 1143 -21789
rect 1541 -21719 1601 -21659
rect 1541 -21849 1601 -21789
rect 1997 -21719 2057 -21659
rect 1997 -21849 2057 -21789
rect 2453 -21719 2513 -21659
rect 2453 -21849 2513 -21789
rect 2911 -21719 2971 -21659
rect 2911 -21849 2971 -21789
rect 3367 -21719 3427 -21659
rect 3367 -21849 3427 -21789
rect 3823 -21719 3883 -21659
rect 3823 -21849 3883 -21789
rect 4281 -21719 4341 -21659
rect 4281 -21849 4341 -21789
rect 4737 -21719 4797 -21659
rect 4737 -21849 4797 -21789
rect 5193 -21719 5253 -21659
rect 5193 -21849 5253 -21789
rect 5651 -21719 5711 -21659
rect 5651 -21849 5711 -21789
rect 6107 -21719 6167 -21659
rect 6107 -21849 6167 -21789
rect 6563 -21719 6623 -21659
rect 6563 -21849 6623 -21789
rect 7021 -21719 7081 -21659
rect 7021 -21849 7081 -21789
rect 7477 -21719 7537 -21659
rect 7477 -21849 7537 -21789
rect 7933 -21719 7993 -21659
rect 7933 -21849 7993 -21789
rect 8407 -21719 8467 -21659
rect 8407 -21849 8467 -21789
rect 8863 -21719 8923 -21659
rect 8863 -21849 8923 -21789
rect 9321 -21719 9381 -21659
rect 9321 -21849 9381 -21789
rect 9777 -21719 9837 -21659
rect 9777 -21849 9837 -21789
rect 10233 -21719 10293 -21659
rect 10233 -21849 10293 -21789
rect 10691 -21719 10751 -21659
rect 10691 -21849 10751 -21789
rect 11147 -21719 11207 -21659
rect 11147 -21849 11207 -21789
rect 11603 -21719 11663 -21659
rect 11603 -21849 11663 -21789
rect 12061 -21719 12121 -21659
rect 12061 -21849 12121 -21789
rect 12517 -21719 12577 -21659
rect 12517 -21849 12577 -21789
rect 12973 -21719 13033 -21659
rect 12973 -21849 13033 -21789
rect 13431 -21719 13491 -21659
rect 13431 -21849 13491 -21789
rect 13887 -21719 13947 -21659
rect 13887 -21849 13947 -21789
rect 14343 -21719 14403 -21659
rect 14343 -21849 14403 -21789
rect 14801 -21719 14861 -21659
rect 14801 -21849 14861 -21789
rect 15257 -21719 15317 -21659
rect 15257 -21849 15317 -21789
rect 171 -22211 231 -22151
rect 171 -22341 231 -22281
rect 627 -22211 687 -22151
rect 627 -22341 687 -22281
rect 1083 -22211 1143 -22151
rect 1083 -22341 1143 -22281
rect 1541 -22211 1601 -22151
rect 1541 -22341 1601 -22281
rect 1997 -22211 2057 -22151
rect 1997 -22341 2057 -22281
rect 2453 -22211 2513 -22151
rect 2453 -22341 2513 -22281
rect 2911 -22211 2971 -22151
rect 2911 -22341 2971 -22281
rect 3367 -22211 3427 -22151
rect 3367 -22341 3427 -22281
rect 3823 -22211 3883 -22151
rect 3823 -22341 3883 -22281
rect 4281 -22211 4341 -22151
rect 4281 -22341 4341 -22281
rect 4737 -22211 4797 -22151
rect 4737 -22341 4797 -22281
rect 5193 -22211 5253 -22151
rect 5193 -22341 5253 -22281
rect 5651 -22211 5711 -22151
rect 5651 -22341 5711 -22281
rect 6107 -22211 6167 -22151
rect 6107 -22341 6167 -22281
rect 6563 -22211 6623 -22151
rect 6563 -22341 6623 -22281
rect 7021 -22211 7081 -22151
rect 7021 -22341 7081 -22281
rect 7477 -22211 7537 -22151
rect 7477 -22341 7537 -22281
rect 7933 -22211 7993 -22151
rect 7933 -22341 7993 -22281
rect 8407 -22211 8467 -22151
rect 8407 -22341 8467 -22281
rect 8863 -22211 8923 -22151
rect 8863 -22341 8923 -22281
rect 9321 -22211 9381 -22151
rect 9321 -22341 9381 -22281
rect 9777 -22211 9837 -22151
rect 9777 -22341 9837 -22281
rect 10233 -22211 10293 -22151
rect 10233 -22341 10293 -22281
rect 10691 -22211 10751 -22151
rect 10691 -22341 10751 -22281
rect 11147 -22211 11207 -22151
rect 11147 -22341 11207 -22281
rect 11603 -22211 11663 -22151
rect 11603 -22341 11663 -22281
rect 12061 -22211 12121 -22151
rect 12061 -22341 12121 -22281
rect 12517 -22211 12577 -22151
rect 12517 -22341 12577 -22281
rect 12973 -22211 13033 -22151
rect 12973 -22341 13033 -22281
rect 13431 -22211 13491 -22151
rect 13431 -22341 13491 -22281
rect 13887 -22211 13947 -22151
rect 13887 -22341 13947 -22281
rect 14343 -22211 14403 -22151
rect 14343 -22341 14403 -22281
rect 14801 -22211 14861 -22151
rect 14801 -22341 14861 -22281
rect 15257 -22211 15317 -22151
rect 15257 -22341 15317 -22281
rect 171 -22698 231 -22638
rect 171 -22828 231 -22768
rect 627 -22698 687 -22638
rect 627 -22828 687 -22768
rect 1083 -22698 1143 -22638
rect 1083 -22828 1143 -22768
rect 1541 -22698 1601 -22638
rect 1541 -22828 1601 -22768
rect 1997 -22698 2057 -22638
rect 1997 -22828 2057 -22768
rect 2453 -22698 2513 -22638
rect 2453 -22828 2513 -22768
rect 2911 -22698 2971 -22638
rect 2911 -22828 2971 -22768
rect 3367 -22698 3427 -22638
rect 3367 -22828 3427 -22768
rect 3823 -22698 3883 -22638
rect 3823 -22828 3883 -22768
rect 4281 -22698 4341 -22638
rect 4281 -22828 4341 -22768
rect 4737 -22698 4797 -22638
rect 4737 -22828 4797 -22768
rect 5193 -22698 5253 -22638
rect 5193 -22828 5253 -22768
rect 5651 -22698 5711 -22638
rect 5651 -22828 5711 -22768
rect 6107 -22698 6167 -22638
rect 6107 -22828 6167 -22768
rect 6563 -22698 6623 -22638
rect 6563 -22828 6623 -22768
rect 7021 -22698 7081 -22638
rect 7021 -22828 7081 -22768
rect 7477 -22698 7537 -22638
rect 7477 -22828 7537 -22768
rect 7933 -22698 7993 -22638
rect 7933 -22828 7993 -22768
rect 8407 -22698 8467 -22638
rect 8407 -22828 8467 -22768
rect 8863 -22698 8923 -22638
rect 8863 -22828 8923 -22768
rect 9321 -22698 9381 -22638
rect 9321 -22828 9381 -22768
rect 9777 -22698 9837 -22638
rect 9777 -22828 9837 -22768
rect 10233 -22698 10293 -22638
rect 10233 -22828 10293 -22768
rect 10691 -22698 10751 -22638
rect 10691 -22828 10751 -22768
rect 11147 -22698 11207 -22638
rect 11147 -22828 11207 -22768
rect 11603 -22698 11663 -22638
rect 11603 -22828 11663 -22768
rect 12061 -22698 12121 -22638
rect 12061 -22828 12121 -22768
rect 12517 -22698 12577 -22638
rect 12517 -22828 12577 -22768
rect 12973 -22698 13033 -22638
rect 12973 -22828 13033 -22768
rect 13431 -22698 13491 -22638
rect 13431 -22828 13491 -22768
rect 13887 -22698 13947 -22638
rect 13887 -22828 13947 -22768
rect 14343 -22698 14403 -22638
rect 14343 -22828 14403 -22768
rect 14801 -22698 14861 -22638
rect 14801 -22828 14861 -22768
rect 15257 -22698 15317 -22638
rect 15257 -22828 15317 -22768
rect 171 -23200 231 -23140
rect 171 -23330 231 -23270
rect 627 -23200 687 -23140
rect 627 -23330 687 -23270
rect 1083 -23200 1143 -23140
rect 1083 -23330 1143 -23270
rect 1541 -23200 1601 -23140
rect 1541 -23330 1601 -23270
rect 1997 -23200 2057 -23140
rect 1997 -23330 2057 -23270
rect 2453 -23200 2513 -23140
rect 2453 -23330 2513 -23270
rect 2911 -23200 2971 -23140
rect 2911 -23330 2971 -23270
rect 3367 -23200 3427 -23140
rect 3367 -23330 3427 -23270
rect 3823 -23200 3883 -23140
rect 3823 -23330 3883 -23270
rect 4281 -23200 4341 -23140
rect 4281 -23330 4341 -23270
rect 4737 -23200 4797 -23140
rect 4737 -23330 4797 -23270
rect 5193 -23200 5253 -23140
rect 5193 -23330 5253 -23270
rect 5651 -23200 5711 -23140
rect 5651 -23330 5711 -23270
rect 6107 -23200 6167 -23140
rect 6107 -23330 6167 -23270
rect 6563 -23200 6623 -23140
rect 6563 -23330 6623 -23270
rect 7021 -23200 7081 -23140
rect 7021 -23330 7081 -23270
rect 7477 -23200 7537 -23140
rect 7477 -23330 7537 -23270
rect 7933 -23200 7993 -23140
rect 7933 -23330 7993 -23270
rect 8407 -23200 8467 -23140
rect 8407 -23330 8467 -23270
rect 8863 -23200 8923 -23140
rect 8863 -23330 8923 -23270
rect 9321 -23200 9381 -23140
rect 9321 -23330 9381 -23270
rect 9777 -23200 9837 -23140
rect 9777 -23330 9837 -23270
rect 10233 -23200 10293 -23140
rect 10233 -23330 10293 -23270
rect 10691 -23200 10751 -23140
rect 10691 -23330 10751 -23270
rect 11147 -23200 11207 -23140
rect 11147 -23330 11207 -23270
rect 11603 -23200 11663 -23140
rect 11603 -23330 11663 -23270
rect 12061 -23200 12121 -23140
rect 12061 -23330 12121 -23270
rect 12517 -23200 12577 -23140
rect 12517 -23330 12577 -23270
rect 12973 -23200 13033 -23140
rect 12973 -23330 13033 -23270
rect 13431 -23200 13491 -23140
rect 13431 -23330 13491 -23270
rect 13887 -23200 13947 -23140
rect 13887 -23330 13947 -23270
rect 14343 -23200 14403 -23140
rect 14343 -23330 14403 -23270
rect 14801 -23200 14861 -23140
rect 14801 -23330 14861 -23270
rect 15257 -23200 15317 -23140
rect 15257 -23330 15317 -23270
rect 171 -23694 231 -23634
rect 171 -23824 231 -23764
rect 627 -23694 687 -23634
rect 627 -23824 687 -23764
rect 1083 -23694 1143 -23634
rect 1083 -23824 1143 -23764
rect 1541 -23694 1601 -23634
rect 1541 -23824 1601 -23764
rect 1997 -23694 2057 -23634
rect 1997 -23824 2057 -23764
rect 2453 -23694 2513 -23634
rect 2453 -23824 2513 -23764
rect 2911 -23694 2971 -23634
rect 2911 -23824 2971 -23764
rect 3367 -23694 3427 -23634
rect 3367 -23824 3427 -23764
rect 3823 -23694 3883 -23634
rect 3823 -23824 3883 -23764
rect 4281 -23694 4341 -23634
rect 4281 -23824 4341 -23764
rect 4737 -23694 4797 -23634
rect 4737 -23824 4797 -23764
rect 5193 -23694 5253 -23634
rect 5193 -23824 5253 -23764
rect 5651 -23694 5711 -23634
rect 5651 -23824 5711 -23764
rect 6107 -23694 6167 -23634
rect 6107 -23824 6167 -23764
rect 6563 -23694 6623 -23634
rect 6563 -23824 6623 -23764
rect 7021 -23694 7081 -23634
rect 7021 -23824 7081 -23764
rect 7477 -23694 7537 -23634
rect 7477 -23824 7537 -23764
rect 7933 -23694 7993 -23634
rect 7933 -23824 7993 -23764
rect 8407 -23694 8467 -23634
rect 8407 -23824 8467 -23764
rect 8863 -23694 8923 -23634
rect 8863 -23824 8923 -23764
rect 9321 -23694 9381 -23634
rect 9321 -23824 9381 -23764
rect 9777 -23694 9837 -23634
rect 9777 -23824 9837 -23764
rect 10233 -23694 10293 -23634
rect 10233 -23824 10293 -23764
rect 10691 -23694 10751 -23634
rect 10691 -23824 10751 -23764
rect 11147 -23694 11207 -23634
rect 11147 -23824 11207 -23764
rect 11603 -23694 11663 -23634
rect 11603 -23824 11663 -23764
rect 12061 -23694 12121 -23634
rect 12061 -23824 12121 -23764
rect 12517 -23694 12577 -23634
rect 12517 -23824 12577 -23764
rect 12973 -23694 13033 -23634
rect 12973 -23824 13033 -23764
rect 13431 -23694 13491 -23634
rect 13431 -23824 13491 -23764
rect 13887 -23694 13947 -23634
rect 13887 -23824 13947 -23764
rect 14343 -23694 14403 -23634
rect 14343 -23824 14403 -23764
rect 14801 -23694 14861 -23634
rect 14801 -23824 14861 -23764
rect 15257 -23694 15317 -23634
rect 15257 -23824 15317 -23764
rect 171 -24186 231 -24126
rect 171 -24316 231 -24256
rect 627 -24186 687 -24126
rect 627 -24316 687 -24256
rect 1083 -24186 1143 -24126
rect 1083 -24316 1143 -24256
rect 1541 -24186 1601 -24126
rect 1541 -24316 1601 -24256
rect 1997 -24186 2057 -24126
rect 1997 -24316 2057 -24256
rect 2453 -24186 2513 -24126
rect 2453 -24316 2513 -24256
rect 2911 -24186 2971 -24126
rect 2911 -24316 2971 -24256
rect 3367 -24186 3427 -24126
rect 3367 -24316 3427 -24256
rect 3823 -24186 3883 -24126
rect 3823 -24316 3883 -24256
rect 4281 -24186 4341 -24126
rect 4281 -24316 4341 -24256
rect 4737 -24186 4797 -24126
rect 4737 -24316 4797 -24256
rect 5193 -24186 5253 -24126
rect 5193 -24316 5253 -24256
rect 5651 -24186 5711 -24126
rect 5651 -24316 5711 -24256
rect 6107 -24186 6167 -24126
rect 6107 -24316 6167 -24256
rect 6563 -24186 6623 -24126
rect 6563 -24316 6623 -24256
rect 7021 -24186 7081 -24126
rect 7021 -24316 7081 -24256
rect 7477 -24186 7537 -24126
rect 7477 -24316 7537 -24256
rect 7933 -24186 7993 -24126
rect 7933 -24316 7993 -24256
rect 8407 -24186 8467 -24126
rect 8407 -24316 8467 -24256
rect 8863 -24186 8923 -24126
rect 8863 -24316 8923 -24256
rect 9321 -24186 9381 -24126
rect 9321 -24316 9381 -24256
rect 9777 -24186 9837 -24126
rect 9777 -24316 9837 -24256
rect 10233 -24186 10293 -24126
rect 10233 -24316 10293 -24256
rect 10691 -24186 10751 -24126
rect 10691 -24316 10751 -24256
rect 11147 -24186 11207 -24126
rect 11147 -24316 11207 -24256
rect 11603 -24186 11663 -24126
rect 11603 -24316 11663 -24256
rect 12061 -24186 12121 -24126
rect 12061 -24316 12121 -24256
rect 12517 -24186 12577 -24126
rect 12517 -24316 12577 -24256
rect 12973 -24186 13033 -24126
rect 12973 -24316 13033 -24256
rect 13431 -24186 13491 -24126
rect 13431 -24316 13491 -24256
rect 13887 -24186 13947 -24126
rect 13887 -24316 13947 -24256
rect 14343 -24186 14403 -24126
rect 14343 -24316 14403 -24256
rect 14801 -24186 14861 -24126
rect 14801 -24316 14861 -24256
rect 15257 -24186 15317 -24126
rect 15257 -24316 15317 -24256
rect 171 -24688 231 -24628
rect 171 -24818 231 -24758
rect 627 -24688 687 -24628
rect 627 -24818 687 -24758
rect 1083 -24688 1143 -24628
rect 1083 -24818 1143 -24758
rect 1541 -24688 1601 -24628
rect 1541 -24818 1601 -24758
rect 1997 -24688 2057 -24628
rect 1997 -24818 2057 -24758
rect 2453 -24688 2513 -24628
rect 2453 -24818 2513 -24758
rect 2911 -24688 2971 -24628
rect 2911 -24818 2971 -24758
rect 3367 -24688 3427 -24628
rect 3367 -24818 3427 -24758
rect 3823 -24688 3883 -24628
rect 3823 -24818 3883 -24758
rect 4281 -24688 4341 -24628
rect 4281 -24818 4341 -24758
rect 4737 -24688 4797 -24628
rect 4737 -24818 4797 -24758
rect 5193 -24688 5253 -24628
rect 5193 -24818 5253 -24758
rect 5651 -24688 5711 -24628
rect 5651 -24818 5711 -24758
rect 6107 -24688 6167 -24628
rect 6107 -24818 6167 -24758
rect 6563 -24688 6623 -24628
rect 6563 -24818 6623 -24758
rect 7021 -24688 7081 -24628
rect 7021 -24818 7081 -24758
rect 7477 -24688 7537 -24628
rect 7477 -24818 7537 -24758
rect 7933 -24688 7993 -24628
rect 7933 -24818 7993 -24758
rect 8407 -24688 8467 -24628
rect 8407 -24818 8467 -24758
rect 8863 -24688 8923 -24628
rect 8863 -24818 8923 -24758
rect 9321 -24688 9381 -24628
rect 9321 -24818 9381 -24758
rect 9777 -24688 9837 -24628
rect 9777 -24818 9837 -24758
rect 10233 -24688 10293 -24628
rect 10233 -24818 10293 -24758
rect 10691 -24688 10751 -24628
rect 10691 -24818 10751 -24758
rect 11147 -24688 11207 -24628
rect 11147 -24818 11207 -24758
rect 11603 -24688 11663 -24628
rect 11603 -24818 11663 -24758
rect 12061 -24688 12121 -24628
rect 12061 -24818 12121 -24758
rect 12517 -24688 12577 -24628
rect 12517 -24818 12577 -24758
rect 12973 -24688 13033 -24628
rect 12973 -24818 13033 -24758
rect 13431 -24688 13491 -24628
rect 13431 -24818 13491 -24758
rect 13887 -24688 13947 -24628
rect 13887 -24818 13947 -24758
rect 14343 -24688 14403 -24628
rect 14343 -24818 14403 -24758
rect 14801 -24688 14861 -24628
rect 14801 -24818 14861 -24758
rect 15257 -24688 15317 -24628
rect 15257 -24818 15317 -24758
rect 171 -25204 231 -25144
rect 171 -25334 231 -25274
rect 627 -25204 687 -25144
rect 627 -25334 687 -25274
rect 1083 -25204 1143 -25144
rect 1083 -25334 1143 -25274
rect 1541 -25204 1601 -25144
rect 1541 -25334 1601 -25274
rect 1997 -25204 2057 -25144
rect 1997 -25334 2057 -25274
rect 2453 -25204 2513 -25144
rect 2453 -25334 2513 -25274
rect 2911 -25204 2971 -25144
rect 2911 -25334 2971 -25274
rect 3367 -25204 3427 -25144
rect 3367 -25334 3427 -25274
rect 3823 -25204 3883 -25144
rect 3823 -25334 3883 -25274
rect 4281 -25204 4341 -25144
rect 4281 -25334 4341 -25274
rect 4737 -25204 4797 -25144
rect 4737 -25334 4797 -25274
rect 5193 -25204 5253 -25144
rect 5193 -25334 5253 -25274
rect 5651 -25204 5711 -25144
rect 5651 -25334 5711 -25274
rect 6107 -25204 6167 -25144
rect 6107 -25334 6167 -25274
rect 6563 -25204 6623 -25144
rect 6563 -25334 6623 -25274
rect 7021 -25204 7081 -25144
rect 7021 -25334 7081 -25274
rect 7477 -25204 7537 -25144
rect 7477 -25334 7537 -25274
rect 7933 -25204 7993 -25144
rect 7933 -25334 7993 -25274
rect 8407 -25204 8467 -25144
rect 8407 -25334 8467 -25274
rect 8863 -25204 8923 -25144
rect 8863 -25334 8923 -25274
rect 9321 -25204 9381 -25144
rect 9321 -25334 9381 -25274
rect 9777 -25204 9837 -25144
rect 9777 -25334 9837 -25274
rect 10233 -25204 10293 -25144
rect 10233 -25334 10293 -25274
rect 10691 -25204 10751 -25144
rect 10691 -25334 10751 -25274
rect 11147 -25204 11207 -25144
rect 11147 -25334 11207 -25274
rect 11603 -25204 11663 -25144
rect 11603 -25334 11663 -25274
rect 12061 -25204 12121 -25144
rect 12061 -25334 12121 -25274
rect 12517 -25204 12577 -25144
rect 12517 -25334 12577 -25274
rect 12973 -25204 13033 -25144
rect 12973 -25334 13033 -25274
rect 13431 -25204 13491 -25144
rect 13431 -25334 13491 -25274
rect 13887 -25204 13947 -25144
rect 13887 -25334 13947 -25274
rect 14343 -25204 14403 -25144
rect 14343 -25334 14403 -25274
rect 14801 -25204 14861 -25144
rect 14801 -25334 14861 -25274
rect 15257 -25204 15317 -25144
rect 15257 -25334 15317 -25274
rect 171 -25696 231 -25636
rect 171 -25826 231 -25766
rect 627 -25696 687 -25636
rect 627 -25826 687 -25766
rect 1083 -25696 1143 -25636
rect 1083 -25826 1143 -25766
rect 1541 -25696 1601 -25636
rect 1541 -25826 1601 -25766
rect 1997 -25696 2057 -25636
rect 1997 -25826 2057 -25766
rect 2453 -25696 2513 -25636
rect 2453 -25826 2513 -25766
rect 2911 -25696 2971 -25636
rect 2911 -25826 2971 -25766
rect 3367 -25696 3427 -25636
rect 3367 -25826 3427 -25766
rect 3823 -25696 3883 -25636
rect 3823 -25826 3883 -25766
rect 4281 -25696 4341 -25636
rect 4281 -25826 4341 -25766
rect 4737 -25696 4797 -25636
rect 4737 -25826 4797 -25766
rect 5193 -25696 5253 -25636
rect 5193 -25826 5253 -25766
rect 5651 -25696 5711 -25636
rect 5651 -25826 5711 -25766
rect 6107 -25696 6167 -25636
rect 6107 -25826 6167 -25766
rect 6563 -25696 6623 -25636
rect 6563 -25826 6623 -25766
rect 7021 -25696 7081 -25636
rect 7021 -25826 7081 -25766
rect 7477 -25696 7537 -25636
rect 7477 -25826 7537 -25766
rect 7933 -25696 7993 -25636
rect 7933 -25826 7993 -25766
rect 8407 -25696 8467 -25636
rect 8407 -25826 8467 -25766
rect 8863 -25696 8923 -25636
rect 8863 -25826 8923 -25766
rect 9321 -25696 9381 -25636
rect 9321 -25826 9381 -25766
rect 9777 -25696 9837 -25636
rect 9777 -25826 9837 -25766
rect 10233 -25696 10293 -25636
rect 10233 -25826 10293 -25766
rect 10691 -25696 10751 -25636
rect 10691 -25826 10751 -25766
rect 11147 -25696 11207 -25636
rect 11147 -25826 11207 -25766
rect 11603 -25696 11663 -25636
rect 11603 -25826 11663 -25766
rect 12061 -25696 12121 -25636
rect 12061 -25826 12121 -25766
rect 12517 -25696 12577 -25636
rect 12517 -25826 12577 -25766
rect 12973 -25696 13033 -25636
rect 12973 -25826 13033 -25766
rect 13431 -25696 13491 -25636
rect 13431 -25826 13491 -25766
rect 13887 -25696 13947 -25636
rect 13887 -25826 13947 -25766
rect 14343 -25696 14403 -25636
rect 14343 -25826 14403 -25766
rect 14801 -25696 14861 -25636
rect 14801 -25826 14861 -25766
rect 15257 -25696 15317 -25636
rect 15257 -25826 15317 -25766
rect 170 -26193 230 -26133
rect 170 -26323 230 -26263
rect 626 -26193 686 -26133
rect 626 -26323 686 -26263
rect 1082 -26193 1142 -26133
rect 1082 -26323 1142 -26263
rect 1540 -26193 1600 -26133
rect 1540 -26323 1600 -26263
rect 1996 -26193 2056 -26133
rect 1996 -26323 2056 -26263
rect 2452 -26193 2512 -26133
rect 2452 -26323 2512 -26263
rect 2910 -26193 2970 -26133
rect 2910 -26323 2970 -26263
rect 3366 -26193 3426 -26133
rect 3366 -26323 3426 -26263
rect 3822 -26193 3882 -26133
rect 3822 -26323 3882 -26263
rect 4280 -26193 4340 -26133
rect 4280 -26323 4340 -26263
rect 4736 -26193 4796 -26133
rect 4736 -26323 4796 -26263
rect 5192 -26193 5252 -26133
rect 5192 -26323 5252 -26263
rect 5650 -26193 5710 -26133
rect 5650 -26323 5710 -26263
rect 6106 -26193 6166 -26133
rect 6106 -26323 6166 -26263
rect 6562 -26193 6622 -26133
rect 6562 -26323 6622 -26263
rect 7020 -26193 7080 -26133
rect 7020 -26323 7080 -26263
rect 7476 -26193 7536 -26133
rect 7476 -26323 7536 -26263
rect 7932 -26193 7992 -26133
rect 7932 -26323 7992 -26263
rect 8406 -26193 8466 -26133
rect 8406 -26323 8466 -26263
rect 8862 -26193 8922 -26133
rect 8862 -26323 8922 -26263
rect 9320 -26193 9380 -26133
rect 9320 -26323 9380 -26263
rect 9776 -26193 9836 -26133
rect 9776 -26323 9836 -26263
rect 10232 -26193 10292 -26133
rect 10232 -26323 10292 -26263
rect 10690 -26193 10750 -26133
rect 10690 -26323 10750 -26263
rect 11146 -26193 11206 -26133
rect 11146 -26323 11206 -26263
rect 11602 -26193 11662 -26133
rect 11602 -26323 11662 -26263
rect 12060 -26193 12120 -26133
rect 12060 -26323 12120 -26263
rect 12516 -26193 12576 -26133
rect 12516 -26323 12576 -26263
rect 12972 -26193 13032 -26133
rect 12972 -26323 13032 -26263
rect 13430 -26193 13490 -26133
rect 13430 -26323 13490 -26263
rect 13886 -26193 13946 -26133
rect 13886 -26323 13946 -26263
rect 14342 -26193 14402 -26133
rect 14342 -26323 14402 -26263
rect 14800 -26193 14860 -26133
rect 14800 -26323 14860 -26263
rect 15256 -26193 15316 -26133
rect 15256 -26323 15316 -26263
rect 170 -26685 230 -26625
rect 170 -26815 230 -26755
rect 626 -26685 686 -26625
rect 626 -26815 686 -26755
rect 1082 -26685 1142 -26625
rect 1082 -26815 1142 -26755
rect 1540 -26685 1600 -26625
rect 1540 -26815 1600 -26755
rect 1996 -26685 2056 -26625
rect 1996 -26815 2056 -26755
rect 2452 -26685 2512 -26625
rect 2452 -26815 2512 -26755
rect 2910 -26685 2970 -26625
rect 2910 -26815 2970 -26755
rect 3366 -26685 3426 -26625
rect 3366 -26815 3426 -26755
rect 3822 -26685 3882 -26625
rect 3822 -26815 3882 -26755
rect 4280 -26685 4340 -26625
rect 4280 -26815 4340 -26755
rect 4736 -26685 4796 -26625
rect 4736 -26815 4796 -26755
rect 5192 -26685 5252 -26625
rect 5192 -26815 5252 -26755
rect 5650 -26685 5710 -26625
rect 5650 -26815 5710 -26755
rect 6106 -26685 6166 -26625
rect 6106 -26815 6166 -26755
rect 6562 -26685 6622 -26625
rect 6562 -26815 6622 -26755
rect 7020 -26685 7080 -26625
rect 7020 -26815 7080 -26755
rect 7476 -26685 7536 -26625
rect 7476 -26815 7536 -26755
rect 7932 -26685 7992 -26625
rect 7932 -26815 7992 -26755
rect 8406 -26685 8466 -26625
rect 8406 -26815 8466 -26755
rect 8862 -26685 8922 -26625
rect 8862 -26815 8922 -26755
rect 9320 -26685 9380 -26625
rect 9320 -26815 9380 -26755
rect 9776 -26685 9836 -26625
rect 9776 -26815 9836 -26755
rect 10232 -26685 10292 -26625
rect 10232 -26815 10292 -26755
rect 10690 -26685 10750 -26625
rect 10690 -26815 10750 -26755
rect 11146 -26685 11206 -26625
rect 11146 -26815 11206 -26755
rect 11602 -26685 11662 -26625
rect 11602 -26815 11662 -26755
rect 12060 -26685 12120 -26625
rect 12060 -26815 12120 -26755
rect 12516 -26685 12576 -26625
rect 12516 -26815 12576 -26755
rect 12972 -26685 13032 -26625
rect 12972 -26815 13032 -26755
rect 13430 -26685 13490 -26625
rect 13430 -26815 13490 -26755
rect 13886 -26685 13946 -26625
rect 13886 -26815 13946 -26755
rect 14342 -26685 14402 -26625
rect 14342 -26815 14402 -26755
rect 14800 -26685 14860 -26625
rect 14800 -26815 14860 -26755
rect 15256 -26685 15316 -26625
rect 15256 -26815 15316 -26755
rect 170 -27187 230 -27127
rect 170 -27317 230 -27257
rect 626 -27187 686 -27127
rect 626 -27317 686 -27257
rect 1082 -27187 1142 -27127
rect 1082 -27317 1142 -27257
rect 1540 -27187 1600 -27127
rect 1540 -27317 1600 -27257
rect 1996 -27187 2056 -27127
rect 1996 -27317 2056 -27257
rect 2452 -27187 2512 -27127
rect 2452 -27317 2512 -27257
rect 2910 -27187 2970 -27127
rect 2910 -27317 2970 -27257
rect 3366 -27187 3426 -27127
rect 3366 -27317 3426 -27257
rect 3822 -27187 3882 -27127
rect 3822 -27317 3882 -27257
rect 4280 -27187 4340 -27127
rect 4280 -27317 4340 -27257
rect 4736 -27187 4796 -27127
rect 4736 -27317 4796 -27257
rect 5192 -27187 5252 -27127
rect 5192 -27317 5252 -27257
rect 5650 -27187 5710 -27127
rect 5650 -27317 5710 -27257
rect 6106 -27187 6166 -27127
rect 6106 -27317 6166 -27257
rect 6562 -27187 6622 -27127
rect 6562 -27317 6622 -27257
rect 7020 -27187 7080 -27127
rect 7020 -27317 7080 -27257
rect 7476 -27187 7536 -27127
rect 7476 -27317 7536 -27257
rect 7932 -27187 7992 -27127
rect 7932 -27317 7992 -27257
rect 8406 -27187 8466 -27127
rect 8406 -27317 8466 -27257
rect 8862 -27187 8922 -27127
rect 8862 -27317 8922 -27257
rect 9320 -27187 9380 -27127
rect 9320 -27317 9380 -27257
rect 9776 -27187 9836 -27127
rect 9776 -27317 9836 -27257
rect 10232 -27187 10292 -27127
rect 10232 -27317 10292 -27257
rect 10690 -27187 10750 -27127
rect 10690 -27317 10750 -27257
rect 11146 -27187 11206 -27127
rect 11146 -27317 11206 -27257
rect 11602 -27187 11662 -27127
rect 11602 -27317 11662 -27257
rect 12060 -27187 12120 -27127
rect 12060 -27317 12120 -27257
rect 12516 -27187 12576 -27127
rect 12516 -27317 12576 -27257
rect 12972 -27187 13032 -27127
rect 12972 -27317 13032 -27257
rect 13430 -27187 13490 -27127
rect 13430 -27317 13490 -27257
rect 13886 -27187 13946 -27127
rect 13886 -27317 13946 -27257
rect 14342 -27187 14402 -27127
rect 14342 -27317 14402 -27257
rect 14800 -27187 14860 -27127
rect 14800 -27317 14860 -27257
rect 15256 -27187 15316 -27127
rect 15256 -27317 15316 -27257
rect 170 -27703 230 -27643
rect 170 -27833 230 -27773
rect 626 -27703 686 -27643
rect 626 -27833 686 -27773
rect 1082 -27703 1142 -27643
rect 1082 -27833 1142 -27773
rect 1540 -27703 1600 -27643
rect 1540 -27833 1600 -27773
rect 1996 -27703 2056 -27643
rect 1996 -27833 2056 -27773
rect 2452 -27703 2512 -27643
rect 2452 -27833 2512 -27773
rect 2910 -27703 2970 -27643
rect 2910 -27833 2970 -27773
rect 3366 -27703 3426 -27643
rect 3366 -27833 3426 -27773
rect 3822 -27703 3882 -27643
rect 3822 -27833 3882 -27773
rect 4280 -27703 4340 -27643
rect 4280 -27833 4340 -27773
rect 4736 -27703 4796 -27643
rect 4736 -27833 4796 -27773
rect 5192 -27703 5252 -27643
rect 5192 -27833 5252 -27773
rect 5650 -27703 5710 -27643
rect 5650 -27833 5710 -27773
rect 6106 -27703 6166 -27643
rect 6106 -27833 6166 -27773
rect 6562 -27703 6622 -27643
rect 6562 -27833 6622 -27773
rect 7020 -27703 7080 -27643
rect 7020 -27833 7080 -27773
rect 7476 -27703 7536 -27643
rect 7476 -27833 7536 -27773
rect 7932 -27703 7992 -27643
rect 7932 -27833 7992 -27773
rect 8406 -27703 8466 -27643
rect 8406 -27833 8466 -27773
rect 8862 -27703 8922 -27643
rect 8862 -27833 8922 -27773
rect 9320 -27703 9380 -27643
rect 9320 -27833 9380 -27773
rect 9776 -27703 9836 -27643
rect 9776 -27833 9836 -27773
rect 10232 -27703 10292 -27643
rect 10232 -27833 10292 -27773
rect 10690 -27703 10750 -27643
rect 10690 -27833 10750 -27773
rect 11146 -27703 11206 -27643
rect 11146 -27833 11206 -27773
rect 11602 -27703 11662 -27643
rect 11602 -27833 11662 -27773
rect 12060 -27703 12120 -27643
rect 12060 -27833 12120 -27773
rect 12516 -27703 12576 -27643
rect 12516 -27833 12576 -27773
rect 12972 -27703 13032 -27643
rect 12972 -27833 13032 -27773
rect 13430 -27703 13490 -27643
rect 13430 -27833 13490 -27773
rect 13886 -27703 13946 -27643
rect 13886 -27833 13946 -27773
rect 14342 -27703 14402 -27643
rect 14342 -27833 14402 -27773
rect 14800 -27703 14860 -27643
rect 14800 -27833 14860 -27773
rect 15256 -27703 15316 -27643
rect 15256 -27833 15316 -27773
rect 170 -28195 230 -28135
rect 170 -28325 230 -28265
rect 626 -28195 686 -28135
rect 626 -28325 686 -28265
rect 1082 -28195 1142 -28135
rect 1082 -28325 1142 -28265
rect 1540 -28195 1600 -28135
rect 1540 -28325 1600 -28265
rect 1996 -28195 2056 -28135
rect 1996 -28325 2056 -28265
rect 2452 -28195 2512 -28135
rect 2452 -28325 2512 -28265
rect 2910 -28195 2970 -28135
rect 2910 -28325 2970 -28265
rect 3366 -28195 3426 -28135
rect 3366 -28325 3426 -28265
rect 3822 -28195 3882 -28135
rect 3822 -28325 3882 -28265
rect 4280 -28195 4340 -28135
rect 4280 -28325 4340 -28265
rect 4736 -28195 4796 -28135
rect 4736 -28325 4796 -28265
rect 5192 -28195 5252 -28135
rect 5192 -28325 5252 -28265
rect 5650 -28195 5710 -28135
rect 5650 -28325 5710 -28265
rect 6106 -28195 6166 -28135
rect 6106 -28325 6166 -28265
rect 6562 -28195 6622 -28135
rect 6562 -28325 6622 -28265
rect 7020 -28195 7080 -28135
rect 7020 -28325 7080 -28265
rect 7476 -28195 7536 -28135
rect 7476 -28325 7536 -28265
rect 7932 -28195 7992 -28135
rect 7932 -28325 7992 -28265
rect 8406 -28195 8466 -28135
rect 8406 -28325 8466 -28265
rect 8862 -28195 8922 -28135
rect 8862 -28325 8922 -28265
rect 9320 -28195 9380 -28135
rect 9320 -28325 9380 -28265
rect 9776 -28195 9836 -28135
rect 9776 -28325 9836 -28265
rect 10232 -28195 10292 -28135
rect 10232 -28325 10292 -28265
rect 10690 -28195 10750 -28135
rect 10690 -28325 10750 -28265
rect 11146 -28195 11206 -28135
rect 11146 -28325 11206 -28265
rect 11602 -28195 11662 -28135
rect 11602 -28325 11662 -28265
rect 12060 -28195 12120 -28135
rect 12060 -28325 12120 -28265
rect 12516 -28195 12576 -28135
rect 12516 -28325 12576 -28265
rect 12972 -28195 13032 -28135
rect 12972 -28325 13032 -28265
rect 13430 -28195 13490 -28135
rect 13430 -28325 13490 -28265
rect 13886 -28195 13946 -28135
rect 13886 -28325 13946 -28265
rect 14342 -28195 14402 -28135
rect 14342 -28325 14402 -28265
rect 14800 -28195 14860 -28135
rect 14800 -28325 14860 -28265
rect 15256 -28195 15316 -28135
rect 15256 -28325 15316 -28265
rect 170 -28697 230 -28637
rect 170 -28827 230 -28767
rect 626 -28697 686 -28637
rect 626 -28827 686 -28767
rect 1082 -28697 1142 -28637
rect 1082 -28827 1142 -28767
rect 1540 -28697 1600 -28637
rect 1540 -28827 1600 -28767
rect 1996 -28697 2056 -28637
rect 1996 -28827 2056 -28767
rect 2452 -28697 2512 -28637
rect 2452 -28827 2512 -28767
rect 2910 -28697 2970 -28637
rect 2910 -28827 2970 -28767
rect 3366 -28697 3426 -28637
rect 3366 -28827 3426 -28767
rect 3822 -28697 3882 -28637
rect 3822 -28827 3882 -28767
rect 4280 -28697 4340 -28637
rect 4280 -28827 4340 -28767
rect 4736 -28697 4796 -28637
rect 4736 -28827 4796 -28767
rect 5192 -28697 5252 -28637
rect 5192 -28827 5252 -28767
rect 5650 -28697 5710 -28637
rect 5650 -28827 5710 -28767
rect 6106 -28697 6166 -28637
rect 6106 -28827 6166 -28767
rect 6562 -28697 6622 -28637
rect 6562 -28827 6622 -28767
rect 7020 -28697 7080 -28637
rect 7020 -28827 7080 -28767
rect 7476 -28697 7536 -28637
rect 7476 -28827 7536 -28767
rect 7932 -28697 7992 -28637
rect 7932 -28827 7992 -28767
rect 8406 -28697 8466 -28637
rect 8406 -28827 8466 -28767
rect 8862 -28697 8922 -28637
rect 8862 -28827 8922 -28767
rect 9320 -28697 9380 -28637
rect 9320 -28827 9380 -28767
rect 9776 -28697 9836 -28637
rect 9776 -28827 9836 -28767
rect 10232 -28697 10292 -28637
rect 10232 -28827 10292 -28767
rect 10690 -28697 10750 -28637
rect 10690 -28827 10750 -28767
rect 11146 -28697 11206 -28637
rect 11146 -28827 11206 -28767
rect 11602 -28697 11662 -28637
rect 11602 -28827 11662 -28767
rect 12060 -28697 12120 -28637
rect 12060 -28827 12120 -28767
rect 12516 -28697 12576 -28637
rect 12516 -28827 12576 -28767
rect 12972 -28697 13032 -28637
rect 12972 -28827 13032 -28767
rect 13430 -28697 13490 -28637
rect 13430 -28827 13490 -28767
rect 13886 -28697 13946 -28637
rect 13886 -28827 13946 -28767
rect 14342 -28697 14402 -28637
rect 14342 -28827 14402 -28767
rect 14800 -28697 14860 -28637
rect 14800 -28827 14860 -28767
rect 15256 -28697 15316 -28637
rect 15256 -28827 15316 -28767
rect 170 -29191 230 -29131
rect 170 -29321 230 -29261
rect 626 -29191 686 -29131
rect 626 -29321 686 -29261
rect 1082 -29191 1142 -29131
rect 1082 -29321 1142 -29261
rect 1540 -29191 1600 -29131
rect 1540 -29321 1600 -29261
rect 1996 -29191 2056 -29131
rect 1996 -29321 2056 -29261
rect 2452 -29191 2512 -29131
rect 2452 -29321 2512 -29261
rect 2910 -29191 2970 -29131
rect 2910 -29321 2970 -29261
rect 3366 -29191 3426 -29131
rect 3366 -29321 3426 -29261
rect 3822 -29191 3882 -29131
rect 3822 -29321 3882 -29261
rect 4280 -29191 4340 -29131
rect 4280 -29321 4340 -29261
rect 4736 -29191 4796 -29131
rect 4736 -29321 4796 -29261
rect 5192 -29191 5252 -29131
rect 5192 -29321 5252 -29261
rect 5650 -29191 5710 -29131
rect 5650 -29321 5710 -29261
rect 6106 -29191 6166 -29131
rect 6106 -29321 6166 -29261
rect 6562 -29191 6622 -29131
rect 6562 -29321 6622 -29261
rect 7020 -29191 7080 -29131
rect 7020 -29321 7080 -29261
rect 7476 -29191 7536 -29131
rect 7476 -29321 7536 -29261
rect 7932 -29191 7992 -29131
rect 7932 -29321 7992 -29261
rect 8406 -29191 8466 -29131
rect 8406 -29321 8466 -29261
rect 8862 -29191 8922 -29131
rect 8862 -29321 8922 -29261
rect 9320 -29191 9380 -29131
rect 9320 -29321 9380 -29261
rect 9776 -29191 9836 -29131
rect 9776 -29321 9836 -29261
rect 10232 -29191 10292 -29131
rect 10232 -29321 10292 -29261
rect 10690 -29191 10750 -29131
rect 10690 -29321 10750 -29261
rect 11146 -29191 11206 -29131
rect 11146 -29321 11206 -29261
rect 11602 -29191 11662 -29131
rect 11602 -29321 11662 -29261
rect 12060 -29191 12120 -29131
rect 12060 -29321 12120 -29261
rect 12516 -29191 12576 -29131
rect 12516 -29321 12576 -29261
rect 12972 -29191 13032 -29131
rect 12972 -29321 13032 -29261
rect 13430 -29191 13490 -29131
rect 13430 -29321 13490 -29261
rect 13886 -29191 13946 -29131
rect 13886 -29321 13946 -29261
rect 14342 -29191 14402 -29131
rect 14342 -29321 14402 -29261
rect 14800 -29191 14860 -29131
rect 14800 -29321 14860 -29261
rect 15256 -29191 15316 -29131
rect 15256 -29321 15316 -29261
rect 170 -29683 230 -29623
rect 170 -29813 230 -29753
rect 626 -29683 686 -29623
rect 626 -29813 686 -29753
rect 1082 -29683 1142 -29623
rect 1082 -29813 1142 -29753
rect 1540 -29683 1600 -29623
rect 1540 -29813 1600 -29753
rect 1996 -29683 2056 -29623
rect 1996 -29813 2056 -29753
rect 2452 -29683 2512 -29623
rect 2452 -29813 2512 -29753
rect 2910 -29683 2970 -29623
rect 2910 -29813 2970 -29753
rect 3366 -29683 3426 -29623
rect 3366 -29813 3426 -29753
rect 3822 -29683 3882 -29623
rect 3822 -29813 3882 -29753
rect 4280 -29683 4340 -29623
rect 4280 -29813 4340 -29753
rect 4736 -29683 4796 -29623
rect 4736 -29813 4796 -29753
rect 5192 -29683 5252 -29623
rect 5192 -29813 5252 -29753
rect 5650 -29683 5710 -29623
rect 5650 -29813 5710 -29753
rect 6106 -29683 6166 -29623
rect 6106 -29813 6166 -29753
rect 6562 -29683 6622 -29623
rect 6562 -29813 6622 -29753
rect 7020 -29683 7080 -29623
rect 7020 -29813 7080 -29753
rect 7476 -29683 7536 -29623
rect 7476 -29813 7536 -29753
rect 7932 -29683 7992 -29623
rect 7932 -29813 7992 -29753
rect 8406 -29683 8466 -29623
rect 8406 -29813 8466 -29753
rect 8862 -29683 8922 -29623
rect 8862 -29813 8922 -29753
rect 9320 -29683 9380 -29623
rect 9320 -29813 9380 -29753
rect 9776 -29683 9836 -29623
rect 9776 -29813 9836 -29753
rect 10232 -29683 10292 -29623
rect 10232 -29813 10292 -29753
rect 10690 -29683 10750 -29623
rect 10690 -29813 10750 -29753
rect 11146 -29683 11206 -29623
rect 11146 -29813 11206 -29753
rect 11602 -29683 11662 -29623
rect 11602 -29813 11662 -29753
rect 12060 -29683 12120 -29623
rect 12060 -29813 12120 -29753
rect 12516 -29683 12576 -29623
rect 12516 -29813 12576 -29753
rect 12972 -29683 13032 -29623
rect 12972 -29813 13032 -29753
rect 13430 -29683 13490 -29623
rect 13430 -29813 13490 -29753
rect 13886 -29683 13946 -29623
rect 13886 -29813 13946 -29753
rect 14342 -29683 14402 -29623
rect 14342 -29813 14402 -29753
rect 14800 -29683 14860 -29623
rect 14800 -29813 14860 -29753
rect 15256 -29683 15316 -29623
rect 15256 -29813 15316 -29753
rect 170 -30185 230 -30125
rect 170 -30315 230 -30255
rect 626 -30185 686 -30125
rect 626 -30315 686 -30255
rect 1082 -30185 1142 -30125
rect 1082 -30315 1142 -30255
rect 1540 -30185 1600 -30125
rect 1540 -30315 1600 -30255
rect 1996 -30185 2056 -30125
rect 1996 -30315 2056 -30255
rect 2452 -30185 2512 -30125
rect 2452 -30315 2512 -30255
rect 2910 -30185 2970 -30125
rect 2910 -30315 2970 -30255
rect 3366 -30185 3426 -30125
rect 3366 -30315 3426 -30255
rect 3822 -30185 3882 -30125
rect 3822 -30315 3882 -30255
rect 4280 -30185 4340 -30125
rect 4280 -30315 4340 -30255
rect 4736 -30185 4796 -30125
rect 4736 -30315 4796 -30255
rect 5192 -30185 5252 -30125
rect 5192 -30315 5252 -30255
rect 5650 -30185 5710 -30125
rect 5650 -30315 5710 -30255
rect 6106 -30185 6166 -30125
rect 6106 -30315 6166 -30255
rect 6562 -30185 6622 -30125
rect 6562 -30315 6622 -30255
rect 7020 -30185 7080 -30125
rect 7020 -30315 7080 -30255
rect 7476 -30185 7536 -30125
rect 7476 -30315 7536 -30255
rect 7932 -30185 7992 -30125
rect 7932 -30315 7992 -30255
rect 8406 -30185 8466 -30125
rect 8406 -30315 8466 -30255
rect 8862 -30185 8922 -30125
rect 8862 -30315 8922 -30255
rect 9320 -30185 9380 -30125
rect 9320 -30315 9380 -30255
rect 9776 -30185 9836 -30125
rect 9776 -30315 9836 -30255
rect 10232 -30185 10292 -30125
rect 10232 -30315 10292 -30255
rect 10690 -30185 10750 -30125
rect 10690 -30315 10750 -30255
rect 11146 -30185 11206 -30125
rect 11146 -30315 11206 -30255
rect 11602 -30185 11662 -30125
rect 11602 -30315 11662 -30255
rect 12060 -30185 12120 -30125
rect 12060 -30315 12120 -30255
rect 12516 -30185 12576 -30125
rect 12516 -30315 12576 -30255
rect 12972 -30185 13032 -30125
rect 12972 -30315 13032 -30255
rect 13430 -30185 13490 -30125
rect 13430 -30315 13490 -30255
rect 13886 -30185 13946 -30125
rect 13886 -30315 13946 -30255
rect 14342 -30185 14402 -30125
rect 14342 -30315 14402 -30255
rect 14800 -30185 14860 -30125
rect 14800 -30315 14860 -30255
rect 15256 -30185 15316 -30125
rect 15256 -30315 15316 -30255
rect 170 -30701 230 -30641
rect 170 -30831 230 -30771
rect 626 -30701 686 -30641
rect 626 -30831 686 -30771
rect 1082 -30701 1142 -30641
rect 1082 -30831 1142 -30771
rect 1540 -30701 1600 -30641
rect 1540 -30831 1600 -30771
rect 1996 -30701 2056 -30641
rect 1996 -30831 2056 -30771
rect 2452 -30701 2512 -30641
rect 2452 -30831 2512 -30771
rect 2910 -30701 2970 -30641
rect 2910 -30831 2970 -30771
rect 3366 -30701 3426 -30641
rect 3366 -30831 3426 -30771
rect 3822 -30701 3882 -30641
rect 3822 -30831 3882 -30771
rect 4280 -30701 4340 -30641
rect 4280 -30831 4340 -30771
rect 4736 -30701 4796 -30641
rect 4736 -30831 4796 -30771
rect 5192 -30701 5252 -30641
rect 5192 -30831 5252 -30771
rect 5650 -30701 5710 -30641
rect 5650 -30831 5710 -30771
rect 6106 -30701 6166 -30641
rect 6106 -30831 6166 -30771
rect 6562 -30701 6622 -30641
rect 6562 -30831 6622 -30771
rect 7020 -30701 7080 -30641
rect 7020 -30831 7080 -30771
rect 7476 -30701 7536 -30641
rect 7476 -30831 7536 -30771
rect 7932 -30701 7992 -30641
rect 7932 -30831 7992 -30771
rect 8406 -30701 8466 -30641
rect 8406 -30831 8466 -30771
rect 8862 -30701 8922 -30641
rect 8862 -30831 8922 -30771
rect 9320 -30701 9380 -30641
rect 9320 -30831 9380 -30771
rect 9776 -30701 9836 -30641
rect 9776 -30831 9836 -30771
rect 10232 -30701 10292 -30641
rect 10232 -30831 10292 -30771
rect 10690 -30701 10750 -30641
rect 10690 -30831 10750 -30771
rect 11146 -30701 11206 -30641
rect 11146 -30831 11206 -30771
rect 11602 -30701 11662 -30641
rect 11602 -30831 11662 -30771
rect 12060 -30701 12120 -30641
rect 12060 -30831 12120 -30771
rect 12516 -30701 12576 -30641
rect 12516 -30831 12576 -30771
rect 12972 -30701 13032 -30641
rect 12972 -30831 13032 -30771
rect 13430 -30701 13490 -30641
rect 13430 -30831 13490 -30771
rect 13886 -30701 13946 -30641
rect 13886 -30831 13946 -30771
rect 14342 -30701 14402 -30641
rect 14342 -30831 14402 -30771
rect 14800 -30701 14860 -30641
rect 14800 -30831 14860 -30771
rect 15256 -30701 15316 -30641
rect 15256 -30831 15316 -30771
rect 170 -31193 230 -31133
rect 170 -31323 230 -31263
rect 626 -31193 686 -31133
rect 626 -31323 686 -31263
rect 1082 -31193 1142 -31133
rect 1082 -31323 1142 -31263
rect 1540 -31193 1600 -31133
rect 1540 -31323 1600 -31263
rect 1996 -31193 2056 -31133
rect 1996 -31323 2056 -31263
rect 2452 -31193 2512 -31133
rect 2452 -31323 2512 -31263
rect 2910 -31193 2970 -31133
rect 2910 -31323 2970 -31263
rect 3366 -31193 3426 -31133
rect 3366 -31323 3426 -31263
rect 3822 -31193 3882 -31133
rect 3822 -31323 3882 -31263
rect 4280 -31193 4340 -31133
rect 4280 -31323 4340 -31263
rect 4736 -31193 4796 -31133
rect 4736 -31323 4796 -31263
rect 5192 -31193 5252 -31133
rect 5192 -31323 5252 -31263
rect 5650 -31193 5710 -31133
rect 5650 -31323 5710 -31263
rect 6106 -31193 6166 -31133
rect 6106 -31323 6166 -31263
rect 6562 -31193 6622 -31133
rect 6562 -31323 6622 -31263
rect 7020 -31193 7080 -31133
rect 7020 -31323 7080 -31263
rect 7476 -31193 7536 -31133
rect 7476 -31323 7536 -31263
rect 7932 -31193 7992 -31133
rect 7932 -31323 7992 -31263
rect 8406 -31193 8466 -31133
rect 8406 -31323 8466 -31263
rect 8862 -31193 8922 -31133
rect 8862 -31323 8922 -31263
rect 9320 -31193 9380 -31133
rect 9320 -31323 9380 -31263
rect 9776 -31193 9836 -31133
rect 9776 -31323 9836 -31263
rect 10232 -31193 10292 -31133
rect 10232 -31323 10292 -31263
rect 10690 -31193 10750 -31133
rect 10690 -31323 10750 -31263
rect 11146 -31193 11206 -31133
rect 11146 -31323 11206 -31263
rect 11602 -31193 11662 -31133
rect 11602 -31323 11662 -31263
rect 12060 -31193 12120 -31133
rect 12060 -31323 12120 -31263
rect 12516 -31193 12576 -31133
rect 12516 -31323 12576 -31263
rect 12972 -31193 13032 -31133
rect 12972 -31323 13032 -31263
rect 13430 -31193 13490 -31133
rect 13430 -31323 13490 -31263
rect 13886 -31193 13946 -31133
rect 13886 -31323 13946 -31263
rect 14342 -31193 14402 -31133
rect 14342 -31323 14402 -31263
rect 14800 -31193 14860 -31133
rect 14800 -31323 14860 -31263
rect 15256 -31193 15316 -31133
rect 15256 -31323 15316 -31263
rect 170 -31695 230 -31635
rect 170 -31825 230 -31765
rect 626 -31695 686 -31635
rect 626 -31825 686 -31765
rect 1082 -31695 1142 -31635
rect 1082 -31825 1142 -31765
rect 1540 -31695 1600 -31635
rect 1540 -31825 1600 -31765
rect 1996 -31695 2056 -31635
rect 1996 -31825 2056 -31765
rect 2452 -31695 2512 -31635
rect 2452 -31825 2512 -31765
rect 2910 -31695 2970 -31635
rect 2910 -31825 2970 -31765
rect 3366 -31695 3426 -31635
rect 3366 -31825 3426 -31765
rect 3822 -31695 3882 -31635
rect 3822 -31825 3882 -31765
rect 4280 -31695 4340 -31635
rect 4280 -31825 4340 -31765
rect 4736 -31695 4796 -31635
rect 4736 -31825 4796 -31765
rect 5192 -31695 5252 -31635
rect 5192 -31825 5252 -31765
rect 5650 -31695 5710 -31635
rect 5650 -31825 5710 -31765
rect 6106 -31695 6166 -31635
rect 6106 -31825 6166 -31765
rect 6562 -31695 6622 -31635
rect 6562 -31825 6622 -31765
rect 7020 -31695 7080 -31635
rect 7020 -31825 7080 -31765
rect 7476 -31695 7536 -31635
rect 7476 -31825 7536 -31765
rect 7932 -31695 7992 -31635
rect 7932 -31825 7992 -31765
rect 8406 -31695 8466 -31635
rect 8406 -31825 8466 -31765
rect 8862 -31695 8922 -31635
rect 8862 -31825 8922 -31765
rect 9320 -31695 9380 -31635
rect 9320 -31825 9380 -31765
rect 9776 -31695 9836 -31635
rect 9776 -31825 9836 -31765
rect 10232 -31695 10292 -31635
rect 10232 -31825 10292 -31765
rect 10690 -31695 10750 -31635
rect 10690 -31825 10750 -31765
rect 11146 -31695 11206 -31635
rect 11146 -31825 11206 -31765
rect 11602 -31695 11662 -31635
rect 11602 -31825 11662 -31765
rect 12060 -31695 12120 -31635
rect 12060 -31825 12120 -31765
rect 12516 -31695 12576 -31635
rect 12516 -31825 12576 -31765
rect 12972 -31695 13032 -31635
rect 12972 -31825 13032 -31765
rect 13430 -31695 13490 -31635
rect 13430 -31825 13490 -31765
rect 13886 -31695 13946 -31635
rect 13886 -31825 13946 -31765
rect 14342 -31695 14402 -31635
rect 14342 -31825 14402 -31765
rect 14800 -31695 14860 -31635
rect 14800 -31825 14860 -31765
rect 15256 -31695 15316 -31635
rect 15256 -31825 15316 -31765
rect 170 -32187 230 -32127
rect 170 -32317 230 -32257
rect 626 -32187 686 -32127
rect 626 -32317 686 -32257
rect 1082 -32187 1142 -32127
rect 1082 -32317 1142 -32257
rect 1540 -32187 1600 -32127
rect 1540 -32317 1600 -32257
rect 1996 -32187 2056 -32127
rect 1996 -32317 2056 -32257
rect 2452 -32187 2512 -32127
rect 2452 -32317 2512 -32257
rect 2910 -32187 2970 -32127
rect 2910 -32317 2970 -32257
rect 3366 -32187 3426 -32127
rect 3366 -32317 3426 -32257
rect 3822 -32187 3882 -32127
rect 3822 -32317 3882 -32257
rect 4280 -32187 4340 -32127
rect 4280 -32317 4340 -32257
rect 4736 -32187 4796 -32127
rect 4736 -32317 4796 -32257
rect 5192 -32187 5252 -32127
rect 5192 -32317 5252 -32257
rect 5650 -32187 5710 -32127
rect 5650 -32317 5710 -32257
rect 6106 -32187 6166 -32127
rect 6106 -32317 6166 -32257
rect 6562 -32187 6622 -32127
rect 6562 -32317 6622 -32257
rect 7020 -32187 7080 -32127
rect 7020 -32317 7080 -32257
rect 7476 -32187 7536 -32127
rect 7476 -32317 7536 -32257
rect 7932 -32187 7992 -32127
rect 7932 -32317 7992 -32257
rect 8406 -32187 8466 -32127
rect 8406 -32317 8466 -32257
rect 8862 -32187 8922 -32127
rect 8862 -32317 8922 -32257
rect 9320 -32187 9380 -32127
rect 9320 -32317 9380 -32257
rect 9776 -32187 9836 -32127
rect 9776 -32317 9836 -32257
rect 10232 -32187 10292 -32127
rect 10232 -32317 10292 -32257
rect 10690 -32187 10750 -32127
rect 10690 -32317 10750 -32257
rect 11146 -32187 11206 -32127
rect 11146 -32317 11206 -32257
rect 11602 -32187 11662 -32127
rect 11602 -32317 11662 -32257
rect 12060 -32187 12120 -32127
rect 12060 -32317 12120 -32257
rect 12516 -32187 12576 -32127
rect 12516 -32317 12576 -32257
rect 12972 -32187 13032 -32127
rect 12972 -32317 13032 -32257
rect 13430 -32187 13490 -32127
rect 13430 -32317 13490 -32257
rect 13886 -32187 13946 -32127
rect 13886 -32317 13946 -32257
rect 14342 -32187 14402 -32127
rect 14342 -32317 14402 -32257
rect 14800 -32187 14860 -32127
rect 14800 -32317 14860 -32257
rect 15256 -32187 15316 -32127
rect 15256 -32317 15316 -32257
<< metal4 >>
rect 78 651 321 661
rect 78 590 89 651
rect 150 590 250 651
rect 311 590 321 651
rect 15111 622 15452 623
rect 78 580 321 590
rect 170 330 230 580
rect 15110 551 15127 622
rect 15200 621 15452 622
rect 15200 612 15357 621
rect 15201 551 15357 612
rect 15430 611 15452 621
rect 15432 551 15452 611
rect 15110 550 15357 551
rect 15430 550 15452 551
rect 15110 539 15452 550
rect 1540 364 1600 460
rect 1996 364 2056 460
rect 2452 364 2512 460
rect 2910 364 2970 460
rect 3366 364 3426 460
rect 3822 364 3882 460
rect 4280 364 4340 460
rect 4736 364 4796 460
rect 5192 364 5252 460
rect 5650 364 5710 460
rect 6106 364 6166 460
rect 6562 364 6622 460
rect 7020 364 7080 460
rect 7476 364 7536 460
rect 7932 364 7992 460
rect 8406 364 8466 451
rect 8862 364 8922 451
rect 9320 364 9380 451
rect 9776 364 9836 451
rect 10232 364 10292 451
rect 10690 364 10750 451
rect 11146 364 11206 451
rect 11602 364 11662 451
rect 12060 364 12120 451
rect 12516 364 12576 451
rect 12972 364 13032 451
rect 13430 364 13490 451
rect 13886 364 13946 451
rect 14342 364 14402 451
rect 14800 365 14860 451
rect 580 348 731 360
rect 580 270 614 348
rect 699 270 731 348
rect 580 140 731 270
rect 1035 350 1177 363
rect 1035 271 1066 350
rect 1154 271 1177 350
rect 1035 139 1177 271
rect 1498 350 1640 364
rect 1498 270 1527 350
rect 1612 270 1640 350
rect 1498 200 1640 270
rect 1498 140 1540 200
rect 1600 140 1640 200
rect 1956 350 2098 364
rect 1956 270 1982 350
rect 2067 270 2098 350
rect 1956 200 2098 270
rect 1956 140 1996 200
rect 2056 140 2098 200
rect 2414 350 2556 364
rect 2414 270 2438 350
rect 2523 270 2556 350
rect 2414 200 2556 270
rect 2414 140 2452 200
rect 2512 140 2556 200
rect 2869 350 3011 364
rect 2869 270 2897 350
rect 2982 270 3011 350
rect 2869 200 3011 270
rect 2869 140 2910 200
rect 2970 140 3011 200
rect 3324 350 3466 364
rect 3324 270 3355 350
rect 3440 270 3466 350
rect 3324 200 3466 270
rect 3324 140 3366 200
rect 3426 140 3466 200
rect 3779 350 3921 364
rect 3779 270 3807 350
rect 3892 270 3921 350
rect 3779 200 3921 270
rect 3779 140 3822 200
rect 3882 140 3921 200
rect 4235 350 4377 364
rect 4235 270 4267 350
rect 4352 270 4377 350
rect 4235 200 4377 270
rect 4235 140 4280 200
rect 4340 140 4377 200
rect 4695 350 4837 364
rect 4695 270 4721 350
rect 4806 270 4837 350
rect 4695 200 4837 270
rect 4695 140 4736 200
rect 4796 140 4837 200
rect 5150 350 5292 364
rect 5150 270 5180 350
rect 5265 270 5292 350
rect 5150 200 5292 270
rect 5150 140 5192 200
rect 5252 140 5292 200
rect 5609 350 5751 364
rect 5609 270 5636 350
rect 5721 270 5751 350
rect 5609 200 5751 270
rect 5609 140 5650 200
rect 5710 140 5751 200
rect 6065 350 6207 364
rect 6065 270 6094 350
rect 6179 270 6207 350
rect 6065 200 6207 270
rect 6065 140 6106 200
rect 6166 140 6207 200
rect 6519 350 6661 364
rect 6519 270 6548 350
rect 6633 270 6661 350
rect 6519 200 6661 270
rect 6519 140 6562 200
rect 6622 140 6661 200
rect 6978 350 7120 364
rect 6978 270 7008 350
rect 7093 270 7120 350
rect 6978 200 7120 270
rect 6978 140 7020 200
rect 7080 140 7120 200
rect 7435 350 7577 364
rect 7435 270 7464 350
rect 7549 270 7577 350
rect 7435 200 7577 270
rect 7435 140 7476 200
rect 7536 140 7577 200
rect 7889 350 8031 364
rect 7889 270 7917 350
rect 8002 270 8031 350
rect 7889 200 8031 270
rect 7889 140 7932 200
rect 7992 140 8031 200
rect 8364 350 8506 364
rect 8364 270 8394 350
rect 8479 270 8506 350
rect 8364 200 8506 270
rect 8364 140 8406 200
rect 8466 140 8506 200
rect 8821 350 8963 364
rect 8821 270 8848 350
rect 8933 270 8963 350
rect 8821 200 8963 270
rect 8821 140 8862 200
rect 8922 140 8963 200
rect 9278 350 9420 364
rect 9278 270 9306 350
rect 9391 270 9420 350
rect 9278 200 9420 270
rect 9278 140 9320 200
rect 9380 140 9420 200
rect 9733 350 9875 364
rect 9733 270 9763 350
rect 9848 270 9875 350
rect 9733 200 9875 270
rect 9733 140 9776 200
rect 9836 140 9875 200
rect 10189 350 10331 364
rect 10189 270 10219 350
rect 10304 270 10331 350
rect 10189 200 10331 270
rect 10189 140 10232 200
rect 10292 140 10331 200
rect 10650 350 10792 364
rect 10650 270 10678 350
rect 10763 270 10792 350
rect 10650 200 10792 270
rect 10650 140 10690 200
rect 10750 140 10792 200
rect 11104 350 11246 364
rect 11104 270 11134 350
rect 11219 270 11246 350
rect 11104 200 11246 270
rect 11104 140 11146 200
rect 11206 140 11246 200
rect 11560 350 11702 364
rect 11560 270 11588 350
rect 11673 270 11702 350
rect 11560 200 11702 270
rect 11560 140 11602 200
rect 11662 140 11702 200
rect 12018 350 12160 364
rect 12018 270 12048 350
rect 12133 270 12160 350
rect 12018 200 12160 270
rect 12018 140 12060 200
rect 12120 140 12160 200
rect 12474 350 12616 364
rect 12474 270 12505 350
rect 12590 270 12616 350
rect 12474 200 12616 270
rect 12474 140 12516 200
rect 12576 140 12616 200
rect 12929 350 13071 364
rect 12929 270 12959 350
rect 13044 270 13071 350
rect 12929 200 13071 270
rect 12929 140 12972 200
rect 13032 140 13071 200
rect 13390 350 13532 364
rect 13390 270 13419 350
rect 13504 270 13532 350
rect 13390 200 13532 270
rect 13390 140 13430 200
rect 13490 140 13532 200
rect 13845 350 13987 364
rect 13845 270 13872 350
rect 13957 270 13987 350
rect 13845 200 13987 270
rect 13845 140 13886 200
rect 13946 140 13987 200
rect 14301 350 14443 364
rect 14301 270 14330 350
rect 14415 270 14443 350
rect 14301 200 14443 270
rect 14301 140 14342 200
rect 14402 140 14443 200
rect 14757 350 14899 365
rect 14757 270 14790 350
rect 14875 270 14899 350
rect 15237 343 15330 539
rect 14757 200 14899 270
rect 14757 141 14800 200
rect 14790 140 14800 141
rect 14860 141 14899 200
rect 15209 330 15371 343
rect 15209 270 15256 330
rect 15316 270 15371 330
rect 15209 200 15371 270
rect 14860 140 14870 141
rect 15209 140 15256 200
rect 15316 140 15371 200
rect 1540 8 1600 140
rect 1996 8 2056 140
rect 2452 8 2512 140
rect 2910 8 2970 140
rect 3366 8 3426 140
rect 3822 8 3882 140
rect 4280 8 4340 140
rect 4736 8 4796 140
rect 5192 8 5252 140
rect 5650 8 5710 140
rect 6106 8 6166 140
rect 6562 8 6622 140
rect 170 -162 230 8
rect 1599 6 1600 8
rect 2055 6 2056 8
rect 2511 7 2512 8
rect 160 -222 170 -172
rect 626 -162 686 5
rect 230 -222 240 -172
rect 160 -292 240 -222
rect 160 -352 170 -292
rect 230 -352 240 -292
rect 616 -222 626 -172
rect 1082 -162 1142 6
rect 686 -222 696 -172
rect 616 -292 696 -222
rect 616 -352 626 -292
rect 686 -352 696 -292
rect 1072 -222 1082 -172
rect 1540 -162 1600 6
rect 1142 -222 1152 -172
rect 1072 -292 1152 -222
rect 1072 -352 1082 -292
rect 1142 -352 1152 -292
rect 1530 -222 1540 -172
rect 1996 -162 2056 6
rect 1600 -222 1610 -172
rect 1530 -292 1610 -222
rect 1530 -352 1540 -292
rect 1600 -352 1610 -292
rect 1986 -222 1996 -172
rect 2452 -162 2512 7
rect 2969 6 2970 8
rect 3425 7 3426 8
rect 2056 -222 2066 -172
rect 1986 -292 2066 -222
rect 1986 -352 1996 -292
rect 2056 -352 2066 -292
rect 2442 -222 2452 -172
rect 2910 -162 2970 6
rect 2512 -222 2522 -172
rect 2442 -292 2522 -222
rect 2442 -352 2452 -292
rect 2512 -352 2522 -292
rect 2900 -222 2910 -172
rect 3366 -162 3426 7
rect 3881 6 3882 8
rect 4339 6 4340 8
rect 4795 7 4796 8
rect 2970 -222 2980 -172
rect 2900 -292 2980 -222
rect 2900 -352 2910 -292
rect 2970 -352 2980 -292
rect 3356 -222 3366 -172
rect 3822 -162 3882 6
rect 3426 -222 3436 -172
rect 3356 -292 3436 -222
rect 3356 -352 3366 -292
rect 3426 -352 3436 -292
rect 3812 -222 3822 -172
rect 4280 -162 4340 6
rect 3882 -222 3892 -172
rect 3812 -292 3892 -222
rect 3812 -352 3822 -292
rect 3882 -352 3892 -292
rect 4270 -222 4280 -172
rect 4736 -162 4796 7
rect 5251 6 5252 8
rect 5709 7 5710 8
rect 4340 -222 4350 -172
rect 4270 -292 4350 -222
rect 4270 -352 4280 -292
rect 4340 -352 4350 -292
rect 4726 -222 4736 -172
rect 5192 -162 5252 6
rect 4796 -222 4806 -172
rect 4726 -292 4806 -222
rect 4726 -352 4736 -292
rect 4796 -352 4806 -292
rect 5182 -222 5192 -172
rect 5650 -162 5710 7
rect 6165 6 6166 8
rect 6621 7 6622 8
rect 5252 -222 5262 -172
rect 5182 -292 5262 -222
rect 5182 -352 5192 -292
rect 5252 -352 5262 -292
rect 5640 -222 5650 -172
rect 6106 -162 6166 6
rect 5710 -222 5720 -172
rect 5640 -292 5720 -222
rect 5640 -352 5650 -292
rect 5710 -352 5720 -292
rect 6096 -222 6106 -172
rect 6562 -162 6622 7
rect 6166 -222 6176 -172
rect 6096 -292 6176 -222
rect 6096 -352 6106 -292
rect 6166 -352 6176 -292
rect 6552 -222 6562 -172
rect 7020 -162 7080 140
rect 7476 8 7536 140
rect 7932 8 7992 140
rect 8406 8 8466 140
rect 8862 8 8922 140
rect 9320 8 9380 140
rect 9776 8 9836 140
rect 10232 8 10292 140
rect 10690 8 10750 140
rect 11146 8 11206 140
rect 11602 8 11662 140
rect 12060 8 12120 140
rect 12516 8 12576 140
rect 12972 8 13032 140
rect 13430 8 13490 140
rect 13886 8 13946 140
rect 14342 8 14402 140
rect 14800 8 14860 140
rect 15209 139 15371 140
rect 15256 8 15316 139
rect 7535 7 7536 8
rect 6622 -222 6632 -172
rect 6552 -292 6632 -222
rect 6552 -352 6562 -292
rect 6622 -352 6632 -292
rect 7010 -222 7020 -172
rect 7476 -162 7536 7
rect 7991 6 7992 8
rect 8465 6 8466 8
rect 7080 -222 7090 -172
rect 7010 -292 7090 -222
rect 7010 -352 7020 -292
rect 7080 -352 7090 -292
rect 7466 -222 7476 -172
rect 7932 -162 7992 6
rect 7536 -222 7546 -172
rect 7466 -292 7546 -222
rect 7466 -352 7476 -292
rect 7536 -352 7546 -292
rect 7922 -222 7932 -172
rect 8406 -162 8466 6
rect 8921 5 8922 8
rect 9379 7 9380 8
rect 7992 -222 8002 -172
rect 7922 -292 8002 -222
rect 7922 -352 7932 -292
rect 7992 -352 8002 -292
rect 8396 -222 8406 -172
rect 8862 -162 8922 5
rect 8466 -222 8476 -172
rect 8396 -292 8476 -222
rect 8396 -352 8406 -292
rect 8466 -352 8476 -292
rect 8852 -222 8862 -172
rect 9320 -162 9380 7
rect 9835 6 9836 8
rect 10291 6 10292 8
rect 8922 -222 8932 -172
rect 8852 -292 8932 -222
rect 8852 -352 8862 -292
rect 8922 -352 8932 -292
rect 9310 -222 9320 -172
rect 9776 -162 9836 6
rect 9380 -222 9390 -172
rect 9310 -292 9390 -222
rect 9310 -352 9320 -292
rect 9380 -352 9390 -292
rect 9766 -222 9776 -172
rect 10232 -162 10292 6
rect 10749 5 10750 8
rect 11205 7 11206 8
rect 9836 -222 9846 -172
rect 9766 -292 9846 -222
rect 9766 -352 9776 -292
rect 9836 -352 9846 -292
rect 10222 -222 10232 -172
rect 10690 -162 10750 5
rect 10292 -222 10302 -172
rect 10222 -292 10302 -222
rect 10222 -352 10232 -292
rect 10292 -352 10302 -292
rect 10680 -222 10690 -172
rect 11146 -162 11206 7
rect 11661 6 11662 8
rect 12119 6 12120 8
rect 12575 7 12576 8
rect 10750 -222 10760 -172
rect 10680 -292 10760 -222
rect 10680 -352 10690 -292
rect 10750 -352 10760 -292
rect 11136 -222 11146 -172
rect 11602 -162 11662 6
rect 11206 -222 11216 -172
rect 11136 -292 11216 -222
rect 11136 -352 11146 -292
rect 11206 -352 11216 -292
rect 11592 -222 11602 -172
rect 12060 -162 12120 6
rect 11662 -222 11672 -172
rect 11592 -292 11672 -222
rect 11592 -352 11602 -292
rect 11662 -352 11672 -292
rect 12050 -222 12060 -172
rect 12516 -162 12576 7
rect 13031 6 13032 8
rect 13489 7 13490 8
rect 13945 7 13946 8
rect 14401 7 14402 8
rect 12120 -222 12130 -172
rect 12050 -292 12130 -222
rect 12050 -352 12060 -292
rect 12120 -352 12130 -292
rect 12506 -222 12516 -172
rect 12972 -162 13032 6
rect 12576 -222 12586 -172
rect 12506 -292 12586 -222
rect 12506 -352 12516 -292
rect 12576 -352 12586 -292
rect 12962 -222 12972 -172
rect 13430 -162 13490 7
rect 13032 -222 13042 -172
rect 12962 -292 13042 -222
rect 12962 -352 12972 -292
rect 13032 -352 13042 -292
rect 13420 -222 13430 -172
rect 13886 -162 13946 7
rect 13490 -222 13500 -172
rect 13420 -292 13500 -222
rect 13420 -352 13430 -292
rect 13490 -352 13500 -292
rect 13876 -222 13886 -172
rect 14342 -162 14402 7
rect 14859 6 14860 8
rect 15315 7 15316 8
rect 13946 -222 13956 -172
rect 13876 -292 13956 -222
rect 13876 -352 13886 -292
rect 13946 -352 13956 -292
rect 14332 -222 14342 -172
rect 14800 -162 14860 6
rect 14402 -222 14412 -172
rect 14332 -292 14412 -222
rect 14332 -352 14342 -292
rect 14402 -352 14412 -292
rect 14790 -222 14800 -172
rect 15256 -162 15316 7
rect 14860 -222 14870 -172
rect 14790 -292 14870 -222
rect 14790 -352 14800 -292
rect 14860 -352 14870 -292
rect 15246 -222 15256 -172
rect 15316 -222 15326 -172
rect 15246 -292 15326 -222
rect 15246 -352 15256 -292
rect 15316 -352 15326 -292
rect 170 -664 230 -352
rect 160 -724 170 -674
rect 626 -664 686 -352
rect 230 -724 240 -674
rect 160 -794 240 -724
rect 160 -854 170 -794
rect 230 -854 240 -794
rect 616 -724 626 -674
rect 1082 -664 1142 -352
rect 686 -724 696 -674
rect 616 -794 696 -724
rect 616 -854 626 -794
rect 686 -854 696 -794
rect 1072 -724 1082 -674
rect 1540 -664 1600 -352
rect 1142 -724 1152 -674
rect 1072 -794 1152 -724
rect 1072 -854 1082 -794
rect 1142 -854 1152 -794
rect 1530 -724 1540 -674
rect 1996 -664 2056 -352
rect 1600 -724 1610 -674
rect 1530 -794 1610 -724
rect 1530 -854 1540 -794
rect 1600 -854 1610 -794
rect 1986 -724 1996 -674
rect 2452 -664 2512 -352
rect 2056 -724 2066 -674
rect 1986 -794 2066 -724
rect 1986 -854 1996 -794
rect 2056 -854 2066 -794
rect 2442 -724 2452 -674
rect 2910 -664 2970 -352
rect 2512 -724 2522 -674
rect 2442 -794 2522 -724
rect 2442 -854 2452 -794
rect 2512 -854 2522 -794
rect 2900 -724 2910 -674
rect 3366 -664 3426 -352
rect 2970 -724 2980 -674
rect 2900 -794 2980 -724
rect 2900 -854 2910 -794
rect 2970 -854 2980 -794
rect 3356 -724 3366 -674
rect 3822 -664 3882 -352
rect 3426 -724 3436 -674
rect 3356 -794 3436 -724
rect 3356 -854 3366 -794
rect 3426 -854 3436 -794
rect 3812 -724 3822 -674
rect 4280 -664 4340 -352
rect 3882 -724 3892 -674
rect 3812 -794 3892 -724
rect 3812 -854 3822 -794
rect 3882 -854 3892 -794
rect 4270 -724 4280 -674
rect 4736 -664 4796 -352
rect 4340 -724 4350 -674
rect 4270 -794 4350 -724
rect 4270 -854 4280 -794
rect 4340 -854 4350 -794
rect 4726 -724 4736 -674
rect 5192 -664 5252 -352
rect 4796 -724 4806 -674
rect 4726 -794 4806 -724
rect 4726 -854 4736 -794
rect 4796 -854 4806 -794
rect 5182 -724 5192 -674
rect 5650 -664 5710 -352
rect 5252 -724 5262 -674
rect 5182 -794 5262 -724
rect 5182 -854 5192 -794
rect 5252 -854 5262 -794
rect 5640 -724 5650 -674
rect 6106 -664 6166 -352
rect 5710 -724 5720 -674
rect 5640 -794 5720 -724
rect 5640 -854 5650 -794
rect 5710 -854 5720 -794
rect 6096 -724 6106 -674
rect 6562 -664 6622 -352
rect 6166 -724 6176 -674
rect 6096 -794 6176 -724
rect 6096 -854 6106 -794
rect 6166 -854 6176 -794
rect 6552 -724 6562 -674
rect 7020 -664 7080 -352
rect 6622 -724 6632 -674
rect 6552 -794 6632 -724
rect 6552 -854 6562 -794
rect 6622 -854 6632 -794
rect 7010 -724 7020 -674
rect 7476 -664 7536 -352
rect 7080 -724 7090 -674
rect 7010 -794 7090 -724
rect 7010 -854 7020 -794
rect 7080 -854 7090 -794
rect 7466 -724 7476 -674
rect 7932 -664 7992 -352
rect 7536 -724 7546 -674
rect 7466 -794 7546 -724
rect 7466 -854 7476 -794
rect 7536 -854 7546 -794
rect 7922 -724 7932 -674
rect 8406 -664 8466 -352
rect 7992 -724 8002 -674
rect 7922 -794 8002 -724
rect 7922 -854 7932 -794
rect 7992 -854 8002 -794
rect 8396 -724 8406 -674
rect 8862 -664 8922 -352
rect 8466 -724 8476 -674
rect 8396 -794 8476 -724
rect 8396 -854 8406 -794
rect 8466 -854 8476 -794
rect 8852 -724 8862 -674
rect 9320 -664 9380 -352
rect 8922 -724 8932 -674
rect 8852 -794 8932 -724
rect 8852 -854 8862 -794
rect 8922 -854 8932 -794
rect 9310 -724 9320 -674
rect 9776 -664 9836 -352
rect 9380 -724 9390 -674
rect 9310 -794 9390 -724
rect 9310 -854 9320 -794
rect 9380 -854 9390 -794
rect 9766 -724 9776 -674
rect 10232 -664 10292 -352
rect 9836 -724 9846 -674
rect 9766 -794 9846 -724
rect 9766 -854 9776 -794
rect 9836 -854 9846 -794
rect 10222 -724 10232 -674
rect 10690 -664 10750 -352
rect 10292 -724 10302 -674
rect 10222 -794 10302 -724
rect 10222 -854 10232 -794
rect 10292 -854 10302 -794
rect 10680 -724 10690 -674
rect 11146 -664 11206 -352
rect 10750 -724 10760 -674
rect 10680 -794 10760 -724
rect 10680 -854 10690 -794
rect 10750 -854 10760 -794
rect 11136 -724 11146 -674
rect 11602 -664 11662 -352
rect 11206 -724 11216 -674
rect 11136 -794 11216 -724
rect 11136 -854 11146 -794
rect 11206 -854 11216 -794
rect 11592 -724 11602 -674
rect 12060 -664 12120 -352
rect 11662 -724 11672 -674
rect 11592 -794 11672 -724
rect 11592 -854 11602 -794
rect 11662 -854 11672 -794
rect 12050 -724 12060 -674
rect 12516 -664 12576 -352
rect 12120 -724 12130 -674
rect 12050 -794 12130 -724
rect 12050 -854 12060 -794
rect 12120 -854 12130 -794
rect 12506 -724 12516 -674
rect 12972 -664 13032 -352
rect 12576 -724 12586 -674
rect 12506 -794 12586 -724
rect 12506 -854 12516 -794
rect 12576 -854 12586 -794
rect 12962 -724 12972 -674
rect 13430 -664 13490 -352
rect 13032 -724 13042 -674
rect 12962 -794 13042 -724
rect 12962 -854 12972 -794
rect 13032 -854 13042 -794
rect 13420 -724 13430 -674
rect 13886 -664 13946 -352
rect 13490 -724 13500 -674
rect 13420 -794 13500 -724
rect 13420 -854 13430 -794
rect 13490 -854 13500 -794
rect 13876 -724 13886 -674
rect 14342 -664 14402 -352
rect 13946 -724 13956 -674
rect 13876 -794 13956 -724
rect 13876 -854 13886 -794
rect 13946 -854 13956 -794
rect 14332 -724 14342 -674
rect 14800 -664 14860 -352
rect 14402 -724 14412 -674
rect 14332 -794 14412 -724
rect 14332 -854 14342 -794
rect 14402 -854 14412 -794
rect 14790 -724 14800 -674
rect 15256 -664 15316 -352
rect 14860 -724 14870 -674
rect 14790 -794 14870 -724
rect 14790 -854 14800 -794
rect 14860 -854 14870 -794
rect 15246 -724 15256 -674
rect 15316 -724 15326 -674
rect 15246 -794 15326 -724
rect 15246 -854 15256 -794
rect 15316 -854 15326 -794
rect 170 -1156 230 -854
rect 160 -1216 170 -1166
rect 626 -1156 686 -854
rect 230 -1216 240 -1166
rect 160 -1286 240 -1216
rect 160 -1346 170 -1286
rect 230 -1346 240 -1286
rect 616 -1216 626 -1166
rect 1082 -1156 1142 -854
rect 686 -1216 696 -1166
rect 616 -1286 696 -1216
rect 616 -1346 626 -1286
rect 686 -1346 696 -1286
rect 1072 -1216 1082 -1166
rect 1540 -1156 1600 -854
rect 1142 -1216 1152 -1166
rect 1072 -1286 1152 -1216
rect 1072 -1346 1082 -1286
rect 1142 -1346 1152 -1286
rect 1530 -1216 1540 -1166
rect 1996 -1156 2056 -854
rect 1600 -1216 1610 -1166
rect 1530 -1286 1610 -1216
rect 1530 -1346 1540 -1286
rect 1600 -1346 1610 -1286
rect 1986 -1216 1996 -1166
rect 2452 -1156 2512 -854
rect 2056 -1216 2066 -1166
rect 1986 -1286 2066 -1216
rect 1986 -1346 1996 -1286
rect 2056 -1346 2066 -1286
rect 2442 -1216 2452 -1166
rect 2910 -1156 2970 -854
rect 2512 -1216 2522 -1166
rect 2442 -1286 2522 -1216
rect 2442 -1346 2452 -1286
rect 2512 -1346 2522 -1286
rect 2900 -1216 2910 -1166
rect 3366 -1156 3426 -854
rect 2970 -1216 2980 -1166
rect 2900 -1286 2980 -1216
rect 2900 -1346 2910 -1286
rect 2970 -1346 2980 -1286
rect 3356 -1216 3366 -1166
rect 3822 -1156 3882 -854
rect 3426 -1216 3436 -1166
rect 3356 -1286 3436 -1216
rect 3356 -1346 3366 -1286
rect 3426 -1346 3436 -1286
rect 3812 -1216 3822 -1166
rect 4280 -1156 4340 -854
rect 3882 -1216 3892 -1166
rect 3812 -1286 3892 -1216
rect 3812 -1346 3822 -1286
rect 3882 -1346 3892 -1286
rect 4270 -1216 4280 -1166
rect 4736 -1156 4796 -854
rect 4340 -1216 4350 -1166
rect 4270 -1286 4350 -1216
rect 4270 -1346 4280 -1286
rect 4340 -1346 4350 -1286
rect 4726 -1216 4736 -1166
rect 5192 -1156 5252 -854
rect 4796 -1216 4806 -1166
rect 4726 -1286 4806 -1216
rect 4726 -1346 4736 -1286
rect 4796 -1346 4806 -1286
rect 5182 -1216 5192 -1166
rect 5650 -1156 5710 -854
rect 5252 -1216 5262 -1166
rect 5182 -1286 5262 -1216
rect 5182 -1346 5192 -1286
rect 5252 -1346 5262 -1286
rect 5640 -1216 5650 -1166
rect 6106 -1156 6166 -854
rect 5710 -1216 5720 -1166
rect 5640 -1286 5720 -1216
rect 5640 -1346 5650 -1286
rect 5710 -1346 5720 -1286
rect 6096 -1216 6106 -1166
rect 6562 -1156 6622 -854
rect 6166 -1216 6176 -1166
rect 6096 -1286 6176 -1216
rect 6096 -1346 6106 -1286
rect 6166 -1346 6176 -1286
rect 6552 -1216 6562 -1166
rect 7020 -1156 7080 -854
rect 6622 -1216 6632 -1166
rect 6552 -1286 6632 -1216
rect 6552 -1346 6562 -1286
rect 6622 -1346 6632 -1286
rect 7010 -1216 7020 -1166
rect 7476 -1156 7536 -854
rect 7080 -1216 7090 -1166
rect 7010 -1286 7090 -1216
rect 7010 -1346 7020 -1286
rect 7080 -1346 7090 -1286
rect 7466 -1216 7476 -1166
rect 7932 -1156 7992 -854
rect 7536 -1216 7546 -1166
rect 7466 -1286 7546 -1216
rect 7466 -1346 7476 -1286
rect 7536 -1346 7546 -1286
rect 7922 -1216 7932 -1166
rect 8406 -1156 8466 -854
rect 7992 -1216 8002 -1166
rect 7922 -1286 8002 -1216
rect 7922 -1346 7932 -1286
rect 7992 -1346 8002 -1286
rect 8396 -1216 8406 -1166
rect 8862 -1156 8922 -854
rect 8466 -1216 8476 -1166
rect 8396 -1286 8476 -1216
rect 8396 -1346 8406 -1286
rect 8466 -1346 8476 -1286
rect 8852 -1216 8862 -1166
rect 9320 -1156 9380 -854
rect 8922 -1216 8932 -1166
rect 8852 -1286 8932 -1216
rect 8852 -1346 8862 -1286
rect 8922 -1346 8932 -1286
rect 9310 -1216 9320 -1166
rect 9776 -1156 9836 -854
rect 9380 -1216 9390 -1166
rect 9310 -1286 9390 -1216
rect 9310 -1346 9320 -1286
rect 9380 -1346 9390 -1286
rect 9766 -1216 9776 -1166
rect 10232 -1156 10292 -854
rect 9836 -1216 9846 -1166
rect 9766 -1286 9846 -1216
rect 9766 -1346 9776 -1286
rect 9836 -1346 9846 -1286
rect 10222 -1216 10232 -1166
rect 10690 -1156 10750 -854
rect 10292 -1216 10302 -1166
rect 10222 -1286 10302 -1216
rect 10222 -1346 10232 -1286
rect 10292 -1346 10302 -1286
rect 10680 -1216 10690 -1166
rect 11146 -1156 11206 -854
rect 10750 -1216 10760 -1166
rect 10680 -1286 10760 -1216
rect 10680 -1346 10690 -1286
rect 10750 -1346 10760 -1286
rect 11136 -1216 11146 -1166
rect 11602 -1156 11662 -854
rect 11206 -1216 11216 -1166
rect 11136 -1286 11216 -1216
rect 11136 -1346 11146 -1286
rect 11206 -1346 11216 -1286
rect 11592 -1216 11602 -1166
rect 12060 -1156 12120 -854
rect 11662 -1216 11672 -1166
rect 11592 -1286 11672 -1216
rect 11592 -1346 11602 -1286
rect 11662 -1346 11672 -1286
rect 12050 -1216 12060 -1166
rect 12516 -1156 12576 -854
rect 12120 -1216 12130 -1166
rect 12050 -1286 12130 -1216
rect 12050 -1346 12060 -1286
rect 12120 -1346 12130 -1286
rect 12506 -1216 12516 -1166
rect 12972 -1156 13032 -854
rect 12576 -1216 12586 -1166
rect 12506 -1286 12586 -1216
rect 12506 -1346 12516 -1286
rect 12576 -1346 12586 -1286
rect 12962 -1216 12972 -1166
rect 13430 -1156 13490 -854
rect 13032 -1216 13042 -1166
rect 12962 -1286 13042 -1216
rect 12962 -1346 12972 -1286
rect 13032 -1346 13042 -1286
rect 13420 -1216 13430 -1166
rect 13886 -1156 13946 -854
rect 13490 -1216 13500 -1166
rect 13420 -1286 13500 -1216
rect 13420 -1346 13430 -1286
rect 13490 -1346 13500 -1286
rect 13876 -1216 13886 -1166
rect 14342 -1156 14402 -854
rect 13946 -1216 13956 -1166
rect 13876 -1286 13956 -1216
rect 13876 -1346 13886 -1286
rect 13946 -1346 13956 -1286
rect 14332 -1216 14342 -1166
rect 14800 -1156 14860 -854
rect 14402 -1216 14412 -1166
rect 14332 -1286 14412 -1216
rect 14332 -1346 14342 -1286
rect 14402 -1346 14412 -1286
rect 14790 -1216 14800 -1166
rect 15256 -1156 15316 -854
rect 14860 -1216 14870 -1166
rect 14790 -1286 14870 -1216
rect 14790 -1346 14800 -1286
rect 14860 -1346 14870 -1286
rect 15246 -1216 15256 -1166
rect 15316 -1216 15326 -1166
rect 15246 -1286 15326 -1216
rect 15246 -1346 15256 -1286
rect 15316 -1346 15326 -1286
rect 170 -1672 230 -1346
rect 160 -1732 170 -1682
rect 626 -1672 686 -1346
rect 230 -1732 240 -1682
rect 160 -1802 240 -1732
rect 160 -1862 170 -1802
rect 230 -1862 240 -1802
rect 616 -1732 626 -1682
rect 1082 -1672 1142 -1346
rect 686 -1732 696 -1682
rect 616 -1802 696 -1732
rect 616 -1862 626 -1802
rect 686 -1862 696 -1802
rect 1072 -1732 1082 -1682
rect 1540 -1672 1600 -1346
rect 1142 -1732 1152 -1682
rect 1072 -1802 1152 -1732
rect 1072 -1862 1082 -1802
rect 1142 -1862 1152 -1802
rect 1530 -1732 1540 -1682
rect 1996 -1672 2056 -1346
rect 1600 -1732 1610 -1682
rect 1530 -1802 1610 -1732
rect 1530 -1862 1540 -1802
rect 1600 -1862 1610 -1802
rect 1986 -1732 1996 -1682
rect 2452 -1672 2512 -1346
rect 2056 -1732 2066 -1682
rect 1986 -1802 2066 -1732
rect 1986 -1862 1996 -1802
rect 2056 -1862 2066 -1802
rect 2442 -1732 2452 -1682
rect 2910 -1672 2970 -1346
rect 2512 -1732 2522 -1682
rect 2442 -1802 2522 -1732
rect 2442 -1862 2452 -1802
rect 2512 -1862 2522 -1802
rect 2900 -1732 2910 -1682
rect 3366 -1672 3426 -1346
rect 2970 -1732 2980 -1682
rect 2900 -1802 2980 -1732
rect 2900 -1862 2910 -1802
rect 2970 -1862 2980 -1802
rect 3356 -1732 3366 -1682
rect 3822 -1672 3882 -1346
rect 3426 -1732 3436 -1682
rect 3356 -1802 3436 -1732
rect 3356 -1862 3366 -1802
rect 3426 -1862 3436 -1802
rect 3812 -1732 3822 -1682
rect 4280 -1672 4340 -1346
rect 3882 -1732 3892 -1682
rect 3812 -1802 3892 -1732
rect 3812 -1862 3822 -1802
rect 3882 -1862 3892 -1802
rect 4270 -1732 4280 -1682
rect 4736 -1672 4796 -1346
rect 4340 -1732 4350 -1682
rect 4270 -1802 4350 -1732
rect 4270 -1862 4280 -1802
rect 4340 -1862 4350 -1802
rect 4726 -1732 4736 -1682
rect 5192 -1672 5252 -1346
rect 4796 -1732 4806 -1682
rect 4726 -1802 4806 -1732
rect 4726 -1862 4736 -1802
rect 4796 -1862 4806 -1802
rect 5182 -1732 5192 -1682
rect 5650 -1672 5710 -1346
rect 5252 -1732 5262 -1682
rect 5182 -1802 5262 -1732
rect 5182 -1862 5192 -1802
rect 5252 -1862 5262 -1802
rect 5640 -1732 5650 -1682
rect 6106 -1672 6166 -1346
rect 5710 -1732 5720 -1682
rect 5640 -1802 5720 -1732
rect 5640 -1862 5650 -1802
rect 5710 -1862 5720 -1802
rect 6096 -1732 6106 -1682
rect 6562 -1672 6622 -1346
rect 6166 -1732 6176 -1682
rect 6096 -1802 6176 -1732
rect 6096 -1862 6106 -1802
rect 6166 -1862 6176 -1802
rect 6552 -1732 6562 -1682
rect 7020 -1672 7080 -1346
rect 6622 -1732 6632 -1682
rect 6552 -1802 6632 -1732
rect 6552 -1862 6562 -1802
rect 6622 -1862 6632 -1802
rect 7010 -1732 7020 -1682
rect 7476 -1672 7536 -1346
rect 7080 -1732 7090 -1682
rect 7010 -1802 7090 -1732
rect 7010 -1862 7020 -1802
rect 7080 -1862 7090 -1802
rect 7466 -1732 7476 -1682
rect 7932 -1672 7992 -1346
rect 7536 -1732 7546 -1682
rect 7466 -1802 7546 -1732
rect 7466 -1862 7476 -1802
rect 7536 -1862 7546 -1802
rect 7922 -1732 7932 -1682
rect 8406 -1672 8466 -1346
rect 7992 -1732 8002 -1682
rect 7922 -1802 8002 -1732
rect 7922 -1862 7932 -1802
rect 7992 -1862 8002 -1802
rect 8396 -1732 8406 -1682
rect 8862 -1672 8922 -1346
rect 8466 -1732 8476 -1682
rect 8396 -1802 8476 -1732
rect 8396 -1862 8406 -1802
rect 8466 -1862 8476 -1802
rect 8852 -1732 8862 -1682
rect 9320 -1672 9380 -1346
rect 8922 -1732 8932 -1682
rect 8852 -1802 8932 -1732
rect 8852 -1862 8862 -1802
rect 8922 -1862 8932 -1802
rect 9310 -1732 9320 -1682
rect 9776 -1672 9836 -1346
rect 9380 -1732 9390 -1682
rect 9310 -1802 9390 -1732
rect 9310 -1862 9320 -1802
rect 9380 -1862 9390 -1802
rect 9766 -1732 9776 -1682
rect 10232 -1672 10292 -1346
rect 9836 -1732 9846 -1682
rect 9766 -1802 9846 -1732
rect 9766 -1862 9776 -1802
rect 9836 -1862 9846 -1802
rect 10222 -1732 10232 -1682
rect 10690 -1672 10750 -1346
rect 10292 -1732 10302 -1682
rect 10222 -1802 10302 -1732
rect 10222 -1862 10232 -1802
rect 10292 -1862 10302 -1802
rect 10680 -1732 10690 -1682
rect 11146 -1672 11206 -1346
rect 10750 -1732 10760 -1682
rect 10680 -1802 10760 -1732
rect 10680 -1862 10690 -1802
rect 10750 -1862 10760 -1802
rect 11136 -1732 11146 -1682
rect 11602 -1672 11662 -1346
rect 11206 -1732 11216 -1682
rect 11136 -1802 11216 -1732
rect 11136 -1862 11146 -1802
rect 11206 -1862 11216 -1802
rect 11592 -1732 11602 -1682
rect 12060 -1672 12120 -1346
rect 11662 -1732 11672 -1682
rect 11592 -1802 11672 -1732
rect 11592 -1862 11602 -1802
rect 11662 -1862 11672 -1802
rect 12050 -1732 12060 -1682
rect 12516 -1672 12576 -1346
rect 12120 -1732 12130 -1682
rect 12050 -1802 12130 -1732
rect 12050 -1862 12060 -1802
rect 12120 -1862 12130 -1802
rect 12506 -1732 12516 -1682
rect 12972 -1672 13032 -1346
rect 12576 -1732 12586 -1682
rect 12506 -1802 12586 -1732
rect 12506 -1862 12516 -1802
rect 12576 -1862 12586 -1802
rect 12962 -1732 12972 -1682
rect 13430 -1672 13490 -1346
rect 13032 -1732 13042 -1682
rect 12962 -1802 13042 -1732
rect 12962 -1862 12972 -1802
rect 13032 -1862 13042 -1802
rect 13420 -1732 13430 -1682
rect 13886 -1672 13946 -1346
rect 13490 -1732 13500 -1682
rect 13420 -1802 13500 -1732
rect 13420 -1862 13430 -1802
rect 13490 -1862 13500 -1802
rect 13876 -1732 13886 -1682
rect 14342 -1672 14402 -1346
rect 13946 -1732 13956 -1682
rect 13876 -1802 13956 -1732
rect 13876 -1862 13886 -1802
rect 13946 -1862 13956 -1802
rect 14332 -1732 14342 -1682
rect 14800 -1672 14860 -1346
rect 14402 -1732 14412 -1682
rect 14332 -1802 14412 -1732
rect 14332 -1862 14342 -1802
rect 14402 -1862 14412 -1802
rect 14790 -1732 14800 -1682
rect 15256 -1672 15316 -1346
rect 14860 -1732 14870 -1682
rect 14790 -1802 14870 -1732
rect 14790 -1862 14800 -1802
rect 14860 -1862 14870 -1802
rect 15246 -1732 15256 -1682
rect 15316 -1732 15326 -1682
rect 15246 -1802 15326 -1732
rect 15246 -1862 15256 -1802
rect 15316 -1862 15326 -1802
rect 170 -2174 230 -1862
rect 160 -2234 170 -2184
rect 626 -2174 686 -1862
rect 230 -2234 240 -2184
rect 160 -2304 240 -2234
rect 160 -2364 170 -2304
rect 230 -2364 240 -2304
rect 616 -2234 626 -2184
rect 1082 -2174 1142 -1862
rect 686 -2234 696 -2184
rect 616 -2304 696 -2234
rect 616 -2364 626 -2304
rect 686 -2364 696 -2304
rect 1072 -2234 1082 -2184
rect 1540 -2174 1600 -1862
rect 1142 -2234 1152 -2184
rect 1072 -2304 1152 -2234
rect 1072 -2364 1082 -2304
rect 1142 -2364 1152 -2304
rect 1530 -2234 1540 -2184
rect 1996 -2174 2056 -1862
rect 1600 -2234 1610 -2184
rect 1530 -2304 1610 -2234
rect 1530 -2364 1540 -2304
rect 1600 -2364 1610 -2304
rect 1986 -2234 1996 -2184
rect 2452 -2174 2512 -1862
rect 2056 -2234 2066 -2184
rect 1986 -2304 2066 -2234
rect 1986 -2364 1996 -2304
rect 2056 -2364 2066 -2304
rect 2442 -2234 2452 -2184
rect 2910 -2174 2970 -1862
rect 2512 -2234 2522 -2184
rect 2442 -2304 2522 -2234
rect 2442 -2364 2452 -2304
rect 2512 -2364 2522 -2304
rect 2900 -2234 2910 -2184
rect 3366 -2174 3426 -1862
rect 2970 -2234 2980 -2184
rect 2900 -2304 2980 -2234
rect 2900 -2364 2910 -2304
rect 2970 -2364 2980 -2304
rect 3356 -2234 3366 -2184
rect 3822 -2174 3882 -1862
rect 3426 -2234 3436 -2184
rect 3356 -2304 3436 -2234
rect 3356 -2364 3366 -2304
rect 3426 -2364 3436 -2304
rect 3812 -2234 3822 -2184
rect 4280 -2174 4340 -1862
rect 3882 -2234 3892 -2184
rect 3812 -2304 3892 -2234
rect 3812 -2364 3822 -2304
rect 3882 -2364 3892 -2304
rect 4270 -2234 4280 -2184
rect 4736 -2174 4796 -1862
rect 4340 -2234 4350 -2184
rect 4270 -2304 4350 -2234
rect 4270 -2364 4280 -2304
rect 4340 -2364 4350 -2304
rect 4726 -2234 4736 -2184
rect 5192 -2174 5252 -1862
rect 4796 -2234 4806 -2184
rect 4726 -2304 4806 -2234
rect 4726 -2364 4736 -2304
rect 4796 -2364 4806 -2304
rect 5182 -2234 5192 -2184
rect 5650 -2174 5710 -1862
rect 5252 -2234 5262 -2184
rect 5182 -2304 5262 -2234
rect 5182 -2364 5192 -2304
rect 5252 -2364 5262 -2304
rect 5640 -2234 5650 -2184
rect 6106 -2174 6166 -1862
rect 5710 -2234 5720 -2184
rect 5640 -2304 5720 -2234
rect 5640 -2364 5650 -2304
rect 5710 -2364 5720 -2304
rect 6096 -2234 6106 -2184
rect 6562 -2174 6622 -1862
rect 6166 -2234 6176 -2184
rect 6096 -2304 6176 -2234
rect 6096 -2364 6106 -2304
rect 6166 -2364 6176 -2304
rect 6552 -2234 6562 -2184
rect 7020 -2174 7080 -1862
rect 6622 -2234 6632 -2184
rect 6552 -2304 6632 -2234
rect 6552 -2364 6562 -2304
rect 6622 -2364 6632 -2304
rect 7010 -2234 7020 -2184
rect 7476 -2174 7536 -1862
rect 7080 -2234 7090 -2184
rect 7010 -2304 7090 -2234
rect 7010 -2364 7020 -2304
rect 7080 -2364 7090 -2304
rect 7466 -2234 7476 -2184
rect 7932 -2174 7992 -1862
rect 7536 -2234 7546 -2184
rect 7466 -2304 7546 -2234
rect 7466 -2364 7476 -2304
rect 7536 -2364 7546 -2304
rect 7922 -2234 7932 -2184
rect 8406 -2174 8466 -1862
rect 7992 -2234 8002 -2184
rect 7922 -2304 8002 -2234
rect 7922 -2364 7932 -2304
rect 7992 -2364 8002 -2304
rect 8396 -2234 8406 -2184
rect 8862 -2174 8922 -1862
rect 8466 -2234 8476 -2184
rect 8396 -2304 8476 -2234
rect 8396 -2364 8406 -2304
rect 8466 -2364 8476 -2304
rect 8852 -2234 8862 -2184
rect 9320 -2174 9380 -1862
rect 8922 -2234 8932 -2184
rect 8852 -2304 8932 -2234
rect 8852 -2364 8862 -2304
rect 8922 -2364 8932 -2304
rect 9310 -2234 9320 -2184
rect 9776 -2174 9836 -1862
rect 9380 -2234 9390 -2184
rect 9310 -2304 9390 -2234
rect 9310 -2364 9320 -2304
rect 9380 -2364 9390 -2304
rect 9766 -2234 9776 -2184
rect 10232 -2174 10292 -1862
rect 9836 -2234 9846 -2184
rect 9766 -2304 9846 -2234
rect 9766 -2364 9776 -2304
rect 9836 -2364 9846 -2304
rect 10222 -2234 10232 -2184
rect 10690 -2174 10750 -1862
rect 10292 -2234 10302 -2184
rect 10222 -2304 10302 -2234
rect 10222 -2364 10232 -2304
rect 10292 -2364 10302 -2304
rect 10680 -2234 10690 -2184
rect 11146 -2174 11206 -1862
rect 10750 -2234 10760 -2184
rect 10680 -2304 10760 -2234
rect 10680 -2364 10690 -2304
rect 10750 -2364 10760 -2304
rect 11136 -2234 11146 -2184
rect 11602 -2174 11662 -1862
rect 11206 -2234 11216 -2184
rect 11136 -2304 11216 -2234
rect 11136 -2364 11146 -2304
rect 11206 -2364 11216 -2304
rect 11592 -2234 11602 -2184
rect 12060 -2174 12120 -1862
rect 11662 -2234 11672 -2184
rect 11592 -2304 11672 -2234
rect 11592 -2364 11602 -2304
rect 11662 -2364 11672 -2304
rect 12050 -2234 12060 -2184
rect 12516 -2174 12576 -1862
rect 12120 -2234 12130 -2184
rect 12050 -2304 12130 -2234
rect 12050 -2364 12060 -2304
rect 12120 -2364 12130 -2304
rect 12506 -2234 12516 -2184
rect 12972 -2174 13032 -1862
rect 12576 -2234 12586 -2184
rect 12506 -2304 12586 -2234
rect 12506 -2364 12516 -2304
rect 12576 -2364 12586 -2304
rect 12962 -2234 12972 -2184
rect 13430 -2174 13490 -1862
rect 13032 -2234 13042 -2184
rect 12962 -2304 13042 -2234
rect 12962 -2364 12972 -2304
rect 13032 -2364 13042 -2304
rect 13420 -2234 13430 -2184
rect 13886 -2174 13946 -1862
rect 13490 -2234 13500 -2184
rect 13420 -2304 13500 -2234
rect 13420 -2364 13430 -2304
rect 13490 -2364 13500 -2304
rect 13876 -2234 13886 -2184
rect 14342 -2174 14402 -1862
rect 13946 -2234 13956 -2184
rect 13876 -2304 13956 -2234
rect 13876 -2364 13886 -2304
rect 13946 -2364 13956 -2304
rect 14332 -2234 14342 -2184
rect 14800 -2174 14860 -1862
rect 14402 -2234 14412 -2184
rect 14332 -2304 14412 -2234
rect 14332 -2364 14342 -2304
rect 14402 -2364 14412 -2304
rect 14790 -2234 14800 -2184
rect 15256 -2174 15316 -1862
rect 14860 -2234 14870 -2184
rect 14790 -2304 14870 -2234
rect 14790 -2364 14800 -2304
rect 14860 -2364 14870 -2304
rect 15246 -2234 15256 -2184
rect 15316 -2234 15326 -2184
rect 15246 -2304 15326 -2234
rect 15246 -2364 15256 -2304
rect 15316 -2364 15326 -2304
rect 170 -2666 230 -2364
rect 160 -2726 170 -2676
rect 626 -2666 686 -2364
rect 230 -2726 240 -2676
rect 160 -2796 240 -2726
rect 160 -2856 170 -2796
rect 230 -2856 240 -2796
rect 616 -2726 626 -2676
rect 1082 -2666 1142 -2364
rect 686 -2726 696 -2676
rect 616 -2796 696 -2726
rect 616 -2856 626 -2796
rect 686 -2856 696 -2796
rect 1072 -2726 1082 -2676
rect 1540 -2666 1600 -2364
rect 1142 -2726 1152 -2676
rect 1072 -2796 1152 -2726
rect 1072 -2856 1082 -2796
rect 1142 -2856 1152 -2796
rect 1530 -2726 1540 -2676
rect 1996 -2666 2056 -2364
rect 1600 -2726 1610 -2676
rect 1530 -2796 1610 -2726
rect 1530 -2856 1540 -2796
rect 1600 -2856 1610 -2796
rect 1986 -2726 1996 -2676
rect 2452 -2666 2512 -2364
rect 2056 -2726 2066 -2676
rect 1986 -2796 2066 -2726
rect 1986 -2856 1996 -2796
rect 2056 -2856 2066 -2796
rect 2442 -2726 2452 -2676
rect 2910 -2666 2970 -2364
rect 2512 -2726 2522 -2676
rect 2442 -2796 2522 -2726
rect 2442 -2856 2452 -2796
rect 2512 -2856 2522 -2796
rect 2900 -2726 2910 -2676
rect 3366 -2666 3426 -2364
rect 2970 -2726 2980 -2676
rect 2900 -2796 2980 -2726
rect 2900 -2856 2910 -2796
rect 2970 -2856 2980 -2796
rect 3356 -2726 3366 -2676
rect 3822 -2666 3882 -2364
rect 3426 -2726 3436 -2676
rect 3356 -2796 3436 -2726
rect 3356 -2856 3366 -2796
rect 3426 -2856 3436 -2796
rect 3812 -2726 3822 -2676
rect 4280 -2666 4340 -2364
rect 3882 -2726 3892 -2676
rect 3812 -2796 3892 -2726
rect 3812 -2856 3822 -2796
rect 3882 -2856 3892 -2796
rect 4270 -2726 4280 -2676
rect 4736 -2666 4796 -2364
rect 4340 -2726 4350 -2676
rect 4270 -2796 4350 -2726
rect 4270 -2856 4280 -2796
rect 4340 -2856 4350 -2796
rect 4726 -2726 4736 -2676
rect 5192 -2666 5252 -2364
rect 4796 -2726 4806 -2676
rect 4726 -2796 4806 -2726
rect 4726 -2856 4736 -2796
rect 4796 -2856 4806 -2796
rect 5182 -2726 5192 -2676
rect 5650 -2666 5710 -2364
rect 5252 -2726 5262 -2676
rect 5182 -2796 5262 -2726
rect 5182 -2856 5192 -2796
rect 5252 -2856 5262 -2796
rect 5640 -2726 5650 -2676
rect 6106 -2666 6166 -2364
rect 5710 -2726 5720 -2676
rect 5640 -2796 5720 -2726
rect 5640 -2856 5650 -2796
rect 5710 -2856 5720 -2796
rect 6096 -2726 6106 -2676
rect 6562 -2666 6622 -2364
rect 6166 -2726 6176 -2676
rect 6096 -2796 6176 -2726
rect 6096 -2856 6106 -2796
rect 6166 -2856 6176 -2796
rect 6552 -2726 6562 -2676
rect 7020 -2666 7080 -2364
rect 6622 -2726 6632 -2676
rect 6552 -2796 6632 -2726
rect 6552 -2856 6562 -2796
rect 6622 -2856 6632 -2796
rect 7010 -2726 7020 -2676
rect 7476 -2666 7536 -2364
rect 7080 -2726 7090 -2676
rect 7010 -2796 7090 -2726
rect 7010 -2856 7020 -2796
rect 7080 -2856 7090 -2796
rect 7466 -2726 7476 -2676
rect 7932 -2666 7992 -2364
rect 7536 -2726 7546 -2676
rect 7466 -2796 7546 -2726
rect 7466 -2856 7476 -2796
rect 7536 -2856 7546 -2796
rect 7922 -2726 7932 -2676
rect 8406 -2666 8466 -2364
rect 7992 -2726 8002 -2676
rect 7922 -2796 8002 -2726
rect 7922 -2856 7932 -2796
rect 7992 -2856 8002 -2796
rect 8396 -2726 8406 -2676
rect 8862 -2666 8922 -2364
rect 8466 -2726 8476 -2676
rect 8396 -2796 8476 -2726
rect 8396 -2856 8406 -2796
rect 8466 -2856 8476 -2796
rect 8852 -2726 8862 -2676
rect 9320 -2666 9380 -2364
rect 8922 -2726 8932 -2676
rect 8852 -2796 8932 -2726
rect 8852 -2856 8862 -2796
rect 8922 -2856 8932 -2796
rect 9310 -2726 9320 -2676
rect 9776 -2666 9836 -2364
rect 9380 -2726 9390 -2676
rect 9310 -2796 9390 -2726
rect 9310 -2856 9320 -2796
rect 9380 -2856 9390 -2796
rect 9766 -2726 9776 -2676
rect 10232 -2666 10292 -2364
rect 9836 -2726 9846 -2676
rect 9766 -2796 9846 -2726
rect 9766 -2856 9776 -2796
rect 9836 -2856 9846 -2796
rect 10222 -2726 10232 -2676
rect 10690 -2666 10750 -2364
rect 10292 -2726 10302 -2676
rect 10222 -2796 10302 -2726
rect 10222 -2856 10232 -2796
rect 10292 -2856 10302 -2796
rect 10680 -2726 10690 -2676
rect 11146 -2666 11206 -2364
rect 10750 -2726 10760 -2676
rect 10680 -2796 10760 -2726
rect 10680 -2856 10690 -2796
rect 10750 -2856 10760 -2796
rect 11136 -2726 11146 -2676
rect 11602 -2666 11662 -2364
rect 11206 -2726 11216 -2676
rect 11136 -2796 11216 -2726
rect 11136 -2856 11146 -2796
rect 11206 -2856 11216 -2796
rect 11592 -2726 11602 -2676
rect 12060 -2666 12120 -2364
rect 11662 -2726 11672 -2676
rect 11592 -2796 11672 -2726
rect 11592 -2856 11602 -2796
rect 11662 -2856 11672 -2796
rect 12050 -2726 12060 -2676
rect 12516 -2666 12576 -2364
rect 12120 -2726 12130 -2676
rect 12050 -2796 12130 -2726
rect 12050 -2856 12060 -2796
rect 12120 -2856 12130 -2796
rect 12506 -2726 12516 -2676
rect 12972 -2666 13032 -2364
rect 12576 -2726 12586 -2676
rect 12506 -2796 12586 -2726
rect 12506 -2856 12516 -2796
rect 12576 -2856 12586 -2796
rect 12962 -2726 12972 -2676
rect 13430 -2666 13490 -2364
rect 13032 -2726 13042 -2676
rect 12962 -2796 13042 -2726
rect 12962 -2856 12972 -2796
rect 13032 -2856 13042 -2796
rect 13420 -2726 13430 -2676
rect 13886 -2666 13946 -2364
rect 13490 -2726 13500 -2676
rect 13420 -2796 13500 -2726
rect 13420 -2856 13430 -2796
rect 13490 -2856 13500 -2796
rect 13876 -2726 13886 -2676
rect 14342 -2666 14402 -2364
rect 13946 -2726 13956 -2676
rect 13876 -2796 13956 -2726
rect 13876 -2856 13886 -2796
rect 13946 -2856 13956 -2796
rect 14332 -2726 14342 -2676
rect 14800 -2666 14860 -2364
rect 14402 -2726 14412 -2676
rect 14332 -2796 14412 -2726
rect 14332 -2856 14342 -2796
rect 14402 -2856 14412 -2796
rect 14790 -2726 14800 -2676
rect 15256 -2666 15316 -2364
rect 14860 -2726 14870 -2676
rect 14790 -2796 14870 -2726
rect 14790 -2856 14800 -2796
rect 14860 -2856 14870 -2796
rect 15246 -2726 15256 -2676
rect 15316 -2726 15326 -2676
rect 15246 -2796 15326 -2726
rect 15246 -2856 15256 -2796
rect 15316 -2856 15326 -2796
rect 170 -3034 230 -2856
rect 626 -3034 686 -2856
rect 1082 -3034 1142 -2856
rect 1540 -3035 1600 -2856
rect 1996 -3032 2056 -2856
rect 2452 -3033 2512 -2856
rect 2910 -3033 2970 -2856
rect 3366 -3033 3426 -2856
rect 3822 -3034 3882 -2856
rect 4280 -3033 4340 -2856
rect 4736 -3034 4796 -2856
rect 5192 -3034 5252 -2856
rect 5650 -3034 5710 -2856
rect 6106 -3034 6166 -2856
rect 6562 -3034 6622 -2856
rect 7020 -3035 7080 -2856
rect 7476 -3034 7536 -2856
rect 7932 -3034 7992 -2856
rect 8406 -3034 8466 -2856
rect 8862 -3035 8922 -2856
rect 9320 -3034 9380 -2856
rect 9776 -3035 9836 -2856
rect 10232 -3034 10292 -2856
rect 10690 -3034 10750 -2856
rect 11146 -3033 11206 -2856
rect 11602 -3034 11662 -2856
rect 12060 -3034 12120 -2856
rect 12516 -3034 12576 -2856
rect 12972 -3034 13032 -2856
rect 13430 -3034 13490 -2856
rect 13886 -3034 13946 -2856
rect 14342 -3034 14402 -2856
rect 14800 -3033 14860 -2856
rect 15256 -3034 15316 -2856
rect 170 -3662 230 -3470
rect 160 -3722 170 -3672
rect 626 -3662 686 -3470
rect 230 -3722 240 -3672
rect 160 -3792 240 -3722
rect 160 -3852 170 -3792
rect 230 -3852 240 -3792
rect 616 -3722 626 -3672
rect 1082 -3662 1142 -3470
rect 686 -3722 696 -3672
rect 616 -3792 696 -3722
rect 616 -3852 626 -3792
rect 686 -3852 696 -3792
rect 1072 -3722 1082 -3672
rect 1540 -3662 1600 -3470
rect 1142 -3722 1152 -3672
rect 1072 -3792 1152 -3722
rect 1072 -3852 1082 -3792
rect 1142 -3852 1152 -3792
rect 1530 -3722 1540 -3672
rect 1996 -3662 2056 -3470
rect 1600 -3722 1610 -3672
rect 1530 -3792 1610 -3722
rect 1530 -3852 1540 -3792
rect 1600 -3852 1610 -3792
rect 1986 -3722 1996 -3672
rect 2452 -3662 2512 -3470
rect 2056 -3722 2066 -3672
rect 1986 -3792 2066 -3722
rect 1986 -3852 1996 -3792
rect 2056 -3852 2066 -3792
rect 2442 -3722 2452 -3672
rect 2910 -3662 2970 -3470
rect 2512 -3722 2522 -3672
rect 2442 -3792 2522 -3722
rect 2442 -3852 2452 -3792
rect 2512 -3852 2522 -3792
rect 2900 -3722 2910 -3672
rect 3366 -3662 3426 -3470
rect 2970 -3722 2980 -3672
rect 2900 -3792 2980 -3722
rect 2900 -3852 2910 -3792
rect 2970 -3852 2980 -3792
rect 3356 -3722 3366 -3672
rect 3822 -3662 3882 -3470
rect 3426 -3722 3436 -3672
rect 3356 -3792 3436 -3722
rect 3356 -3852 3366 -3792
rect 3426 -3852 3436 -3792
rect 3812 -3722 3822 -3672
rect 4280 -3662 4340 -3470
rect 3882 -3722 3892 -3672
rect 3812 -3792 3892 -3722
rect 3812 -3852 3822 -3792
rect 3882 -3852 3892 -3792
rect 4270 -3722 4280 -3672
rect 4736 -3662 4796 -3470
rect 4340 -3722 4350 -3672
rect 4270 -3792 4350 -3722
rect 4270 -3852 4280 -3792
rect 4340 -3852 4350 -3792
rect 4726 -3722 4736 -3672
rect 5192 -3662 5252 -3470
rect 4796 -3722 4806 -3672
rect 4726 -3792 4806 -3722
rect 4726 -3852 4736 -3792
rect 4796 -3852 4806 -3792
rect 5182 -3722 5192 -3672
rect 5650 -3662 5710 -3470
rect 5252 -3722 5262 -3672
rect 5182 -3792 5262 -3722
rect 5182 -3852 5192 -3792
rect 5252 -3852 5262 -3792
rect 5640 -3722 5650 -3672
rect 6106 -3662 6166 -3470
rect 5710 -3722 5720 -3672
rect 5640 -3792 5720 -3722
rect 5640 -3852 5650 -3792
rect 5710 -3852 5720 -3792
rect 6096 -3722 6106 -3672
rect 6562 -3662 6622 -3470
rect 6166 -3722 6176 -3672
rect 6096 -3792 6176 -3722
rect 6096 -3852 6106 -3792
rect 6166 -3852 6176 -3792
rect 6552 -3722 6562 -3672
rect 7020 -3662 7080 -3470
rect 6622 -3722 6632 -3672
rect 6552 -3792 6632 -3722
rect 6552 -3852 6562 -3792
rect 6622 -3852 6632 -3792
rect 7010 -3722 7020 -3672
rect 7476 -3662 7536 -3470
rect 7080 -3722 7090 -3672
rect 7010 -3792 7090 -3722
rect 7010 -3852 7020 -3792
rect 7080 -3852 7090 -3792
rect 7466 -3722 7476 -3672
rect 7932 -3662 7992 -3470
rect 7536 -3722 7546 -3672
rect 7466 -3792 7546 -3722
rect 7466 -3852 7476 -3792
rect 7536 -3852 7546 -3792
rect 7922 -3722 7932 -3672
rect 8406 -3662 8466 -3470
rect 7992 -3722 8002 -3672
rect 7922 -3792 8002 -3722
rect 7922 -3852 7932 -3792
rect 7992 -3852 8002 -3792
rect 8396 -3722 8406 -3672
rect 8862 -3662 8922 -3470
rect 8466 -3722 8476 -3672
rect 8396 -3792 8476 -3722
rect 8396 -3852 8406 -3792
rect 8466 -3852 8476 -3792
rect 8852 -3722 8862 -3672
rect 9320 -3662 9380 -3470
rect 8922 -3722 8932 -3672
rect 8852 -3792 8932 -3722
rect 8852 -3852 8862 -3792
rect 8922 -3852 8932 -3792
rect 9310 -3722 9320 -3672
rect 9776 -3662 9836 -3470
rect 9380 -3722 9390 -3672
rect 9310 -3792 9390 -3722
rect 9310 -3852 9320 -3792
rect 9380 -3852 9390 -3792
rect 9766 -3722 9776 -3672
rect 10232 -3662 10292 -3470
rect 9836 -3722 9846 -3672
rect 9766 -3792 9846 -3722
rect 9766 -3852 9776 -3792
rect 9836 -3852 9846 -3792
rect 10222 -3722 10232 -3672
rect 10690 -3662 10750 -3470
rect 10292 -3722 10302 -3672
rect 10222 -3792 10302 -3722
rect 10222 -3852 10232 -3792
rect 10292 -3852 10302 -3792
rect 10680 -3722 10690 -3672
rect 11146 -3662 11206 -3470
rect 10750 -3722 10760 -3672
rect 10680 -3792 10760 -3722
rect 10680 -3852 10690 -3792
rect 10750 -3852 10760 -3792
rect 11136 -3722 11146 -3672
rect 11602 -3662 11662 -3470
rect 11206 -3722 11216 -3672
rect 11136 -3792 11216 -3722
rect 11136 -3852 11146 -3792
rect 11206 -3852 11216 -3792
rect 11592 -3722 11602 -3672
rect 12060 -3662 12120 -3470
rect 11662 -3722 11672 -3672
rect 11592 -3792 11672 -3722
rect 11592 -3852 11602 -3792
rect 11662 -3852 11672 -3792
rect 12050 -3722 12060 -3672
rect 12516 -3662 12576 -3470
rect 12120 -3722 12130 -3672
rect 12050 -3792 12130 -3722
rect 12050 -3852 12060 -3792
rect 12120 -3852 12130 -3792
rect 12506 -3722 12516 -3672
rect 12972 -3662 13032 -3470
rect 12576 -3722 12586 -3672
rect 12506 -3792 12586 -3722
rect 12506 -3852 12516 -3792
rect 12576 -3852 12586 -3792
rect 12962 -3722 12972 -3672
rect 13430 -3662 13490 -3470
rect 13032 -3722 13042 -3672
rect 12962 -3792 13042 -3722
rect 12962 -3852 12972 -3792
rect 13032 -3852 13042 -3792
rect 13420 -3722 13430 -3672
rect 13886 -3662 13946 -3470
rect 13490 -3722 13500 -3672
rect 13420 -3792 13500 -3722
rect 13420 -3852 13430 -3792
rect 13490 -3852 13500 -3792
rect 13876 -3722 13886 -3672
rect 14342 -3662 14402 -3470
rect 13946 -3722 13956 -3672
rect 13876 -3792 13956 -3722
rect 13876 -3852 13886 -3792
rect 13946 -3852 13956 -3792
rect 14332 -3722 14342 -3672
rect 14800 -3662 14860 -3470
rect 14402 -3722 14412 -3672
rect 14332 -3792 14412 -3722
rect 14332 -3852 14342 -3792
rect 14402 -3852 14412 -3792
rect 14790 -3722 14800 -3672
rect 15256 -3662 15316 -3470
rect 14860 -3722 14870 -3672
rect 14790 -3792 14870 -3722
rect 14790 -3852 14800 -3792
rect 14860 -3852 14870 -3792
rect 15246 -3722 15256 -3672
rect 15316 -3722 15326 -3672
rect 15246 -3792 15326 -3722
rect 15246 -3852 15256 -3792
rect 15316 -3852 15326 -3792
rect 170 -4154 230 -3852
rect 160 -4214 170 -4164
rect 626 -4154 686 -3852
rect 230 -4214 240 -4164
rect 160 -4284 240 -4214
rect 160 -4344 170 -4284
rect 230 -4344 240 -4284
rect 616 -4214 626 -4164
rect 1082 -4154 1142 -3852
rect 686 -4214 696 -4164
rect 616 -4284 696 -4214
rect 616 -4344 626 -4284
rect 686 -4344 696 -4284
rect 1072 -4214 1082 -4164
rect 1540 -4154 1600 -3852
rect 1142 -4214 1152 -4164
rect 1072 -4284 1152 -4214
rect 1072 -4344 1082 -4284
rect 1142 -4344 1152 -4284
rect 1530 -4214 1540 -4164
rect 1996 -4154 2056 -3852
rect 1600 -4214 1610 -4164
rect 1530 -4284 1610 -4214
rect 1530 -4344 1540 -4284
rect 1600 -4344 1610 -4284
rect 1986 -4214 1996 -4164
rect 2452 -4154 2512 -3852
rect 2056 -4214 2066 -4164
rect 1986 -4284 2066 -4214
rect 1986 -4344 1996 -4284
rect 2056 -4344 2066 -4284
rect 2442 -4214 2452 -4164
rect 2910 -4154 2970 -3852
rect 2512 -4214 2522 -4164
rect 2442 -4284 2522 -4214
rect 2442 -4344 2452 -4284
rect 2512 -4344 2522 -4284
rect 2900 -4214 2910 -4164
rect 3366 -4154 3426 -3852
rect 2970 -4214 2980 -4164
rect 2900 -4284 2980 -4214
rect 2900 -4344 2910 -4284
rect 2970 -4344 2980 -4284
rect 3356 -4214 3366 -4164
rect 3822 -4154 3882 -3852
rect 3426 -4214 3436 -4164
rect 3356 -4284 3436 -4214
rect 3356 -4344 3366 -4284
rect 3426 -4344 3436 -4284
rect 3812 -4214 3822 -4164
rect 4280 -4154 4340 -3852
rect 3882 -4214 3892 -4164
rect 3812 -4284 3892 -4214
rect 3812 -4344 3822 -4284
rect 3882 -4344 3892 -4284
rect 4270 -4214 4280 -4164
rect 4736 -4154 4796 -3852
rect 4340 -4214 4350 -4164
rect 4270 -4284 4350 -4214
rect 4270 -4344 4280 -4284
rect 4340 -4344 4350 -4284
rect 4726 -4214 4736 -4164
rect 5192 -4154 5252 -3852
rect 4796 -4214 4806 -4164
rect 4726 -4284 4806 -4214
rect 4726 -4344 4736 -4284
rect 4796 -4344 4806 -4284
rect 5182 -4214 5192 -4164
rect 5650 -4154 5710 -3852
rect 5252 -4214 5262 -4164
rect 5182 -4284 5262 -4214
rect 5182 -4344 5192 -4284
rect 5252 -4344 5262 -4284
rect 5640 -4214 5650 -4164
rect 6106 -4154 6166 -3852
rect 5710 -4214 5720 -4164
rect 5640 -4284 5720 -4214
rect 5640 -4344 5650 -4284
rect 5710 -4344 5720 -4284
rect 6096 -4214 6106 -4164
rect 6562 -4154 6622 -3852
rect 6166 -4214 6176 -4164
rect 6096 -4284 6176 -4214
rect 6096 -4344 6106 -4284
rect 6166 -4344 6176 -4284
rect 6552 -4214 6562 -4164
rect 7020 -4154 7080 -3852
rect 6622 -4214 6632 -4164
rect 6552 -4284 6632 -4214
rect 6552 -4344 6562 -4284
rect 6622 -4344 6632 -4284
rect 7010 -4214 7020 -4164
rect 7476 -4154 7536 -3852
rect 7080 -4214 7090 -4164
rect 7010 -4284 7090 -4214
rect 7010 -4344 7020 -4284
rect 7080 -4344 7090 -4284
rect 7466 -4214 7476 -4164
rect 7932 -4154 7992 -3852
rect 7536 -4214 7546 -4164
rect 7466 -4284 7546 -4214
rect 7466 -4344 7476 -4284
rect 7536 -4344 7546 -4284
rect 7922 -4214 7932 -4164
rect 8406 -4154 8466 -3852
rect 7992 -4214 8002 -4164
rect 7922 -4284 8002 -4214
rect 7922 -4344 7932 -4284
rect 7992 -4344 8002 -4284
rect 8396 -4214 8406 -4164
rect 8862 -4154 8922 -3852
rect 8466 -4214 8476 -4164
rect 8396 -4284 8476 -4214
rect 8396 -4344 8406 -4284
rect 8466 -4344 8476 -4284
rect 8852 -4214 8862 -4164
rect 9320 -4154 9380 -3852
rect 8922 -4214 8932 -4164
rect 8852 -4284 8932 -4214
rect 8852 -4344 8862 -4284
rect 8922 -4344 8932 -4284
rect 9310 -4214 9320 -4164
rect 9776 -4154 9836 -3852
rect 9380 -4214 9390 -4164
rect 9310 -4284 9390 -4214
rect 9310 -4344 9320 -4284
rect 9380 -4344 9390 -4284
rect 9766 -4214 9776 -4164
rect 10232 -4154 10292 -3852
rect 9836 -4214 9846 -4164
rect 9766 -4284 9846 -4214
rect 9766 -4344 9776 -4284
rect 9836 -4344 9846 -4284
rect 10222 -4214 10232 -4164
rect 10690 -4154 10750 -3852
rect 10292 -4214 10302 -4164
rect 10222 -4284 10302 -4214
rect 10222 -4344 10232 -4284
rect 10292 -4344 10302 -4284
rect 10680 -4214 10690 -4164
rect 11146 -4154 11206 -3852
rect 10750 -4214 10760 -4164
rect 10680 -4284 10760 -4214
rect 10680 -4344 10690 -4284
rect 10750 -4344 10760 -4284
rect 11136 -4214 11146 -4164
rect 11602 -4154 11662 -3852
rect 11206 -4214 11216 -4164
rect 11136 -4284 11216 -4214
rect 11136 -4344 11146 -4284
rect 11206 -4344 11216 -4284
rect 11592 -4214 11602 -4164
rect 12060 -4154 12120 -3852
rect 11662 -4214 11672 -4164
rect 11592 -4284 11672 -4214
rect 11592 -4344 11602 -4284
rect 11662 -4344 11672 -4284
rect 12050 -4214 12060 -4164
rect 12516 -4154 12576 -3852
rect 12120 -4214 12130 -4164
rect 12050 -4284 12130 -4214
rect 12050 -4344 12060 -4284
rect 12120 -4344 12130 -4284
rect 12506 -4214 12516 -4164
rect 12972 -4154 13032 -3852
rect 12576 -4214 12586 -4164
rect 12506 -4284 12586 -4214
rect 12506 -4344 12516 -4284
rect 12576 -4344 12586 -4284
rect 12962 -4214 12972 -4164
rect 13430 -4154 13490 -3852
rect 13032 -4214 13042 -4164
rect 12962 -4284 13042 -4214
rect 12962 -4344 12972 -4284
rect 13032 -4344 13042 -4284
rect 13420 -4214 13430 -4164
rect 13886 -4154 13946 -3852
rect 13490 -4214 13500 -4164
rect 13420 -4284 13500 -4214
rect 13420 -4344 13430 -4284
rect 13490 -4344 13500 -4284
rect 13876 -4214 13886 -4164
rect 14342 -4154 14402 -3852
rect 13946 -4214 13956 -4164
rect 13876 -4284 13956 -4214
rect 13876 -4344 13886 -4284
rect 13946 -4344 13956 -4284
rect 14332 -4214 14342 -4164
rect 14800 -4154 14860 -3852
rect 14402 -4214 14412 -4164
rect 14332 -4284 14412 -4214
rect 14332 -4344 14342 -4284
rect 14402 -4344 14412 -4284
rect 14790 -4214 14800 -4164
rect 15256 -4154 15316 -3852
rect 14860 -4214 14870 -4164
rect 14790 -4284 14870 -4214
rect 14790 -4344 14800 -4284
rect 14860 -4344 14870 -4284
rect 15246 -4214 15256 -4164
rect 15316 -4214 15326 -4164
rect 15246 -4284 15326 -4214
rect 15246 -4344 15256 -4284
rect 15316 -4344 15326 -4284
rect 170 -4670 230 -4344
rect 160 -4730 170 -4680
rect 626 -4670 686 -4344
rect 230 -4730 240 -4680
rect 160 -4800 240 -4730
rect 160 -4860 170 -4800
rect 230 -4860 240 -4800
rect 616 -4730 626 -4680
rect 1082 -4670 1142 -4344
rect 686 -4730 696 -4680
rect 616 -4800 696 -4730
rect 616 -4860 626 -4800
rect 686 -4860 696 -4800
rect 1072 -4730 1082 -4680
rect 1540 -4670 1600 -4344
rect 1142 -4730 1152 -4680
rect 1072 -4800 1152 -4730
rect 1072 -4860 1082 -4800
rect 1142 -4860 1152 -4800
rect 1530 -4730 1540 -4680
rect 1996 -4670 2056 -4344
rect 1600 -4730 1610 -4680
rect 1530 -4800 1610 -4730
rect 1530 -4860 1540 -4800
rect 1600 -4860 1610 -4800
rect 1986 -4730 1996 -4680
rect 2452 -4670 2512 -4344
rect 2056 -4730 2066 -4680
rect 1986 -4800 2066 -4730
rect 1986 -4860 1996 -4800
rect 2056 -4860 2066 -4800
rect 2442 -4730 2452 -4680
rect 2910 -4670 2970 -4344
rect 2512 -4730 2522 -4680
rect 2442 -4800 2522 -4730
rect 2442 -4860 2452 -4800
rect 2512 -4860 2522 -4800
rect 2900 -4730 2910 -4680
rect 3366 -4670 3426 -4344
rect 2970 -4730 2980 -4680
rect 2900 -4800 2980 -4730
rect 2900 -4860 2910 -4800
rect 2970 -4860 2980 -4800
rect 3356 -4730 3366 -4680
rect 3822 -4670 3882 -4344
rect 3426 -4730 3436 -4680
rect 3356 -4800 3436 -4730
rect 3356 -4860 3366 -4800
rect 3426 -4860 3436 -4800
rect 3812 -4730 3822 -4680
rect 4280 -4670 4340 -4344
rect 3882 -4730 3892 -4680
rect 3812 -4800 3892 -4730
rect 3812 -4860 3822 -4800
rect 3882 -4860 3892 -4800
rect 4270 -4730 4280 -4680
rect 4736 -4670 4796 -4344
rect 4340 -4730 4350 -4680
rect 4270 -4800 4350 -4730
rect 4270 -4860 4280 -4800
rect 4340 -4860 4350 -4800
rect 4726 -4730 4736 -4680
rect 5192 -4670 5252 -4344
rect 4796 -4730 4806 -4680
rect 4726 -4800 4806 -4730
rect 4726 -4860 4736 -4800
rect 4796 -4860 4806 -4800
rect 5182 -4730 5192 -4680
rect 5650 -4670 5710 -4344
rect 5252 -4730 5262 -4680
rect 5182 -4800 5262 -4730
rect 5182 -4860 5192 -4800
rect 5252 -4860 5262 -4800
rect 5640 -4730 5650 -4680
rect 6106 -4670 6166 -4344
rect 5710 -4730 5720 -4680
rect 5640 -4800 5720 -4730
rect 5640 -4860 5650 -4800
rect 5710 -4860 5720 -4800
rect 6096 -4730 6106 -4680
rect 6562 -4670 6622 -4344
rect 6166 -4730 6176 -4680
rect 6096 -4800 6176 -4730
rect 6096 -4860 6106 -4800
rect 6166 -4860 6176 -4800
rect 6552 -4730 6562 -4680
rect 7020 -4670 7080 -4344
rect 6622 -4730 6632 -4680
rect 6552 -4800 6632 -4730
rect 6552 -4860 6562 -4800
rect 6622 -4860 6632 -4800
rect 7010 -4730 7020 -4680
rect 7476 -4670 7536 -4344
rect 7080 -4730 7090 -4680
rect 7010 -4800 7090 -4730
rect 7010 -4860 7020 -4800
rect 7080 -4860 7090 -4800
rect 7466 -4730 7476 -4680
rect 7932 -4670 7992 -4344
rect 7536 -4730 7546 -4680
rect 7466 -4800 7546 -4730
rect 7466 -4860 7476 -4800
rect 7536 -4860 7546 -4800
rect 7922 -4730 7932 -4680
rect 8406 -4670 8466 -4344
rect 7992 -4730 8002 -4680
rect 7922 -4800 8002 -4730
rect 7922 -4860 7932 -4800
rect 7992 -4860 8002 -4800
rect 8396 -4730 8406 -4680
rect 8862 -4670 8922 -4344
rect 8466 -4730 8476 -4680
rect 8396 -4800 8476 -4730
rect 8396 -4860 8406 -4800
rect 8466 -4860 8476 -4800
rect 8852 -4730 8862 -4680
rect 9320 -4670 9380 -4344
rect 8922 -4730 8932 -4680
rect 8852 -4800 8932 -4730
rect 8852 -4860 8862 -4800
rect 8922 -4860 8932 -4800
rect 9310 -4730 9320 -4680
rect 9776 -4670 9836 -4344
rect 9380 -4730 9390 -4680
rect 9310 -4800 9390 -4730
rect 9310 -4860 9320 -4800
rect 9380 -4860 9390 -4800
rect 9766 -4730 9776 -4680
rect 10232 -4670 10292 -4344
rect 9836 -4730 9846 -4680
rect 9766 -4800 9846 -4730
rect 9766 -4860 9776 -4800
rect 9836 -4860 9846 -4800
rect 10222 -4730 10232 -4680
rect 10690 -4670 10750 -4344
rect 10292 -4730 10302 -4680
rect 10222 -4800 10302 -4730
rect 10222 -4860 10232 -4800
rect 10292 -4860 10302 -4800
rect 10680 -4730 10690 -4680
rect 11146 -4670 11206 -4344
rect 10750 -4730 10760 -4680
rect 10680 -4800 10760 -4730
rect 10680 -4860 10690 -4800
rect 10750 -4860 10760 -4800
rect 11136 -4730 11146 -4680
rect 11602 -4670 11662 -4344
rect 11206 -4730 11216 -4680
rect 11136 -4800 11216 -4730
rect 11136 -4860 11146 -4800
rect 11206 -4860 11216 -4800
rect 11592 -4730 11602 -4680
rect 12060 -4670 12120 -4344
rect 11662 -4730 11672 -4680
rect 11592 -4800 11672 -4730
rect 11592 -4860 11602 -4800
rect 11662 -4860 11672 -4800
rect 12050 -4730 12060 -4680
rect 12516 -4670 12576 -4344
rect 12120 -4730 12130 -4680
rect 12050 -4800 12130 -4730
rect 12050 -4860 12060 -4800
rect 12120 -4860 12130 -4800
rect 12506 -4730 12516 -4680
rect 12972 -4670 13032 -4344
rect 12576 -4730 12586 -4680
rect 12506 -4800 12586 -4730
rect 12506 -4860 12516 -4800
rect 12576 -4860 12586 -4800
rect 12962 -4730 12972 -4680
rect 13430 -4670 13490 -4344
rect 13032 -4730 13042 -4680
rect 12962 -4800 13042 -4730
rect 12962 -4860 12972 -4800
rect 13032 -4860 13042 -4800
rect 13420 -4730 13430 -4680
rect 13886 -4670 13946 -4344
rect 13490 -4730 13500 -4680
rect 13420 -4800 13500 -4730
rect 13420 -4860 13430 -4800
rect 13490 -4860 13500 -4800
rect 13876 -4730 13886 -4680
rect 14342 -4670 14402 -4344
rect 13946 -4730 13956 -4680
rect 13876 -4800 13956 -4730
rect 13876 -4860 13886 -4800
rect 13946 -4860 13956 -4800
rect 14332 -4730 14342 -4680
rect 14800 -4670 14860 -4344
rect 14402 -4730 14412 -4680
rect 14332 -4800 14412 -4730
rect 14332 -4860 14342 -4800
rect 14402 -4860 14412 -4800
rect 14790 -4730 14800 -4680
rect 15256 -4670 15316 -4344
rect 14860 -4730 14870 -4680
rect 14790 -4800 14870 -4730
rect 14790 -4860 14800 -4800
rect 14860 -4860 14870 -4800
rect 15246 -4730 15256 -4680
rect 15316 -4730 15326 -4680
rect 15246 -4800 15326 -4730
rect 15246 -4860 15256 -4800
rect 15316 -4860 15326 -4800
rect 170 -5172 230 -4860
rect 160 -5232 170 -5182
rect 626 -5172 686 -4860
rect 230 -5232 240 -5182
rect 160 -5302 240 -5232
rect 160 -5362 170 -5302
rect 230 -5362 240 -5302
rect 616 -5232 626 -5182
rect 1082 -5172 1142 -4860
rect 686 -5232 696 -5182
rect 616 -5302 696 -5232
rect 616 -5362 626 -5302
rect 686 -5362 696 -5302
rect 1072 -5232 1082 -5182
rect 1540 -5172 1600 -4860
rect 1142 -5232 1152 -5182
rect 1072 -5302 1152 -5232
rect 1072 -5362 1082 -5302
rect 1142 -5362 1152 -5302
rect 1530 -5232 1540 -5182
rect 1996 -5172 2056 -4860
rect 1600 -5232 1610 -5182
rect 1530 -5302 1610 -5232
rect 1530 -5362 1540 -5302
rect 1600 -5362 1610 -5302
rect 1986 -5232 1996 -5182
rect 2452 -5172 2512 -4860
rect 2056 -5232 2066 -5182
rect 1986 -5302 2066 -5232
rect 1986 -5362 1996 -5302
rect 2056 -5362 2066 -5302
rect 2442 -5232 2452 -5182
rect 2910 -5172 2970 -4860
rect 2512 -5232 2522 -5182
rect 2442 -5302 2522 -5232
rect 2442 -5362 2452 -5302
rect 2512 -5362 2522 -5302
rect 2900 -5232 2910 -5182
rect 3366 -5172 3426 -4860
rect 2970 -5232 2980 -5182
rect 2900 -5302 2980 -5232
rect 2900 -5362 2910 -5302
rect 2970 -5362 2980 -5302
rect 3356 -5232 3366 -5182
rect 3822 -5172 3882 -4860
rect 3426 -5232 3436 -5182
rect 3356 -5302 3436 -5232
rect 3356 -5362 3366 -5302
rect 3426 -5362 3436 -5302
rect 3812 -5232 3822 -5182
rect 4280 -5172 4340 -4860
rect 3882 -5232 3892 -5182
rect 3812 -5302 3892 -5232
rect 3812 -5362 3822 -5302
rect 3882 -5362 3892 -5302
rect 4270 -5232 4280 -5182
rect 4736 -5172 4796 -4860
rect 4340 -5232 4350 -5182
rect 4270 -5302 4350 -5232
rect 4270 -5362 4280 -5302
rect 4340 -5362 4350 -5302
rect 4726 -5232 4736 -5182
rect 5192 -5172 5252 -4860
rect 4796 -5232 4806 -5182
rect 4726 -5302 4806 -5232
rect 4726 -5362 4736 -5302
rect 4796 -5362 4806 -5302
rect 5182 -5232 5192 -5182
rect 5650 -5172 5710 -4860
rect 5252 -5232 5262 -5182
rect 5182 -5302 5262 -5232
rect 5182 -5362 5192 -5302
rect 5252 -5362 5262 -5302
rect 5640 -5232 5650 -5182
rect 6106 -5172 6166 -4860
rect 5710 -5232 5720 -5182
rect 5640 -5302 5720 -5232
rect 5640 -5362 5650 -5302
rect 5710 -5362 5720 -5302
rect 6096 -5232 6106 -5182
rect 6562 -5172 6622 -4860
rect 6166 -5232 6176 -5182
rect 6096 -5302 6176 -5232
rect 6096 -5362 6106 -5302
rect 6166 -5362 6176 -5302
rect 6552 -5232 6562 -5182
rect 7020 -5172 7080 -4860
rect 6622 -5232 6632 -5182
rect 6552 -5302 6632 -5232
rect 6552 -5362 6562 -5302
rect 6622 -5362 6632 -5302
rect 7010 -5232 7020 -5182
rect 7476 -5172 7536 -4860
rect 7080 -5232 7090 -5182
rect 7010 -5302 7090 -5232
rect 7010 -5362 7020 -5302
rect 7080 -5362 7090 -5302
rect 7466 -5232 7476 -5182
rect 7932 -5172 7992 -4860
rect 7536 -5232 7546 -5182
rect 7466 -5302 7546 -5232
rect 7466 -5362 7476 -5302
rect 7536 -5362 7546 -5302
rect 7922 -5232 7932 -5182
rect 8406 -5172 8466 -4860
rect 7992 -5232 8002 -5182
rect 7922 -5302 8002 -5232
rect 7922 -5362 7932 -5302
rect 7992 -5362 8002 -5302
rect 8396 -5232 8406 -5182
rect 8862 -5172 8922 -4860
rect 8466 -5232 8476 -5182
rect 8396 -5302 8476 -5232
rect 8396 -5362 8406 -5302
rect 8466 -5362 8476 -5302
rect 8852 -5232 8862 -5182
rect 9320 -5172 9380 -4860
rect 8922 -5232 8932 -5182
rect 8852 -5302 8932 -5232
rect 8852 -5362 8862 -5302
rect 8922 -5362 8932 -5302
rect 9310 -5232 9320 -5182
rect 9776 -5172 9836 -4860
rect 9380 -5232 9390 -5182
rect 9310 -5302 9390 -5232
rect 9310 -5362 9320 -5302
rect 9380 -5362 9390 -5302
rect 9766 -5232 9776 -5182
rect 10232 -5172 10292 -4860
rect 9836 -5232 9846 -5182
rect 9766 -5302 9846 -5232
rect 9766 -5362 9776 -5302
rect 9836 -5362 9846 -5302
rect 10222 -5232 10232 -5182
rect 10690 -5172 10750 -4860
rect 10292 -5232 10302 -5182
rect 10222 -5302 10302 -5232
rect 10222 -5362 10232 -5302
rect 10292 -5362 10302 -5302
rect 10680 -5232 10690 -5182
rect 11146 -5172 11206 -4860
rect 10750 -5232 10760 -5182
rect 10680 -5302 10760 -5232
rect 10680 -5362 10690 -5302
rect 10750 -5362 10760 -5302
rect 11136 -5232 11146 -5182
rect 11602 -5172 11662 -4860
rect 11206 -5232 11216 -5182
rect 11136 -5302 11216 -5232
rect 11136 -5362 11146 -5302
rect 11206 -5362 11216 -5302
rect 11592 -5232 11602 -5182
rect 12060 -5172 12120 -4860
rect 11662 -5232 11672 -5182
rect 11592 -5302 11672 -5232
rect 11592 -5362 11602 -5302
rect 11662 -5362 11672 -5302
rect 12050 -5232 12060 -5182
rect 12516 -5172 12576 -4860
rect 12120 -5232 12130 -5182
rect 12050 -5302 12130 -5232
rect 12050 -5362 12060 -5302
rect 12120 -5362 12130 -5302
rect 12506 -5232 12516 -5182
rect 12972 -5172 13032 -4860
rect 12576 -5232 12586 -5182
rect 12506 -5302 12586 -5232
rect 12506 -5362 12516 -5302
rect 12576 -5362 12586 -5302
rect 12962 -5232 12972 -5182
rect 13430 -5172 13490 -4860
rect 13032 -5232 13042 -5182
rect 12962 -5302 13042 -5232
rect 12962 -5362 12972 -5302
rect 13032 -5362 13042 -5302
rect 13420 -5232 13430 -5182
rect 13886 -5172 13946 -4860
rect 13490 -5232 13500 -5182
rect 13420 -5302 13500 -5232
rect 13420 -5362 13430 -5302
rect 13490 -5362 13500 -5302
rect 13876 -5232 13886 -5182
rect 14342 -5172 14402 -4860
rect 13946 -5232 13956 -5182
rect 13876 -5302 13956 -5232
rect 13876 -5362 13886 -5302
rect 13946 -5362 13956 -5302
rect 14332 -5232 14342 -5182
rect 14800 -5172 14860 -4860
rect 14402 -5232 14412 -5182
rect 14332 -5302 14412 -5232
rect 14332 -5362 14342 -5302
rect 14402 -5362 14412 -5302
rect 14790 -5232 14800 -5182
rect 15256 -5172 15316 -4860
rect 14860 -5232 14870 -5182
rect 14790 -5302 14870 -5232
rect 14790 -5362 14800 -5302
rect 14860 -5362 14870 -5302
rect 15246 -5232 15256 -5182
rect 15316 -5232 15326 -5182
rect 15246 -5302 15326 -5232
rect 15246 -5362 15256 -5302
rect 15316 -5362 15326 -5302
rect 170 -5664 230 -5362
rect 160 -5724 170 -5674
rect 626 -5664 686 -5362
rect 230 -5724 240 -5674
rect 160 -5794 240 -5724
rect 160 -5854 170 -5794
rect 230 -5854 240 -5794
rect 616 -5724 626 -5674
rect 1082 -5664 1142 -5362
rect 686 -5724 696 -5674
rect 616 -5794 696 -5724
rect 616 -5854 626 -5794
rect 686 -5854 696 -5794
rect 1072 -5724 1082 -5674
rect 1540 -5664 1600 -5362
rect 1142 -5724 1152 -5674
rect 1072 -5794 1152 -5724
rect 1072 -5854 1082 -5794
rect 1142 -5854 1152 -5794
rect 1530 -5724 1540 -5674
rect 1996 -5664 2056 -5362
rect 1600 -5724 1610 -5674
rect 1530 -5794 1610 -5724
rect 1530 -5854 1540 -5794
rect 1600 -5854 1610 -5794
rect 1986 -5724 1996 -5674
rect 2452 -5664 2512 -5362
rect 2056 -5724 2066 -5674
rect 1986 -5794 2066 -5724
rect 1986 -5854 1996 -5794
rect 2056 -5854 2066 -5794
rect 2442 -5724 2452 -5674
rect 2910 -5664 2970 -5362
rect 2512 -5724 2522 -5674
rect 2442 -5794 2522 -5724
rect 2442 -5854 2452 -5794
rect 2512 -5854 2522 -5794
rect 2900 -5724 2910 -5674
rect 3366 -5664 3426 -5362
rect 2970 -5724 2980 -5674
rect 2900 -5794 2980 -5724
rect 2900 -5854 2910 -5794
rect 2970 -5854 2980 -5794
rect 3356 -5724 3366 -5674
rect 3822 -5664 3882 -5362
rect 3426 -5724 3436 -5674
rect 3356 -5794 3436 -5724
rect 3356 -5854 3366 -5794
rect 3426 -5854 3436 -5794
rect 3812 -5724 3822 -5674
rect 4280 -5664 4340 -5362
rect 3882 -5724 3892 -5674
rect 3812 -5794 3892 -5724
rect 3812 -5854 3822 -5794
rect 3882 -5854 3892 -5794
rect 4270 -5724 4280 -5674
rect 4736 -5664 4796 -5362
rect 4340 -5724 4350 -5674
rect 4270 -5794 4350 -5724
rect 4270 -5854 4280 -5794
rect 4340 -5854 4350 -5794
rect 4726 -5724 4736 -5674
rect 5192 -5664 5252 -5362
rect 4796 -5724 4806 -5674
rect 4726 -5794 4806 -5724
rect 4726 -5854 4736 -5794
rect 4796 -5854 4806 -5794
rect 5182 -5724 5192 -5674
rect 5650 -5664 5710 -5362
rect 5252 -5724 5262 -5674
rect 5182 -5794 5262 -5724
rect 5182 -5854 5192 -5794
rect 5252 -5854 5262 -5794
rect 5640 -5724 5650 -5674
rect 6106 -5664 6166 -5362
rect 5710 -5724 5720 -5674
rect 5640 -5794 5720 -5724
rect 5640 -5854 5650 -5794
rect 5710 -5854 5720 -5794
rect 6096 -5724 6106 -5674
rect 6562 -5664 6622 -5362
rect 6166 -5724 6176 -5674
rect 6096 -5794 6176 -5724
rect 6096 -5854 6106 -5794
rect 6166 -5854 6176 -5794
rect 6552 -5724 6562 -5674
rect 7020 -5664 7080 -5362
rect 6622 -5724 6632 -5674
rect 6552 -5794 6632 -5724
rect 6552 -5854 6562 -5794
rect 6622 -5854 6632 -5794
rect 7010 -5724 7020 -5674
rect 7476 -5664 7536 -5362
rect 7080 -5724 7090 -5674
rect 7010 -5794 7090 -5724
rect 7010 -5854 7020 -5794
rect 7080 -5854 7090 -5794
rect 7466 -5724 7476 -5674
rect 7932 -5664 7992 -5362
rect 7536 -5724 7546 -5674
rect 7466 -5794 7546 -5724
rect 7466 -5854 7476 -5794
rect 7536 -5854 7546 -5794
rect 7922 -5724 7932 -5674
rect 8406 -5664 8466 -5362
rect 7992 -5724 8002 -5674
rect 7922 -5794 8002 -5724
rect 7922 -5854 7932 -5794
rect 7992 -5854 8002 -5794
rect 8396 -5724 8406 -5674
rect 8862 -5664 8922 -5362
rect 8466 -5724 8476 -5674
rect 8396 -5794 8476 -5724
rect 8396 -5854 8406 -5794
rect 8466 -5854 8476 -5794
rect 8852 -5724 8862 -5674
rect 9320 -5664 9380 -5362
rect 8922 -5724 8932 -5674
rect 8852 -5794 8932 -5724
rect 8852 -5854 8862 -5794
rect 8922 -5854 8932 -5794
rect 9310 -5724 9320 -5674
rect 9776 -5664 9836 -5362
rect 9380 -5724 9390 -5674
rect 9310 -5794 9390 -5724
rect 9310 -5854 9320 -5794
rect 9380 -5854 9390 -5794
rect 9766 -5724 9776 -5674
rect 10232 -5664 10292 -5362
rect 9836 -5724 9846 -5674
rect 9766 -5794 9846 -5724
rect 9766 -5854 9776 -5794
rect 9836 -5854 9846 -5794
rect 10222 -5724 10232 -5674
rect 10690 -5664 10750 -5362
rect 10292 -5724 10302 -5674
rect 10222 -5794 10302 -5724
rect 10222 -5854 10232 -5794
rect 10292 -5854 10302 -5794
rect 10680 -5724 10690 -5674
rect 11146 -5664 11206 -5362
rect 10750 -5724 10760 -5674
rect 10680 -5794 10760 -5724
rect 10680 -5854 10690 -5794
rect 10750 -5854 10760 -5794
rect 11136 -5724 11146 -5674
rect 11602 -5664 11662 -5362
rect 11206 -5724 11216 -5674
rect 11136 -5794 11216 -5724
rect 11136 -5854 11146 -5794
rect 11206 -5854 11216 -5794
rect 11592 -5724 11602 -5674
rect 12060 -5664 12120 -5362
rect 11662 -5724 11672 -5674
rect 11592 -5794 11672 -5724
rect 11592 -5854 11602 -5794
rect 11662 -5854 11672 -5794
rect 12050 -5724 12060 -5674
rect 12516 -5664 12576 -5362
rect 12120 -5724 12130 -5674
rect 12050 -5794 12130 -5724
rect 12050 -5854 12060 -5794
rect 12120 -5854 12130 -5794
rect 12506 -5724 12516 -5674
rect 12972 -5664 13032 -5362
rect 12576 -5724 12586 -5674
rect 12506 -5794 12586 -5724
rect 12506 -5854 12516 -5794
rect 12576 -5854 12586 -5794
rect 12962 -5724 12972 -5674
rect 13430 -5664 13490 -5362
rect 13032 -5724 13042 -5674
rect 12962 -5794 13042 -5724
rect 12962 -5854 12972 -5794
rect 13032 -5854 13042 -5794
rect 13420 -5724 13430 -5674
rect 13886 -5664 13946 -5362
rect 13490 -5724 13500 -5674
rect 13420 -5794 13500 -5724
rect 13420 -5854 13430 -5794
rect 13490 -5854 13500 -5794
rect 13876 -5724 13886 -5674
rect 14342 -5664 14402 -5362
rect 13946 -5724 13956 -5674
rect 13876 -5794 13956 -5724
rect 13876 -5854 13886 -5794
rect 13946 -5854 13956 -5794
rect 14332 -5724 14342 -5674
rect 14800 -5664 14860 -5362
rect 14402 -5724 14412 -5674
rect 14332 -5794 14412 -5724
rect 14332 -5854 14342 -5794
rect 14402 -5854 14412 -5794
rect 14790 -5724 14800 -5674
rect 15256 -5664 15316 -5362
rect 14860 -5724 14870 -5674
rect 14790 -5794 14870 -5724
rect 14790 -5854 14800 -5794
rect 14860 -5854 14870 -5794
rect 15246 -5724 15256 -5674
rect 15316 -5724 15326 -5674
rect 15246 -5794 15326 -5724
rect 15246 -5854 15256 -5794
rect 15316 -5854 15326 -5794
rect 170 -5990 230 -5854
rect 626 -5990 686 -5854
rect 1082 -5990 1142 -5854
rect 1540 -5990 1600 -5854
rect 1996 -5990 2056 -5854
rect 2452 -5990 2512 -5854
rect 2910 -5990 2970 -5854
rect 3366 -5990 3426 -5854
rect 3822 -5990 3882 -5854
rect 4280 -5990 4340 -5854
rect 4736 -5990 4796 -5854
rect 5192 -5990 5252 -5854
rect 5650 -5990 5710 -5854
rect 6106 -5990 6166 -5854
rect 6562 -5990 6622 -5854
rect 7020 -5990 7080 -5854
rect 7476 -5990 7536 -5854
rect 7932 -5990 7992 -5854
rect 8406 -5990 8466 -5854
rect 8862 -5990 8922 -5854
rect 9320 -5990 9380 -5854
rect 9776 -5990 9836 -5854
rect 10232 -5990 10292 -5854
rect 10690 -5990 10750 -5854
rect 11146 -5990 11206 -5854
rect 11602 -5990 11662 -5854
rect 12060 -5990 12120 -5854
rect 12516 -5990 12576 -5854
rect 12972 -5990 13032 -5854
rect 13430 -5990 13490 -5854
rect 13886 -5990 13946 -5854
rect 14342 -5990 14402 -5854
rect 14800 -5990 14860 -5854
rect 15256 -5990 15316 -5854
rect 170 -5994 231 -5990
rect 626 -5994 687 -5990
rect 1082 -5994 1143 -5990
rect 1540 -5994 1601 -5990
rect 1996 -5994 2057 -5990
rect 2452 -5994 2513 -5990
rect 2910 -5994 2971 -5990
rect 3366 -5994 3427 -5990
rect 3822 -5994 3883 -5990
rect 4280 -5994 4341 -5990
rect 4736 -5994 4797 -5990
rect 5192 -5994 5253 -5990
rect 5650 -5994 5711 -5990
rect 6106 -5994 6167 -5990
rect 6562 -5994 6623 -5990
rect 7020 -5994 7081 -5990
rect 7476 -5994 7537 -5990
rect 7932 -5994 7993 -5990
rect 8406 -5994 8467 -5990
rect 8862 -5994 8923 -5990
rect 9320 -5994 9381 -5990
rect 9776 -5994 9837 -5990
rect 10232 -5994 10293 -5990
rect 10690 -5994 10751 -5990
rect 11146 -5994 11207 -5990
rect 11602 -5994 11663 -5990
rect 12060 -5994 12121 -5990
rect 12516 -5994 12577 -5990
rect 12972 -5994 13033 -5990
rect 13430 -5994 13491 -5990
rect 13886 -5994 13947 -5990
rect 14342 -5994 14403 -5990
rect 14800 -5994 14861 -5990
rect 15256 -5994 15317 -5990
rect 171 -6161 231 -5994
rect 161 -6221 171 -6171
rect 627 -6161 687 -5994
rect 231 -6221 241 -6171
rect 161 -6291 241 -6221
rect 161 -6351 171 -6291
rect 231 -6351 241 -6291
rect 617 -6221 627 -6171
rect 1083 -6161 1143 -5994
rect 687 -6221 697 -6171
rect 617 -6291 697 -6221
rect 617 -6351 627 -6291
rect 687 -6351 697 -6291
rect 1073 -6221 1083 -6171
rect 1541 -6161 1601 -5994
rect 1143 -6221 1153 -6171
rect 1073 -6291 1153 -6221
rect 1073 -6351 1083 -6291
rect 1143 -6351 1153 -6291
rect 1531 -6221 1541 -6171
rect 1997 -6161 2057 -5994
rect 1601 -6221 1611 -6171
rect 1531 -6291 1611 -6221
rect 1531 -6351 1541 -6291
rect 1601 -6351 1611 -6291
rect 1987 -6221 1997 -6171
rect 2453 -6161 2513 -5994
rect 2057 -6221 2067 -6171
rect 1987 -6291 2067 -6221
rect 1987 -6351 1997 -6291
rect 2057 -6351 2067 -6291
rect 2443 -6221 2453 -6171
rect 2911 -6161 2971 -5994
rect 2513 -6221 2523 -6171
rect 2443 -6291 2523 -6221
rect 2443 -6351 2453 -6291
rect 2513 -6351 2523 -6291
rect 2901 -6221 2911 -6171
rect 3367 -6161 3427 -5994
rect 2971 -6221 2981 -6171
rect 2901 -6291 2981 -6221
rect 2901 -6351 2911 -6291
rect 2971 -6351 2981 -6291
rect 3357 -6221 3367 -6171
rect 3823 -6161 3883 -5994
rect 3427 -6221 3437 -6171
rect 3357 -6291 3437 -6221
rect 3357 -6351 3367 -6291
rect 3427 -6351 3437 -6291
rect 3813 -6221 3823 -6171
rect 4281 -6161 4341 -5994
rect 3883 -6221 3893 -6171
rect 3813 -6291 3893 -6221
rect 3813 -6351 3823 -6291
rect 3883 -6351 3893 -6291
rect 4271 -6221 4281 -6171
rect 4737 -6161 4797 -5994
rect 4341 -6221 4351 -6171
rect 4271 -6291 4351 -6221
rect 4271 -6351 4281 -6291
rect 4341 -6351 4351 -6291
rect 4727 -6221 4737 -6171
rect 5193 -6161 5253 -5994
rect 4797 -6221 4807 -6171
rect 4727 -6291 4807 -6221
rect 4727 -6351 4737 -6291
rect 4797 -6351 4807 -6291
rect 5183 -6221 5193 -6171
rect 5651 -6161 5711 -5994
rect 5253 -6221 5263 -6171
rect 5183 -6291 5263 -6221
rect 5183 -6351 5193 -6291
rect 5253 -6351 5263 -6291
rect 5641 -6221 5651 -6171
rect 6107 -6161 6167 -5994
rect 5711 -6221 5721 -6171
rect 5641 -6291 5721 -6221
rect 5641 -6351 5651 -6291
rect 5711 -6351 5721 -6291
rect 6097 -6221 6107 -6171
rect 6563 -6161 6623 -5994
rect 6167 -6221 6177 -6171
rect 6097 -6291 6177 -6221
rect 6097 -6351 6107 -6291
rect 6167 -6351 6177 -6291
rect 6553 -6221 6563 -6171
rect 7021 -6161 7081 -5994
rect 6623 -6221 6633 -6171
rect 6553 -6291 6633 -6221
rect 6553 -6351 6563 -6291
rect 6623 -6351 6633 -6291
rect 7011 -6221 7021 -6171
rect 7477 -6161 7537 -5994
rect 7081 -6221 7091 -6171
rect 7011 -6291 7091 -6221
rect 7011 -6351 7021 -6291
rect 7081 -6351 7091 -6291
rect 7467 -6221 7477 -6171
rect 7933 -6161 7993 -5994
rect 7537 -6221 7547 -6171
rect 7467 -6291 7547 -6221
rect 7467 -6351 7477 -6291
rect 7537 -6351 7547 -6291
rect 7923 -6221 7933 -6171
rect 8407 -6161 8467 -5994
rect 7993 -6221 8003 -6171
rect 7923 -6291 8003 -6221
rect 7923 -6351 7933 -6291
rect 7993 -6351 8003 -6291
rect 8397 -6221 8407 -6171
rect 8863 -6161 8923 -5994
rect 8467 -6221 8477 -6171
rect 8397 -6291 8477 -6221
rect 8397 -6351 8407 -6291
rect 8467 -6351 8477 -6291
rect 8853 -6221 8863 -6171
rect 9321 -6161 9381 -5994
rect 8923 -6221 8933 -6171
rect 8853 -6291 8933 -6221
rect 8853 -6351 8863 -6291
rect 8923 -6351 8933 -6291
rect 9311 -6221 9321 -6171
rect 9777 -6161 9837 -5994
rect 9381 -6221 9391 -6171
rect 9311 -6291 9391 -6221
rect 9311 -6351 9321 -6291
rect 9381 -6351 9391 -6291
rect 9767 -6221 9777 -6171
rect 10233 -6161 10293 -5994
rect 9837 -6221 9847 -6171
rect 9767 -6291 9847 -6221
rect 9767 -6351 9777 -6291
rect 9837 -6351 9847 -6291
rect 10223 -6221 10233 -6171
rect 10691 -6161 10751 -5994
rect 10293 -6221 10303 -6171
rect 10223 -6291 10303 -6221
rect 10223 -6351 10233 -6291
rect 10293 -6351 10303 -6291
rect 10681 -6221 10691 -6171
rect 11147 -6161 11207 -5994
rect 10751 -6221 10761 -6171
rect 10681 -6291 10761 -6221
rect 10681 -6351 10691 -6291
rect 10751 -6351 10761 -6291
rect 11137 -6221 11147 -6171
rect 11603 -6161 11663 -5994
rect 11207 -6221 11217 -6171
rect 11137 -6291 11217 -6221
rect 11137 -6351 11147 -6291
rect 11207 -6351 11217 -6291
rect 11593 -6221 11603 -6171
rect 12061 -6161 12121 -5994
rect 11663 -6221 11673 -6171
rect 11593 -6291 11673 -6221
rect 11593 -6351 11603 -6291
rect 11663 -6351 11673 -6291
rect 12051 -6221 12061 -6171
rect 12517 -6161 12577 -5994
rect 12121 -6221 12131 -6171
rect 12051 -6291 12131 -6221
rect 12051 -6351 12061 -6291
rect 12121 -6351 12131 -6291
rect 12507 -6221 12517 -6171
rect 12973 -6161 13033 -5994
rect 12577 -6221 12587 -6171
rect 12507 -6291 12587 -6221
rect 12507 -6351 12517 -6291
rect 12577 -6351 12587 -6291
rect 12963 -6221 12973 -6171
rect 13431 -6161 13491 -5994
rect 13033 -6221 13043 -6171
rect 12963 -6291 13043 -6221
rect 12963 -6351 12973 -6291
rect 13033 -6351 13043 -6291
rect 13421 -6221 13431 -6171
rect 13887 -6161 13947 -5994
rect 13491 -6221 13501 -6171
rect 13421 -6291 13501 -6221
rect 13421 -6351 13431 -6291
rect 13491 -6351 13501 -6291
rect 13877 -6221 13887 -6171
rect 14343 -6161 14403 -5994
rect 13947 -6221 13957 -6171
rect 13877 -6291 13957 -6221
rect 13877 -6351 13887 -6291
rect 13947 -6351 13957 -6291
rect 14333 -6221 14343 -6171
rect 14801 -6161 14861 -5994
rect 14403 -6221 14413 -6171
rect 14333 -6291 14413 -6221
rect 14333 -6351 14343 -6291
rect 14403 -6351 14413 -6291
rect 14791 -6221 14801 -6171
rect 15257 -6161 15317 -5994
rect 14861 -6221 14871 -6171
rect 14791 -6291 14871 -6221
rect 14791 -6351 14801 -6291
rect 14861 -6351 14871 -6291
rect 15247 -6221 15257 -6171
rect 15317 -6221 15327 -6171
rect 15247 -6291 15327 -6221
rect 15247 -6351 15257 -6291
rect 15317 -6351 15327 -6291
rect 171 -6653 231 -6351
rect 161 -6713 171 -6663
rect 627 -6653 687 -6351
rect 231 -6713 241 -6663
rect 161 -6783 241 -6713
rect 161 -6843 171 -6783
rect 231 -6843 241 -6783
rect 617 -6713 627 -6663
rect 1083 -6653 1143 -6351
rect 687 -6713 697 -6663
rect 617 -6783 697 -6713
rect 617 -6843 627 -6783
rect 687 -6843 697 -6783
rect 1073 -6713 1083 -6663
rect 1541 -6653 1601 -6351
rect 1143 -6713 1153 -6663
rect 1073 -6783 1153 -6713
rect 1073 -6843 1083 -6783
rect 1143 -6843 1153 -6783
rect 1531 -6713 1541 -6663
rect 1997 -6653 2057 -6351
rect 1601 -6713 1611 -6663
rect 1531 -6783 1611 -6713
rect 1531 -6843 1541 -6783
rect 1601 -6843 1611 -6783
rect 1987 -6713 1997 -6663
rect 2453 -6653 2513 -6351
rect 2057 -6713 2067 -6663
rect 1987 -6783 2067 -6713
rect 1987 -6843 1997 -6783
rect 2057 -6843 2067 -6783
rect 2443 -6713 2453 -6663
rect 2911 -6653 2971 -6351
rect 2513 -6713 2523 -6663
rect 2443 -6783 2523 -6713
rect 2443 -6843 2453 -6783
rect 2513 -6843 2523 -6783
rect 2901 -6713 2911 -6663
rect 3367 -6653 3427 -6351
rect 2971 -6713 2981 -6663
rect 2901 -6783 2981 -6713
rect 2901 -6843 2911 -6783
rect 2971 -6843 2981 -6783
rect 3357 -6713 3367 -6663
rect 3823 -6653 3883 -6351
rect 3427 -6713 3437 -6663
rect 3357 -6783 3437 -6713
rect 3357 -6843 3367 -6783
rect 3427 -6843 3437 -6783
rect 3813 -6713 3823 -6663
rect 4281 -6653 4341 -6351
rect 3883 -6713 3893 -6663
rect 3813 -6783 3893 -6713
rect 3813 -6843 3823 -6783
rect 3883 -6843 3893 -6783
rect 4271 -6713 4281 -6663
rect 4737 -6653 4797 -6351
rect 4341 -6713 4351 -6663
rect 4271 -6783 4351 -6713
rect 4271 -6843 4281 -6783
rect 4341 -6843 4351 -6783
rect 4727 -6713 4737 -6663
rect 5193 -6653 5253 -6351
rect 4797 -6713 4807 -6663
rect 4727 -6783 4807 -6713
rect 4727 -6843 4737 -6783
rect 4797 -6843 4807 -6783
rect 5183 -6713 5193 -6663
rect 5651 -6653 5711 -6351
rect 5253 -6713 5263 -6663
rect 5183 -6783 5263 -6713
rect 5183 -6843 5193 -6783
rect 5253 -6843 5263 -6783
rect 5641 -6713 5651 -6663
rect 6107 -6653 6167 -6351
rect 5711 -6713 5721 -6663
rect 5641 -6783 5721 -6713
rect 5641 -6843 5651 -6783
rect 5711 -6843 5721 -6783
rect 6097 -6713 6107 -6663
rect 6563 -6653 6623 -6351
rect 6167 -6713 6177 -6663
rect 6097 -6783 6177 -6713
rect 6097 -6843 6107 -6783
rect 6167 -6843 6177 -6783
rect 6553 -6713 6563 -6663
rect 7021 -6653 7081 -6351
rect 6623 -6713 6633 -6663
rect 6553 -6783 6633 -6713
rect 6553 -6843 6563 -6783
rect 6623 -6843 6633 -6783
rect 7011 -6713 7021 -6663
rect 7477 -6653 7537 -6351
rect 7081 -6713 7091 -6663
rect 7011 -6783 7091 -6713
rect 7011 -6843 7021 -6783
rect 7081 -6843 7091 -6783
rect 7467 -6713 7477 -6663
rect 7933 -6653 7993 -6351
rect 7537 -6713 7547 -6663
rect 7467 -6783 7547 -6713
rect 7467 -6843 7477 -6783
rect 7537 -6843 7547 -6783
rect 7923 -6713 7933 -6663
rect 8407 -6653 8467 -6351
rect 7993 -6713 8003 -6663
rect 7923 -6783 8003 -6713
rect 7923 -6843 7933 -6783
rect 7993 -6843 8003 -6783
rect 8397 -6713 8407 -6663
rect 8863 -6653 8923 -6351
rect 8467 -6713 8477 -6663
rect 8397 -6783 8477 -6713
rect 8397 -6843 8407 -6783
rect 8467 -6843 8477 -6783
rect 8853 -6713 8863 -6663
rect 9321 -6653 9381 -6351
rect 8923 -6713 8933 -6663
rect 8853 -6783 8933 -6713
rect 8853 -6843 8863 -6783
rect 8923 -6843 8933 -6783
rect 9311 -6713 9321 -6663
rect 9777 -6653 9837 -6351
rect 9381 -6713 9391 -6663
rect 9311 -6783 9391 -6713
rect 9311 -6843 9321 -6783
rect 9381 -6843 9391 -6783
rect 9767 -6713 9777 -6663
rect 10233 -6653 10293 -6351
rect 9837 -6713 9847 -6663
rect 9767 -6783 9847 -6713
rect 9767 -6843 9777 -6783
rect 9837 -6843 9847 -6783
rect 10223 -6713 10233 -6663
rect 10691 -6653 10751 -6351
rect 10293 -6713 10303 -6663
rect 10223 -6783 10303 -6713
rect 10223 -6843 10233 -6783
rect 10293 -6843 10303 -6783
rect 10681 -6713 10691 -6663
rect 11147 -6653 11207 -6351
rect 10751 -6713 10761 -6663
rect 10681 -6783 10761 -6713
rect 10681 -6843 10691 -6783
rect 10751 -6843 10761 -6783
rect 11137 -6713 11147 -6663
rect 11603 -6653 11663 -6351
rect 11207 -6713 11217 -6663
rect 11137 -6783 11217 -6713
rect 11137 -6843 11147 -6783
rect 11207 -6843 11217 -6783
rect 11593 -6713 11603 -6663
rect 12061 -6653 12121 -6351
rect 11663 -6713 11673 -6663
rect 11593 -6783 11673 -6713
rect 11593 -6843 11603 -6783
rect 11663 -6843 11673 -6783
rect 12051 -6713 12061 -6663
rect 12517 -6653 12577 -6351
rect 12121 -6713 12131 -6663
rect 12051 -6783 12131 -6713
rect 12051 -6843 12061 -6783
rect 12121 -6843 12131 -6783
rect 12507 -6713 12517 -6663
rect 12973 -6653 13033 -6351
rect 12577 -6713 12587 -6663
rect 12507 -6783 12587 -6713
rect 12507 -6843 12517 -6783
rect 12577 -6843 12587 -6783
rect 12963 -6713 12973 -6663
rect 13431 -6653 13491 -6351
rect 13033 -6713 13043 -6663
rect 12963 -6783 13043 -6713
rect 12963 -6843 12973 -6783
rect 13033 -6843 13043 -6783
rect 13421 -6713 13431 -6663
rect 13887 -6653 13947 -6351
rect 13491 -6713 13501 -6663
rect 13421 -6783 13501 -6713
rect 13421 -6843 13431 -6783
rect 13491 -6843 13501 -6783
rect 13877 -6713 13887 -6663
rect 14343 -6653 14403 -6351
rect 13947 -6713 13957 -6663
rect 13877 -6783 13957 -6713
rect 13877 -6843 13887 -6783
rect 13947 -6843 13957 -6783
rect 14333 -6713 14343 -6663
rect 14801 -6653 14861 -6351
rect 14403 -6713 14413 -6663
rect 14333 -6783 14413 -6713
rect 14333 -6843 14343 -6783
rect 14403 -6843 14413 -6783
rect 14791 -6713 14801 -6663
rect 15257 -6653 15317 -6351
rect 14861 -6713 14871 -6663
rect 14791 -6783 14871 -6713
rect 14791 -6843 14801 -6783
rect 14861 -6843 14871 -6783
rect 15247 -6713 15257 -6663
rect 15317 -6713 15327 -6663
rect 15247 -6783 15327 -6713
rect 15247 -6843 15257 -6783
rect 15317 -6843 15327 -6783
rect 171 -7169 231 -6843
rect 161 -7229 171 -7179
rect 627 -7169 687 -6843
rect 231 -7229 241 -7179
rect 161 -7299 241 -7229
rect 161 -7359 171 -7299
rect 231 -7359 241 -7299
rect 617 -7229 627 -7179
rect 1083 -7169 1143 -6843
rect 687 -7229 697 -7179
rect 617 -7299 697 -7229
rect 617 -7359 627 -7299
rect 687 -7359 697 -7299
rect 1073 -7229 1083 -7179
rect 1541 -7169 1601 -6843
rect 1143 -7229 1153 -7179
rect 1073 -7299 1153 -7229
rect 1073 -7359 1083 -7299
rect 1143 -7359 1153 -7299
rect 1531 -7229 1541 -7179
rect 1997 -7169 2057 -6843
rect 1601 -7229 1611 -7179
rect 1531 -7299 1611 -7229
rect 1531 -7359 1541 -7299
rect 1601 -7359 1611 -7299
rect 1987 -7229 1997 -7179
rect 2453 -7169 2513 -6843
rect 2057 -7229 2067 -7179
rect 1987 -7299 2067 -7229
rect 1987 -7359 1997 -7299
rect 2057 -7359 2067 -7299
rect 2443 -7229 2453 -7179
rect 2911 -7169 2971 -6843
rect 2513 -7229 2523 -7179
rect 2443 -7299 2523 -7229
rect 2443 -7359 2453 -7299
rect 2513 -7359 2523 -7299
rect 2901 -7229 2911 -7179
rect 3367 -7169 3427 -6843
rect 2971 -7229 2981 -7179
rect 2901 -7299 2981 -7229
rect 2901 -7359 2911 -7299
rect 2971 -7359 2981 -7299
rect 3357 -7229 3367 -7179
rect 3823 -7169 3883 -6843
rect 3427 -7229 3437 -7179
rect 3357 -7299 3437 -7229
rect 3357 -7359 3367 -7299
rect 3427 -7359 3437 -7299
rect 3813 -7229 3823 -7179
rect 4281 -7169 4341 -6843
rect 3883 -7229 3893 -7179
rect 3813 -7299 3893 -7229
rect 3813 -7359 3823 -7299
rect 3883 -7359 3893 -7299
rect 4271 -7229 4281 -7179
rect 4737 -7169 4797 -6843
rect 4341 -7229 4351 -7179
rect 4271 -7299 4351 -7229
rect 4271 -7359 4281 -7299
rect 4341 -7359 4351 -7299
rect 4727 -7229 4737 -7179
rect 5193 -7169 5253 -6843
rect 4797 -7229 4807 -7179
rect 4727 -7299 4807 -7229
rect 4727 -7359 4737 -7299
rect 4797 -7359 4807 -7299
rect 5183 -7229 5193 -7179
rect 5651 -7169 5711 -6843
rect 5253 -7229 5263 -7179
rect 5183 -7299 5263 -7229
rect 5183 -7359 5193 -7299
rect 5253 -7359 5263 -7299
rect 5641 -7229 5651 -7179
rect 6107 -7169 6167 -6843
rect 5711 -7229 5721 -7179
rect 5641 -7299 5721 -7229
rect 5641 -7359 5651 -7299
rect 5711 -7359 5721 -7299
rect 6097 -7229 6107 -7179
rect 6563 -7169 6623 -6843
rect 6167 -7229 6177 -7179
rect 6097 -7299 6177 -7229
rect 6097 -7359 6107 -7299
rect 6167 -7359 6177 -7299
rect 6553 -7229 6563 -7179
rect 7021 -7169 7081 -6843
rect 6623 -7229 6633 -7179
rect 6553 -7299 6633 -7229
rect 6553 -7359 6563 -7299
rect 6623 -7359 6633 -7299
rect 7011 -7229 7021 -7179
rect 7477 -7169 7537 -6843
rect 7081 -7229 7091 -7179
rect 7011 -7299 7091 -7229
rect 7011 -7359 7021 -7299
rect 7081 -7359 7091 -7299
rect 7467 -7229 7477 -7179
rect 7933 -7169 7993 -6843
rect 7537 -7229 7547 -7179
rect 7467 -7299 7547 -7229
rect 7467 -7359 7477 -7299
rect 7537 -7359 7547 -7299
rect 7923 -7229 7933 -7179
rect 8407 -7169 8467 -6843
rect 7993 -7229 8003 -7179
rect 7923 -7299 8003 -7229
rect 7923 -7359 7933 -7299
rect 7993 -7359 8003 -7299
rect 8397 -7229 8407 -7179
rect 8863 -7169 8923 -6843
rect 8467 -7229 8477 -7179
rect 8397 -7299 8477 -7229
rect 8397 -7359 8407 -7299
rect 8467 -7359 8477 -7299
rect 8853 -7229 8863 -7179
rect 9321 -7169 9381 -6843
rect 8923 -7229 8933 -7179
rect 8853 -7299 8933 -7229
rect 8853 -7359 8863 -7299
rect 8923 -7359 8933 -7299
rect 9311 -7229 9321 -7179
rect 9777 -7169 9837 -6843
rect 9381 -7229 9391 -7179
rect 9311 -7299 9391 -7229
rect 9311 -7359 9321 -7299
rect 9381 -7359 9391 -7299
rect 9767 -7229 9777 -7179
rect 10233 -7169 10293 -6843
rect 9837 -7229 9847 -7179
rect 9767 -7299 9847 -7229
rect 9767 -7359 9777 -7299
rect 9837 -7359 9847 -7299
rect 10223 -7229 10233 -7179
rect 10691 -7169 10751 -6843
rect 10293 -7229 10303 -7179
rect 10223 -7299 10303 -7229
rect 10223 -7359 10233 -7299
rect 10293 -7359 10303 -7299
rect 10681 -7229 10691 -7179
rect 11147 -7169 11207 -6843
rect 10751 -7229 10761 -7179
rect 10681 -7299 10761 -7229
rect 10681 -7359 10691 -7299
rect 10751 -7359 10761 -7299
rect 11137 -7229 11147 -7179
rect 11603 -7169 11663 -6843
rect 11207 -7229 11217 -7179
rect 11137 -7299 11217 -7229
rect 11137 -7359 11147 -7299
rect 11207 -7359 11217 -7299
rect 11593 -7229 11603 -7179
rect 12061 -7169 12121 -6843
rect 11663 -7229 11673 -7179
rect 11593 -7299 11673 -7229
rect 11593 -7359 11603 -7299
rect 11663 -7359 11673 -7299
rect 12051 -7229 12061 -7179
rect 12517 -7169 12577 -6843
rect 12121 -7229 12131 -7179
rect 12051 -7299 12131 -7229
rect 12051 -7359 12061 -7299
rect 12121 -7359 12131 -7299
rect 12507 -7229 12517 -7179
rect 12973 -7169 13033 -6843
rect 12577 -7229 12587 -7179
rect 12507 -7299 12587 -7229
rect 12507 -7359 12517 -7299
rect 12577 -7359 12587 -7299
rect 12963 -7229 12973 -7179
rect 13431 -7169 13491 -6843
rect 13033 -7229 13043 -7179
rect 12963 -7299 13043 -7229
rect 12963 -7359 12973 -7299
rect 13033 -7359 13043 -7299
rect 13421 -7229 13431 -7179
rect 13887 -7169 13947 -6843
rect 13491 -7229 13501 -7179
rect 13421 -7299 13501 -7229
rect 13421 -7359 13431 -7299
rect 13491 -7359 13501 -7299
rect 13877 -7229 13887 -7179
rect 14343 -7169 14403 -6843
rect 13947 -7229 13957 -7179
rect 13877 -7299 13957 -7229
rect 13877 -7359 13887 -7299
rect 13947 -7359 13957 -7299
rect 14333 -7229 14343 -7179
rect 14801 -7169 14861 -6843
rect 14403 -7229 14413 -7179
rect 14333 -7299 14413 -7229
rect 14333 -7359 14343 -7299
rect 14403 -7359 14413 -7299
rect 14791 -7229 14801 -7179
rect 15257 -7169 15317 -6843
rect 14861 -7229 14871 -7179
rect 14791 -7299 14871 -7229
rect 14791 -7359 14801 -7299
rect 14861 -7359 14871 -7299
rect 15247 -7229 15257 -7179
rect 15317 -7229 15327 -7179
rect 15247 -7299 15327 -7229
rect 15247 -7359 15257 -7299
rect 15317 -7359 15327 -7299
rect 171 -7671 231 -7359
rect 161 -7731 171 -7681
rect 627 -7671 687 -7359
rect 231 -7731 241 -7681
rect 161 -7801 241 -7731
rect 161 -7861 171 -7801
rect 231 -7861 241 -7801
rect 617 -7731 627 -7681
rect 1083 -7671 1143 -7359
rect 687 -7731 697 -7681
rect 617 -7801 697 -7731
rect 617 -7861 627 -7801
rect 687 -7861 697 -7801
rect 1073 -7731 1083 -7681
rect 1541 -7671 1601 -7359
rect 1143 -7731 1153 -7681
rect 1073 -7801 1153 -7731
rect 1073 -7861 1083 -7801
rect 1143 -7861 1153 -7801
rect 1531 -7731 1541 -7681
rect 1997 -7671 2057 -7359
rect 1601 -7731 1611 -7681
rect 1531 -7801 1611 -7731
rect 1531 -7861 1541 -7801
rect 1601 -7861 1611 -7801
rect 1987 -7731 1997 -7681
rect 2453 -7671 2513 -7359
rect 2057 -7731 2067 -7681
rect 1987 -7801 2067 -7731
rect 1987 -7861 1997 -7801
rect 2057 -7861 2067 -7801
rect 2443 -7731 2453 -7681
rect 2911 -7671 2971 -7359
rect 2513 -7731 2523 -7681
rect 2443 -7801 2523 -7731
rect 2443 -7861 2453 -7801
rect 2513 -7861 2523 -7801
rect 2901 -7731 2911 -7681
rect 3367 -7671 3427 -7359
rect 2971 -7731 2981 -7681
rect 2901 -7801 2981 -7731
rect 2901 -7861 2911 -7801
rect 2971 -7861 2981 -7801
rect 3357 -7731 3367 -7681
rect 3823 -7671 3883 -7359
rect 3427 -7731 3437 -7681
rect 3357 -7801 3437 -7731
rect 3357 -7861 3367 -7801
rect 3427 -7861 3437 -7801
rect 3813 -7731 3823 -7681
rect 4281 -7671 4341 -7359
rect 3883 -7731 3893 -7681
rect 3813 -7801 3893 -7731
rect 3813 -7861 3823 -7801
rect 3883 -7861 3893 -7801
rect 4271 -7731 4281 -7681
rect 4737 -7671 4797 -7359
rect 4341 -7731 4351 -7681
rect 4271 -7801 4351 -7731
rect 4271 -7861 4281 -7801
rect 4341 -7861 4351 -7801
rect 4727 -7731 4737 -7681
rect 5193 -7671 5253 -7359
rect 4797 -7731 4807 -7681
rect 4727 -7801 4807 -7731
rect 4727 -7861 4737 -7801
rect 4797 -7861 4807 -7801
rect 5183 -7731 5193 -7681
rect 5651 -7671 5711 -7359
rect 5253 -7731 5263 -7681
rect 5183 -7801 5263 -7731
rect 5183 -7861 5193 -7801
rect 5253 -7861 5263 -7801
rect 5641 -7731 5651 -7681
rect 6107 -7671 6167 -7359
rect 5711 -7731 5721 -7681
rect 5641 -7801 5721 -7731
rect 5641 -7861 5651 -7801
rect 5711 -7861 5721 -7801
rect 6097 -7731 6107 -7681
rect 6563 -7671 6623 -7359
rect 6167 -7731 6177 -7681
rect 6097 -7801 6177 -7731
rect 6097 -7861 6107 -7801
rect 6167 -7861 6177 -7801
rect 6553 -7731 6563 -7681
rect 7021 -7671 7081 -7359
rect 6623 -7731 6633 -7681
rect 6553 -7801 6633 -7731
rect 6553 -7861 6563 -7801
rect 6623 -7861 6633 -7801
rect 7011 -7731 7021 -7681
rect 7477 -7671 7537 -7359
rect 7081 -7731 7091 -7681
rect 7011 -7801 7091 -7731
rect 7011 -7861 7021 -7801
rect 7081 -7861 7091 -7801
rect 7467 -7731 7477 -7681
rect 7933 -7671 7993 -7359
rect 7537 -7731 7547 -7681
rect 7467 -7801 7547 -7731
rect 7467 -7861 7477 -7801
rect 7537 -7861 7547 -7801
rect 7923 -7731 7933 -7681
rect 8407 -7671 8467 -7359
rect 7993 -7731 8003 -7681
rect 7923 -7801 8003 -7731
rect 7923 -7861 7933 -7801
rect 7993 -7861 8003 -7801
rect 8397 -7731 8407 -7681
rect 8863 -7671 8923 -7359
rect 8467 -7731 8477 -7681
rect 8397 -7801 8477 -7731
rect 8397 -7861 8407 -7801
rect 8467 -7861 8477 -7801
rect 8853 -7731 8863 -7681
rect 9321 -7671 9381 -7359
rect 8923 -7731 8933 -7681
rect 8853 -7801 8933 -7731
rect 8853 -7861 8863 -7801
rect 8923 -7861 8933 -7801
rect 9311 -7731 9321 -7681
rect 9777 -7671 9837 -7359
rect 9381 -7731 9391 -7681
rect 9311 -7801 9391 -7731
rect 9311 -7861 9321 -7801
rect 9381 -7861 9391 -7801
rect 9767 -7731 9777 -7681
rect 10233 -7671 10293 -7359
rect 9837 -7731 9847 -7681
rect 9767 -7801 9847 -7731
rect 9767 -7861 9777 -7801
rect 9837 -7861 9847 -7801
rect 10223 -7731 10233 -7681
rect 10691 -7671 10751 -7359
rect 10293 -7731 10303 -7681
rect 10223 -7801 10303 -7731
rect 10223 -7861 10233 -7801
rect 10293 -7861 10303 -7801
rect 10681 -7731 10691 -7681
rect 11147 -7671 11207 -7359
rect 10751 -7731 10761 -7681
rect 10681 -7801 10761 -7731
rect 10681 -7861 10691 -7801
rect 10751 -7861 10761 -7801
rect 11137 -7731 11147 -7681
rect 11603 -7671 11663 -7359
rect 11207 -7731 11217 -7681
rect 11137 -7801 11217 -7731
rect 11137 -7861 11147 -7801
rect 11207 -7861 11217 -7801
rect 11593 -7731 11603 -7681
rect 12061 -7671 12121 -7359
rect 11663 -7731 11673 -7681
rect 11593 -7801 11673 -7731
rect 11593 -7861 11603 -7801
rect 11663 -7861 11673 -7801
rect 12051 -7731 12061 -7681
rect 12517 -7671 12577 -7359
rect 12121 -7731 12131 -7681
rect 12051 -7801 12131 -7731
rect 12051 -7861 12061 -7801
rect 12121 -7861 12131 -7801
rect 12507 -7731 12517 -7681
rect 12973 -7671 13033 -7359
rect 12577 -7731 12587 -7681
rect 12507 -7801 12587 -7731
rect 12507 -7861 12517 -7801
rect 12577 -7861 12587 -7801
rect 12963 -7731 12973 -7681
rect 13431 -7671 13491 -7359
rect 13033 -7731 13043 -7681
rect 12963 -7801 13043 -7731
rect 12963 -7861 12973 -7801
rect 13033 -7861 13043 -7801
rect 13421 -7731 13431 -7681
rect 13887 -7671 13947 -7359
rect 13491 -7731 13501 -7681
rect 13421 -7801 13501 -7731
rect 13421 -7861 13431 -7801
rect 13491 -7861 13501 -7801
rect 13877 -7731 13887 -7681
rect 14343 -7671 14403 -7359
rect 13947 -7731 13957 -7681
rect 13877 -7801 13957 -7731
rect 13877 -7861 13887 -7801
rect 13947 -7861 13957 -7801
rect 14333 -7731 14343 -7681
rect 14801 -7671 14861 -7359
rect 14403 -7731 14413 -7681
rect 14333 -7801 14413 -7731
rect 14333 -7861 14343 -7801
rect 14403 -7861 14413 -7801
rect 14791 -7731 14801 -7681
rect 15257 -7671 15317 -7359
rect 14861 -7731 14871 -7681
rect 14791 -7801 14871 -7731
rect 14791 -7861 14801 -7801
rect 14861 -7861 14871 -7801
rect 15247 -7731 15257 -7681
rect 15317 -7731 15327 -7681
rect 15247 -7801 15327 -7731
rect 15247 -7861 15257 -7801
rect 15317 -7861 15327 -7801
rect 171 -8163 231 -7861
rect 161 -8223 171 -8173
rect 627 -8163 687 -7861
rect 231 -8223 241 -8173
rect 161 -8293 241 -8223
rect 161 -8353 171 -8293
rect 231 -8353 241 -8293
rect 617 -8223 627 -8173
rect 1083 -8163 1143 -7861
rect 687 -8223 697 -8173
rect 617 -8293 697 -8223
rect 617 -8353 627 -8293
rect 687 -8353 697 -8293
rect 1073 -8223 1083 -8173
rect 1541 -8163 1601 -7861
rect 1143 -8223 1153 -8173
rect 1073 -8293 1153 -8223
rect 1073 -8353 1083 -8293
rect 1143 -8353 1153 -8293
rect 1531 -8223 1541 -8173
rect 1997 -8163 2057 -7861
rect 1601 -8223 1611 -8173
rect 1531 -8293 1611 -8223
rect 1531 -8353 1541 -8293
rect 1601 -8353 1611 -8293
rect 1987 -8223 1997 -8173
rect 2453 -8163 2513 -7861
rect 2057 -8223 2067 -8173
rect 1987 -8293 2067 -8223
rect 1987 -8353 1997 -8293
rect 2057 -8353 2067 -8293
rect 2443 -8223 2453 -8173
rect 2911 -8163 2971 -7861
rect 2513 -8223 2523 -8173
rect 2443 -8293 2523 -8223
rect 2443 -8353 2453 -8293
rect 2513 -8353 2523 -8293
rect 2901 -8223 2911 -8173
rect 3367 -8163 3427 -7861
rect 2971 -8223 2981 -8173
rect 2901 -8293 2981 -8223
rect 2901 -8353 2911 -8293
rect 2971 -8353 2981 -8293
rect 3357 -8223 3367 -8173
rect 3823 -8163 3883 -7861
rect 3427 -8223 3437 -8173
rect 3357 -8293 3437 -8223
rect 3357 -8353 3367 -8293
rect 3427 -8353 3437 -8293
rect 3813 -8223 3823 -8173
rect 4281 -8163 4341 -7861
rect 3883 -8223 3893 -8173
rect 3813 -8293 3893 -8223
rect 3813 -8353 3823 -8293
rect 3883 -8353 3893 -8293
rect 4271 -8223 4281 -8173
rect 4737 -8163 4797 -7861
rect 4341 -8223 4351 -8173
rect 4271 -8293 4351 -8223
rect 4271 -8353 4281 -8293
rect 4341 -8353 4351 -8293
rect 4727 -8223 4737 -8173
rect 5193 -8163 5253 -7861
rect 4797 -8223 4807 -8173
rect 4727 -8293 4807 -8223
rect 4727 -8353 4737 -8293
rect 4797 -8353 4807 -8293
rect 5183 -8223 5193 -8173
rect 5651 -8163 5711 -7861
rect 5253 -8223 5263 -8173
rect 5183 -8293 5263 -8223
rect 5183 -8353 5193 -8293
rect 5253 -8353 5263 -8293
rect 5641 -8223 5651 -8173
rect 6107 -8163 6167 -7861
rect 5711 -8223 5721 -8173
rect 5641 -8293 5721 -8223
rect 5641 -8353 5651 -8293
rect 5711 -8353 5721 -8293
rect 6097 -8223 6107 -8173
rect 6563 -8163 6623 -7861
rect 6167 -8223 6177 -8173
rect 6097 -8293 6177 -8223
rect 6097 -8353 6107 -8293
rect 6167 -8353 6177 -8293
rect 6553 -8223 6563 -8173
rect 7021 -8163 7081 -7861
rect 6623 -8223 6633 -8173
rect 6553 -8293 6633 -8223
rect 6553 -8353 6563 -8293
rect 6623 -8353 6633 -8293
rect 7011 -8223 7021 -8173
rect 7477 -8163 7537 -7861
rect 7081 -8223 7091 -8173
rect 7011 -8293 7091 -8223
rect 7011 -8353 7021 -8293
rect 7081 -8353 7091 -8293
rect 7467 -8223 7477 -8173
rect 7933 -8163 7993 -7861
rect 7537 -8223 7547 -8173
rect 7467 -8293 7547 -8223
rect 7467 -8353 7477 -8293
rect 7537 -8353 7547 -8293
rect 7923 -8223 7933 -8173
rect 8407 -8163 8467 -7861
rect 7993 -8223 8003 -8173
rect 7923 -8293 8003 -8223
rect 7923 -8353 7933 -8293
rect 7993 -8353 8003 -8293
rect 8397 -8223 8407 -8173
rect 8863 -8163 8923 -7861
rect 8467 -8223 8477 -8173
rect 8397 -8293 8477 -8223
rect 8397 -8353 8407 -8293
rect 8467 -8353 8477 -8293
rect 8853 -8223 8863 -8173
rect 9321 -8163 9381 -7861
rect 8923 -8223 8933 -8173
rect 8853 -8293 8933 -8223
rect 8853 -8353 8863 -8293
rect 8923 -8353 8933 -8293
rect 9311 -8223 9321 -8173
rect 9777 -8163 9837 -7861
rect 9381 -8223 9391 -8173
rect 9311 -8293 9391 -8223
rect 9311 -8353 9321 -8293
rect 9381 -8353 9391 -8293
rect 9767 -8223 9777 -8173
rect 10233 -8163 10293 -7861
rect 9837 -8223 9847 -8173
rect 9767 -8293 9847 -8223
rect 9767 -8353 9777 -8293
rect 9837 -8353 9847 -8293
rect 10223 -8223 10233 -8173
rect 10691 -8163 10751 -7861
rect 10293 -8223 10303 -8173
rect 10223 -8293 10303 -8223
rect 10223 -8353 10233 -8293
rect 10293 -8353 10303 -8293
rect 10681 -8223 10691 -8173
rect 11147 -8163 11207 -7861
rect 10751 -8223 10761 -8173
rect 10681 -8293 10761 -8223
rect 10681 -8353 10691 -8293
rect 10751 -8353 10761 -8293
rect 11137 -8223 11147 -8173
rect 11603 -8163 11663 -7861
rect 11207 -8223 11217 -8173
rect 11137 -8293 11217 -8223
rect 11137 -8353 11147 -8293
rect 11207 -8353 11217 -8293
rect 11593 -8223 11603 -8173
rect 12061 -8163 12121 -7861
rect 11663 -8223 11673 -8173
rect 11593 -8293 11673 -8223
rect 11593 -8353 11603 -8293
rect 11663 -8353 11673 -8293
rect 12051 -8223 12061 -8173
rect 12517 -8163 12577 -7861
rect 12121 -8223 12131 -8173
rect 12051 -8293 12131 -8223
rect 12051 -8353 12061 -8293
rect 12121 -8353 12131 -8293
rect 12507 -8223 12517 -8173
rect 12973 -8163 13033 -7861
rect 12577 -8223 12587 -8173
rect 12507 -8293 12587 -8223
rect 12507 -8353 12517 -8293
rect 12577 -8353 12587 -8293
rect 12963 -8223 12973 -8173
rect 13431 -8163 13491 -7861
rect 13033 -8223 13043 -8173
rect 12963 -8293 13043 -8223
rect 12963 -8353 12973 -8293
rect 13033 -8353 13043 -8293
rect 13421 -8223 13431 -8173
rect 13887 -8163 13947 -7861
rect 13491 -8223 13501 -8173
rect 13421 -8293 13501 -8223
rect 13421 -8353 13431 -8293
rect 13491 -8353 13501 -8293
rect 13877 -8223 13887 -8173
rect 14343 -8163 14403 -7861
rect 13947 -8223 13957 -8173
rect 13877 -8293 13957 -8223
rect 13877 -8353 13887 -8293
rect 13947 -8353 13957 -8293
rect 14333 -8223 14343 -8173
rect 14801 -8163 14861 -7861
rect 14403 -8223 14413 -8173
rect 14333 -8293 14413 -8223
rect 14333 -8353 14343 -8293
rect 14403 -8353 14413 -8293
rect 14791 -8223 14801 -8173
rect 15257 -8163 15317 -7861
rect 14861 -8223 14871 -8173
rect 14791 -8293 14871 -8223
rect 14791 -8353 14801 -8293
rect 14861 -8353 14871 -8293
rect 15247 -8223 15257 -8173
rect 15317 -8223 15327 -8173
rect 15247 -8293 15327 -8223
rect 15247 -8353 15257 -8293
rect 15317 -8353 15327 -8293
rect 171 -8657 231 -8353
rect 161 -8717 171 -8667
rect 627 -8657 687 -8353
rect 231 -8717 241 -8667
rect 161 -8787 241 -8717
rect 161 -8847 171 -8787
rect 231 -8847 241 -8787
rect 617 -8717 627 -8667
rect 1083 -8657 1143 -8353
rect 687 -8717 697 -8667
rect 617 -8787 697 -8717
rect 617 -8847 627 -8787
rect 687 -8847 697 -8787
rect 1073 -8717 1083 -8667
rect 1541 -8657 1601 -8353
rect 1143 -8717 1153 -8667
rect 1073 -8787 1153 -8717
rect 1073 -8847 1083 -8787
rect 1143 -8847 1153 -8787
rect 1531 -8717 1541 -8667
rect 1997 -8657 2057 -8353
rect 1601 -8717 1611 -8667
rect 1531 -8787 1611 -8717
rect 1531 -8847 1541 -8787
rect 1601 -8847 1611 -8787
rect 1987 -8717 1997 -8667
rect 2453 -8657 2513 -8353
rect 2057 -8717 2067 -8667
rect 1987 -8787 2067 -8717
rect 1987 -8847 1997 -8787
rect 2057 -8847 2067 -8787
rect 2443 -8717 2453 -8667
rect 2911 -8657 2971 -8353
rect 2513 -8717 2523 -8667
rect 2443 -8787 2523 -8717
rect 2443 -8847 2453 -8787
rect 2513 -8847 2523 -8787
rect 2901 -8717 2911 -8667
rect 3367 -8657 3427 -8353
rect 2971 -8717 2981 -8667
rect 2901 -8787 2981 -8717
rect 2901 -8847 2911 -8787
rect 2971 -8847 2981 -8787
rect 3357 -8717 3367 -8667
rect 3823 -8657 3883 -8353
rect 3427 -8717 3437 -8667
rect 3357 -8787 3437 -8717
rect 3357 -8847 3367 -8787
rect 3427 -8847 3437 -8787
rect 3813 -8717 3823 -8667
rect 4281 -8657 4341 -8353
rect 3883 -8717 3893 -8667
rect 3813 -8787 3893 -8717
rect 3813 -8847 3823 -8787
rect 3883 -8847 3893 -8787
rect 4271 -8717 4281 -8667
rect 4737 -8657 4797 -8353
rect 4341 -8717 4351 -8667
rect 4271 -8787 4351 -8717
rect 4271 -8847 4281 -8787
rect 4341 -8847 4351 -8787
rect 4727 -8717 4737 -8667
rect 5193 -8657 5253 -8353
rect 4797 -8717 4807 -8667
rect 4727 -8787 4807 -8717
rect 4727 -8847 4737 -8787
rect 4797 -8847 4807 -8787
rect 5183 -8717 5193 -8667
rect 5651 -8657 5711 -8353
rect 5253 -8717 5263 -8667
rect 5183 -8787 5263 -8717
rect 5183 -8847 5193 -8787
rect 5253 -8847 5263 -8787
rect 5641 -8717 5651 -8667
rect 6107 -8657 6167 -8353
rect 5711 -8717 5721 -8667
rect 5641 -8787 5721 -8717
rect 5641 -8847 5651 -8787
rect 5711 -8847 5721 -8787
rect 6097 -8717 6107 -8667
rect 6563 -8657 6623 -8353
rect 6167 -8717 6177 -8667
rect 6097 -8787 6177 -8717
rect 6097 -8847 6107 -8787
rect 6167 -8847 6177 -8787
rect 6553 -8717 6563 -8667
rect 7021 -8657 7081 -8353
rect 6623 -8717 6633 -8667
rect 6553 -8787 6633 -8717
rect 6553 -8847 6563 -8787
rect 6623 -8847 6633 -8787
rect 7011 -8717 7021 -8667
rect 7477 -8657 7537 -8353
rect 7081 -8717 7091 -8667
rect 7011 -8787 7091 -8717
rect 7011 -8847 7021 -8787
rect 7081 -8847 7091 -8787
rect 7467 -8717 7477 -8667
rect 7933 -8657 7993 -8353
rect 7537 -8717 7547 -8667
rect 7467 -8787 7547 -8717
rect 7467 -8847 7477 -8787
rect 7537 -8847 7547 -8787
rect 7923 -8717 7933 -8667
rect 8407 -8657 8467 -8353
rect 7993 -8717 8003 -8667
rect 7923 -8787 8003 -8717
rect 7923 -8847 7933 -8787
rect 7993 -8847 8003 -8787
rect 8397 -8717 8407 -8667
rect 8863 -8657 8923 -8353
rect 8467 -8717 8477 -8667
rect 8397 -8787 8477 -8717
rect 8397 -8847 8407 -8787
rect 8467 -8847 8477 -8787
rect 8853 -8717 8863 -8667
rect 9321 -8657 9381 -8353
rect 8923 -8717 8933 -8667
rect 8853 -8787 8933 -8717
rect 8853 -8847 8863 -8787
rect 8923 -8847 8933 -8787
rect 9311 -8717 9321 -8667
rect 9777 -8657 9837 -8353
rect 9381 -8717 9391 -8667
rect 9311 -8787 9391 -8717
rect 9311 -8847 9321 -8787
rect 9381 -8847 9391 -8787
rect 9767 -8717 9777 -8667
rect 10233 -8657 10293 -8353
rect 9837 -8717 9847 -8667
rect 9767 -8787 9847 -8717
rect 9767 -8847 9777 -8787
rect 9837 -8847 9847 -8787
rect 10223 -8717 10233 -8667
rect 10691 -8657 10751 -8353
rect 10293 -8717 10303 -8667
rect 10223 -8787 10303 -8717
rect 10223 -8847 10233 -8787
rect 10293 -8847 10303 -8787
rect 10681 -8717 10691 -8667
rect 11147 -8657 11207 -8353
rect 10751 -8717 10761 -8667
rect 10681 -8787 10761 -8717
rect 10681 -8847 10691 -8787
rect 10751 -8847 10761 -8787
rect 11137 -8717 11147 -8667
rect 11603 -8657 11663 -8353
rect 11207 -8717 11217 -8667
rect 11137 -8787 11217 -8717
rect 11137 -8847 11147 -8787
rect 11207 -8847 11217 -8787
rect 11593 -8717 11603 -8667
rect 12061 -8657 12121 -8353
rect 11663 -8717 11673 -8667
rect 11593 -8787 11673 -8717
rect 11593 -8847 11603 -8787
rect 11663 -8847 11673 -8787
rect 12051 -8717 12061 -8667
rect 12517 -8657 12577 -8353
rect 12121 -8717 12131 -8667
rect 12051 -8787 12131 -8717
rect 12051 -8847 12061 -8787
rect 12121 -8847 12131 -8787
rect 12507 -8717 12517 -8667
rect 12973 -8657 13033 -8353
rect 12577 -8717 12587 -8667
rect 12507 -8787 12587 -8717
rect 12507 -8847 12517 -8787
rect 12577 -8847 12587 -8787
rect 12963 -8717 12973 -8667
rect 13431 -8657 13491 -8353
rect 13033 -8717 13043 -8667
rect 12963 -8787 13043 -8717
rect 12963 -8847 12973 -8787
rect 13033 -8847 13043 -8787
rect 13421 -8717 13431 -8667
rect 13887 -8657 13947 -8353
rect 13491 -8717 13501 -8667
rect 13421 -8787 13501 -8717
rect 13421 -8847 13431 -8787
rect 13491 -8847 13501 -8787
rect 13877 -8717 13887 -8667
rect 14343 -8657 14403 -8353
rect 13947 -8717 13957 -8667
rect 13877 -8787 13957 -8717
rect 13877 -8847 13887 -8787
rect 13947 -8847 13957 -8787
rect 14333 -8717 14343 -8667
rect 14801 -8657 14861 -8353
rect 14403 -8717 14413 -8667
rect 14333 -8787 14413 -8717
rect 14333 -8847 14343 -8787
rect 14403 -8847 14413 -8787
rect 14791 -8717 14801 -8667
rect 15257 -8657 15317 -8353
rect 14861 -8717 14871 -8667
rect 14791 -8787 14871 -8717
rect 14791 -8847 14801 -8787
rect 14861 -8847 14871 -8787
rect 15247 -8717 15257 -8667
rect 15317 -8717 15327 -8667
rect 15247 -8787 15327 -8717
rect 15247 -8847 15257 -8787
rect 15317 -8847 15327 -8787
rect 171 -9159 231 -8847
rect 161 -9219 171 -9169
rect 627 -9159 687 -8847
rect 231 -9219 241 -9169
rect 161 -9289 241 -9219
rect 161 -9349 171 -9289
rect 231 -9349 241 -9289
rect 617 -9219 627 -9169
rect 1083 -9159 1143 -8847
rect 687 -9219 697 -9169
rect 617 -9289 697 -9219
rect 617 -9349 627 -9289
rect 687 -9349 697 -9289
rect 1073 -9219 1083 -9169
rect 1541 -9159 1601 -8847
rect 1143 -9219 1153 -9169
rect 1073 -9289 1153 -9219
rect 1073 -9349 1083 -9289
rect 1143 -9349 1153 -9289
rect 1531 -9219 1541 -9169
rect 1997 -9159 2057 -8847
rect 1601 -9219 1611 -9169
rect 1531 -9289 1611 -9219
rect 1531 -9349 1541 -9289
rect 1601 -9349 1611 -9289
rect 1987 -9219 1997 -9169
rect 2453 -9159 2513 -8847
rect 2057 -9219 2067 -9169
rect 1987 -9289 2067 -9219
rect 1987 -9349 1997 -9289
rect 2057 -9349 2067 -9289
rect 2443 -9219 2453 -9169
rect 2911 -9159 2971 -8847
rect 2513 -9219 2523 -9169
rect 2443 -9289 2523 -9219
rect 2443 -9349 2453 -9289
rect 2513 -9349 2523 -9289
rect 2901 -9219 2911 -9169
rect 3367 -9159 3427 -8847
rect 2971 -9219 2981 -9169
rect 2901 -9289 2981 -9219
rect 2901 -9349 2911 -9289
rect 2971 -9349 2981 -9289
rect 3357 -9219 3367 -9169
rect 3823 -9159 3883 -8847
rect 3427 -9219 3437 -9169
rect 3357 -9289 3437 -9219
rect 3357 -9349 3367 -9289
rect 3427 -9349 3437 -9289
rect 3813 -9219 3823 -9169
rect 4281 -9159 4341 -8847
rect 3883 -9219 3893 -9169
rect 3813 -9289 3893 -9219
rect 3813 -9349 3823 -9289
rect 3883 -9349 3893 -9289
rect 4271 -9219 4281 -9169
rect 4737 -9159 4797 -8847
rect 4341 -9219 4351 -9169
rect 4271 -9289 4351 -9219
rect 4271 -9349 4281 -9289
rect 4341 -9349 4351 -9289
rect 4727 -9219 4737 -9169
rect 5193 -9159 5253 -8847
rect 4797 -9219 4807 -9169
rect 4727 -9289 4807 -9219
rect 4727 -9349 4737 -9289
rect 4797 -9349 4807 -9289
rect 5183 -9219 5193 -9169
rect 5651 -9159 5711 -8847
rect 5253 -9219 5263 -9169
rect 5183 -9289 5263 -9219
rect 5183 -9349 5193 -9289
rect 5253 -9349 5263 -9289
rect 5641 -9219 5651 -9169
rect 6107 -9159 6167 -8847
rect 5711 -9219 5721 -9169
rect 5641 -9289 5721 -9219
rect 5641 -9349 5651 -9289
rect 5711 -9349 5721 -9289
rect 6097 -9219 6107 -9169
rect 6563 -9159 6623 -8847
rect 6167 -9219 6177 -9169
rect 6097 -9289 6177 -9219
rect 6097 -9349 6107 -9289
rect 6167 -9349 6177 -9289
rect 6553 -9219 6563 -9169
rect 7021 -9159 7081 -8847
rect 6623 -9219 6633 -9169
rect 6553 -9289 6633 -9219
rect 6553 -9349 6563 -9289
rect 6623 -9349 6633 -9289
rect 7011 -9219 7021 -9169
rect 7477 -9159 7537 -8847
rect 7081 -9219 7091 -9169
rect 7011 -9289 7091 -9219
rect 7011 -9349 7021 -9289
rect 7081 -9349 7091 -9289
rect 7467 -9219 7477 -9169
rect 7933 -9159 7993 -8847
rect 7537 -9219 7547 -9169
rect 7467 -9289 7547 -9219
rect 7467 -9349 7477 -9289
rect 7537 -9349 7547 -9289
rect 7923 -9219 7933 -9169
rect 8407 -9159 8467 -8847
rect 7993 -9219 8003 -9169
rect 7923 -9289 8003 -9219
rect 7923 -9349 7933 -9289
rect 7993 -9349 8003 -9289
rect 8397 -9219 8407 -9169
rect 8863 -9159 8923 -8847
rect 8467 -9219 8477 -9169
rect 8397 -9289 8477 -9219
rect 8397 -9349 8407 -9289
rect 8467 -9349 8477 -9289
rect 8853 -9219 8863 -9169
rect 9321 -9159 9381 -8847
rect 8923 -9219 8933 -9169
rect 8853 -9289 8933 -9219
rect 8853 -9349 8863 -9289
rect 8923 -9349 8933 -9289
rect 9311 -9219 9321 -9169
rect 9777 -9159 9837 -8847
rect 9381 -9219 9391 -9169
rect 9311 -9289 9391 -9219
rect 9311 -9349 9321 -9289
rect 9381 -9349 9391 -9289
rect 9767 -9219 9777 -9169
rect 10233 -9159 10293 -8847
rect 9837 -9219 9847 -9169
rect 9767 -9289 9847 -9219
rect 9767 -9349 9777 -9289
rect 9837 -9349 9847 -9289
rect 10223 -9219 10233 -9169
rect 10691 -9159 10751 -8847
rect 10293 -9219 10303 -9169
rect 10223 -9289 10303 -9219
rect 10223 -9349 10233 -9289
rect 10293 -9349 10303 -9289
rect 10681 -9219 10691 -9169
rect 11147 -9159 11207 -8847
rect 10751 -9219 10761 -9169
rect 10681 -9289 10761 -9219
rect 10681 -9349 10691 -9289
rect 10751 -9349 10761 -9289
rect 11137 -9219 11147 -9169
rect 11603 -9159 11663 -8847
rect 11207 -9219 11217 -9169
rect 11137 -9289 11217 -9219
rect 11137 -9349 11147 -9289
rect 11207 -9349 11217 -9289
rect 11593 -9219 11603 -9169
rect 12061 -9159 12121 -8847
rect 11663 -9219 11673 -9169
rect 11593 -9289 11673 -9219
rect 11593 -9349 11603 -9289
rect 11663 -9349 11673 -9289
rect 12051 -9219 12061 -9169
rect 12517 -9159 12577 -8847
rect 12121 -9219 12131 -9169
rect 12051 -9289 12131 -9219
rect 12051 -9349 12061 -9289
rect 12121 -9349 12131 -9289
rect 12507 -9219 12517 -9169
rect 12973 -9159 13033 -8847
rect 12577 -9219 12587 -9169
rect 12507 -9289 12587 -9219
rect 12507 -9349 12517 -9289
rect 12577 -9349 12587 -9289
rect 12963 -9219 12973 -9169
rect 13431 -9159 13491 -8847
rect 13033 -9219 13043 -9169
rect 12963 -9289 13043 -9219
rect 12963 -9349 12973 -9289
rect 13033 -9349 13043 -9289
rect 13421 -9219 13431 -9169
rect 13887 -9159 13947 -8847
rect 13491 -9219 13501 -9169
rect 13421 -9289 13501 -9219
rect 13421 -9349 13431 -9289
rect 13491 -9349 13501 -9289
rect 13877 -9219 13887 -9169
rect 14343 -9159 14403 -8847
rect 13947 -9219 13957 -9169
rect 13877 -9289 13957 -9219
rect 13877 -9349 13887 -9289
rect 13947 -9349 13957 -9289
rect 14333 -9219 14343 -9169
rect 14801 -9159 14861 -8847
rect 14403 -9219 14413 -9169
rect 14333 -9289 14413 -9219
rect 14333 -9349 14343 -9289
rect 14403 -9349 14413 -9289
rect 14791 -9219 14801 -9169
rect 15257 -9159 15317 -8847
rect 14861 -9219 14871 -9169
rect 14791 -9289 14871 -9219
rect 14791 -9349 14801 -9289
rect 14861 -9349 14871 -9289
rect 15247 -9219 15257 -9169
rect 15317 -9219 15327 -9169
rect 15247 -9289 15327 -9219
rect 15247 -9349 15257 -9289
rect 15317 -9349 15327 -9289
rect 171 -9651 231 -9349
rect 161 -9711 171 -9661
rect 627 -9651 687 -9349
rect 231 -9711 241 -9661
rect 161 -9781 241 -9711
rect 161 -9841 171 -9781
rect 231 -9841 241 -9781
rect 617 -9711 627 -9661
rect 1083 -9651 1143 -9349
rect 687 -9711 697 -9661
rect 617 -9781 697 -9711
rect 617 -9841 627 -9781
rect 687 -9841 697 -9781
rect 1073 -9711 1083 -9661
rect 1541 -9651 1601 -9349
rect 1143 -9711 1153 -9661
rect 1073 -9781 1153 -9711
rect 1073 -9841 1083 -9781
rect 1143 -9841 1153 -9781
rect 1531 -9711 1541 -9661
rect 1997 -9651 2057 -9349
rect 1601 -9711 1611 -9661
rect 1531 -9781 1611 -9711
rect 1531 -9841 1541 -9781
rect 1601 -9841 1611 -9781
rect 1987 -9711 1997 -9661
rect 2453 -9651 2513 -9349
rect 2057 -9711 2067 -9661
rect 1987 -9781 2067 -9711
rect 1987 -9841 1997 -9781
rect 2057 -9841 2067 -9781
rect 2443 -9711 2453 -9661
rect 2911 -9651 2971 -9349
rect 2513 -9711 2523 -9661
rect 2443 -9781 2523 -9711
rect 2443 -9841 2453 -9781
rect 2513 -9841 2523 -9781
rect 2901 -9711 2911 -9661
rect 3367 -9651 3427 -9349
rect 2971 -9711 2981 -9661
rect 2901 -9781 2981 -9711
rect 2901 -9841 2911 -9781
rect 2971 -9841 2981 -9781
rect 3357 -9711 3367 -9661
rect 3823 -9651 3883 -9349
rect 3427 -9711 3437 -9661
rect 3357 -9781 3437 -9711
rect 3357 -9841 3367 -9781
rect 3427 -9841 3437 -9781
rect 3813 -9711 3823 -9661
rect 4281 -9651 4341 -9349
rect 3883 -9711 3893 -9661
rect 3813 -9781 3893 -9711
rect 3813 -9841 3823 -9781
rect 3883 -9841 3893 -9781
rect 4271 -9711 4281 -9661
rect 4737 -9651 4797 -9349
rect 4341 -9711 4351 -9661
rect 4271 -9781 4351 -9711
rect 4271 -9841 4281 -9781
rect 4341 -9841 4351 -9781
rect 4727 -9711 4737 -9661
rect 5193 -9651 5253 -9349
rect 4797 -9711 4807 -9661
rect 4727 -9781 4807 -9711
rect 4727 -9841 4737 -9781
rect 4797 -9841 4807 -9781
rect 5183 -9711 5193 -9661
rect 5651 -9651 5711 -9349
rect 5253 -9711 5263 -9661
rect 5183 -9781 5263 -9711
rect 5183 -9841 5193 -9781
rect 5253 -9841 5263 -9781
rect 5641 -9711 5651 -9661
rect 6107 -9651 6167 -9349
rect 5711 -9711 5721 -9661
rect 5641 -9781 5721 -9711
rect 5641 -9841 5651 -9781
rect 5711 -9841 5721 -9781
rect 6097 -9711 6107 -9661
rect 6563 -9651 6623 -9349
rect 6167 -9711 6177 -9661
rect 6097 -9781 6177 -9711
rect 6097 -9841 6107 -9781
rect 6167 -9841 6177 -9781
rect 6553 -9711 6563 -9661
rect 7021 -9651 7081 -9349
rect 6623 -9711 6633 -9661
rect 6553 -9781 6633 -9711
rect 6553 -9841 6563 -9781
rect 6623 -9841 6633 -9781
rect 7011 -9711 7021 -9661
rect 7477 -9651 7537 -9349
rect 7081 -9711 7091 -9661
rect 7011 -9781 7091 -9711
rect 7011 -9841 7021 -9781
rect 7081 -9841 7091 -9781
rect 7467 -9711 7477 -9661
rect 7933 -9651 7993 -9349
rect 7537 -9711 7547 -9661
rect 7467 -9781 7547 -9711
rect 7467 -9841 7477 -9781
rect 7537 -9841 7547 -9781
rect 7923 -9711 7933 -9661
rect 8407 -9651 8467 -9349
rect 7993 -9711 8003 -9661
rect 7923 -9781 8003 -9711
rect 7923 -9841 7933 -9781
rect 7993 -9841 8003 -9781
rect 8397 -9711 8407 -9661
rect 8863 -9651 8923 -9349
rect 8467 -9711 8477 -9661
rect 8397 -9781 8477 -9711
rect 8397 -9841 8407 -9781
rect 8467 -9841 8477 -9781
rect 8853 -9711 8863 -9661
rect 9321 -9651 9381 -9349
rect 8923 -9711 8933 -9661
rect 8853 -9781 8933 -9711
rect 8853 -9841 8863 -9781
rect 8923 -9841 8933 -9781
rect 9311 -9711 9321 -9661
rect 9777 -9651 9837 -9349
rect 9381 -9711 9391 -9661
rect 9311 -9781 9391 -9711
rect 9311 -9841 9321 -9781
rect 9381 -9841 9391 -9781
rect 9767 -9711 9777 -9661
rect 10233 -9651 10293 -9349
rect 9837 -9711 9847 -9661
rect 9767 -9781 9847 -9711
rect 9767 -9841 9777 -9781
rect 9837 -9841 9847 -9781
rect 10223 -9711 10233 -9661
rect 10691 -9651 10751 -9349
rect 10293 -9711 10303 -9661
rect 10223 -9781 10303 -9711
rect 10223 -9841 10233 -9781
rect 10293 -9841 10303 -9781
rect 10681 -9711 10691 -9661
rect 11147 -9651 11207 -9349
rect 10751 -9711 10761 -9661
rect 10681 -9781 10761 -9711
rect 10681 -9841 10691 -9781
rect 10751 -9841 10761 -9781
rect 11137 -9711 11147 -9661
rect 11603 -9651 11663 -9349
rect 11207 -9711 11217 -9661
rect 11137 -9781 11217 -9711
rect 11137 -9841 11147 -9781
rect 11207 -9841 11217 -9781
rect 11593 -9711 11603 -9661
rect 12061 -9651 12121 -9349
rect 11663 -9711 11673 -9661
rect 11593 -9781 11673 -9711
rect 11593 -9841 11603 -9781
rect 11663 -9841 11673 -9781
rect 12051 -9711 12061 -9661
rect 12517 -9651 12577 -9349
rect 12121 -9711 12131 -9661
rect 12051 -9781 12131 -9711
rect 12051 -9841 12061 -9781
rect 12121 -9841 12131 -9781
rect 12507 -9711 12517 -9661
rect 12973 -9651 13033 -9349
rect 12577 -9711 12587 -9661
rect 12507 -9781 12587 -9711
rect 12507 -9841 12517 -9781
rect 12577 -9841 12587 -9781
rect 12963 -9711 12973 -9661
rect 13431 -9651 13491 -9349
rect 13033 -9711 13043 -9661
rect 12963 -9781 13043 -9711
rect 12963 -9841 12973 -9781
rect 13033 -9841 13043 -9781
rect 13421 -9711 13431 -9661
rect 13887 -9651 13947 -9349
rect 13491 -9711 13501 -9661
rect 13421 -9781 13501 -9711
rect 13421 -9841 13431 -9781
rect 13491 -9841 13501 -9781
rect 13877 -9711 13887 -9661
rect 14343 -9651 14403 -9349
rect 13947 -9711 13957 -9661
rect 13877 -9781 13957 -9711
rect 13877 -9841 13887 -9781
rect 13947 -9841 13957 -9781
rect 14333 -9711 14343 -9661
rect 14801 -9651 14861 -9349
rect 14403 -9711 14413 -9661
rect 14333 -9781 14413 -9711
rect 14333 -9841 14343 -9781
rect 14403 -9841 14413 -9781
rect 14791 -9711 14801 -9661
rect 15257 -9651 15317 -9349
rect 14861 -9711 14871 -9661
rect 14791 -9781 14871 -9711
rect 14791 -9841 14801 -9781
rect 14861 -9841 14871 -9781
rect 15247 -9711 15257 -9661
rect 15317 -9711 15327 -9661
rect 15247 -9781 15327 -9711
rect 15247 -9841 15257 -9781
rect 15317 -9841 15327 -9781
rect 171 -10167 231 -9841
rect 161 -10227 171 -10177
rect 627 -10167 687 -9841
rect 231 -10227 241 -10177
rect 161 -10297 241 -10227
rect 161 -10357 171 -10297
rect 231 -10357 241 -10297
rect 617 -10227 627 -10177
rect 1083 -10167 1143 -9841
rect 687 -10227 697 -10177
rect 617 -10297 697 -10227
rect 617 -10357 627 -10297
rect 687 -10357 697 -10297
rect 1073 -10227 1083 -10177
rect 1541 -10167 1601 -9841
rect 1143 -10227 1153 -10177
rect 1073 -10297 1153 -10227
rect 1073 -10357 1083 -10297
rect 1143 -10357 1153 -10297
rect 1531 -10227 1541 -10177
rect 1997 -10167 2057 -9841
rect 1601 -10227 1611 -10177
rect 1531 -10297 1611 -10227
rect 1531 -10357 1541 -10297
rect 1601 -10357 1611 -10297
rect 1987 -10227 1997 -10177
rect 2453 -10167 2513 -9841
rect 2057 -10227 2067 -10177
rect 1987 -10297 2067 -10227
rect 1987 -10357 1997 -10297
rect 2057 -10357 2067 -10297
rect 2443 -10227 2453 -10177
rect 2911 -10167 2971 -9841
rect 2513 -10227 2523 -10177
rect 2443 -10297 2523 -10227
rect 2443 -10357 2453 -10297
rect 2513 -10357 2523 -10297
rect 2901 -10227 2911 -10177
rect 3367 -10167 3427 -9841
rect 2971 -10227 2981 -10177
rect 2901 -10297 2981 -10227
rect 2901 -10357 2911 -10297
rect 2971 -10357 2981 -10297
rect 3357 -10227 3367 -10177
rect 3823 -10167 3883 -9841
rect 3427 -10227 3437 -10177
rect 3357 -10297 3437 -10227
rect 3357 -10357 3367 -10297
rect 3427 -10357 3437 -10297
rect 3813 -10227 3823 -10177
rect 4281 -10167 4341 -9841
rect 3883 -10227 3893 -10177
rect 3813 -10297 3893 -10227
rect 3813 -10357 3823 -10297
rect 3883 -10357 3893 -10297
rect 4271 -10227 4281 -10177
rect 4737 -10167 4797 -9841
rect 4341 -10227 4351 -10177
rect 4271 -10297 4351 -10227
rect 4271 -10357 4281 -10297
rect 4341 -10357 4351 -10297
rect 4727 -10227 4737 -10177
rect 5193 -10167 5253 -9841
rect 4797 -10227 4807 -10177
rect 4727 -10297 4807 -10227
rect 4727 -10357 4737 -10297
rect 4797 -10357 4807 -10297
rect 5183 -10227 5193 -10177
rect 5651 -10167 5711 -9841
rect 5253 -10227 5263 -10177
rect 5183 -10297 5263 -10227
rect 5183 -10357 5193 -10297
rect 5253 -10357 5263 -10297
rect 5641 -10227 5651 -10177
rect 6107 -10167 6167 -9841
rect 5711 -10227 5721 -10177
rect 5641 -10297 5721 -10227
rect 5641 -10357 5651 -10297
rect 5711 -10357 5721 -10297
rect 6097 -10227 6107 -10177
rect 6563 -10167 6623 -9841
rect 6167 -10227 6177 -10177
rect 6097 -10297 6177 -10227
rect 6097 -10357 6107 -10297
rect 6167 -10357 6177 -10297
rect 6553 -10227 6563 -10177
rect 7021 -10167 7081 -9841
rect 6623 -10227 6633 -10177
rect 6553 -10297 6633 -10227
rect 6553 -10357 6563 -10297
rect 6623 -10357 6633 -10297
rect 7011 -10227 7021 -10177
rect 7477 -10167 7537 -9841
rect 7081 -10227 7091 -10177
rect 7011 -10297 7091 -10227
rect 7011 -10357 7021 -10297
rect 7081 -10357 7091 -10297
rect 7467 -10227 7477 -10177
rect 7933 -10167 7993 -9841
rect 7537 -10227 7547 -10177
rect 7467 -10297 7547 -10227
rect 7467 -10357 7477 -10297
rect 7537 -10357 7547 -10297
rect 7923 -10227 7933 -10177
rect 8407 -10167 8467 -9841
rect 7993 -10227 8003 -10177
rect 7923 -10297 8003 -10227
rect 7923 -10357 7933 -10297
rect 7993 -10357 8003 -10297
rect 8397 -10227 8407 -10177
rect 8863 -10167 8923 -9841
rect 8467 -10227 8477 -10177
rect 8397 -10297 8477 -10227
rect 8397 -10357 8407 -10297
rect 8467 -10357 8477 -10297
rect 8853 -10227 8863 -10177
rect 9321 -10167 9381 -9841
rect 8923 -10227 8933 -10177
rect 8853 -10297 8933 -10227
rect 8853 -10357 8863 -10297
rect 8923 -10357 8933 -10297
rect 9311 -10227 9321 -10177
rect 9777 -10167 9837 -9841
rect 9381 -10227 9391 -10177
rect 9311 -10297 9391 -10227
rect 9311 -10357 9321 -10297
rect 9381 -10357 9391 -10297
rect 9767 -10227 9777 -10177
rect 10233 -10167 10293 -9841
rect 9837 -10227 9847 -10177
rect 9767 -10297 9847 -10227
rect 9767 -10357 9777 -10297
rect 9837 -10357 9847 -10297
rect 10223 -10227 10233 -10177
rect 10691 -10167 10751 -9841
rect 10293 -10227 10303 -10177
rect 10223 -10297 10303 -10227
rect 10223 -10357 10233 -10297
rect 10293 -10357 10303 -10297
rect 10681 -10227 10691 -10177
rect 11147 -10167 11207 -9841
rect 10751 -10227 10761 -10177
rect 10681 -10297 10761 -10227
rect 10681 -10357 10691 -10297
rect 10751 -10357 10761 -10297
rect 11137 -10227 11147 -10177
rect 11603 -10167 11663 -9841
rect 11207 -10227 11217 -10177
rect 11137 -10297 11217 -10227
rect 11137 -10357 11147 -10297
rect 11207 -10357 11217 -10297
rect 11593 -10227 11603 -10177
rect 12061 -10167 12121 -9841
rect 11663 -10227 11673 -10177
rect 11593 -10297 11673 -10227
rect 11593 -10357 11603 -10297
rect 11663 -10357 11673 -10297
rect 12051 -10227 12061 -10177
rect 12517 -10167 12577 -9841
rect 12121 -10227 12131 -10177
rect 12051 -10297 12131 -10227
rect 12051 -10357 12061 -10297
rect 12121 -10357 12131 -10297
rect 12507 -10227 12517 -10177
rect 12973 -10167 13033 -9841
rect 12577 -10227 12587 -10177
rect 12507 -10297 12587 -10227
rect 12507 -10357 12517 -10297
rect 12577 -10357 12587 -10297
rect 12963 -10227 12973 -10177
rect 13431 -10167 13491 -9841
rect 13033 -10227 13043 -10177
rect 12963 -10297 13043 -10227
rect 12963 -10357 12973 -10297
rect 13033 -10357 13043 -10297
rect 13421 -10227 13431 -10177
rect 13887 -10167 13947 -9841
rect 13491 -10227 13501 -10177
rect 13421 -10297 13501 -10227
rect 13421 -10357 13431 -10297
rect 13491 -10357 13501 -10297
rect 13877 -10227 13887 -10177
rect 14343 -10167 14403 -9841
rect 13947 -10227 13957 -10177
rect 13877 -10297 13957 -10227
rect 13877 -10357 13887 -10297
rect 13947 -10357 13957 -10297
rect 14333 -10227 14343 -10177
rect 14801 -10167 14861 -9841
rect 14403 -10227 14413 -10177
rect 14333 -10297 14413 -10227
rect 14333 -10357 14343 -10297
rect 14403 -10357 14413 -10297
rect 14791 -10227 14801 -10177
rect 15257 -10167 15317 -9841
rect 14861 -10227 14871 -10177
rect 14791 -10297 14871 -10227
rect 14791 -10357 14801 -10297
rect 14861 -10357 14871 -10297
rect 15247 -10227 15257 -10177
rect 15317 -10227 15327 -10177
rect 15247 -10297 15327 -10227
rect 15247 -10357 15257 -10297
rect 15317 -10357 15327 -10297
rect 171 -10669 231 -10357
rect 161 -10729 171 -10679
rect 627 -10669 687 -10357
rect 231 -10729 241 -10679
rect 161 -10799 241 -10729
rect 161 -10859 171 -10799
rect 231 -10859 241 -10799
rect 617 -10729 627 -10679
rect 1083 -10669 1143 -10357
rect 687 -10729 697 -10679
rect 617 -10799 697 -10729
rect 617 -10859 627 -10799
rect 687 -10859 697 -10799
rect 1073 -10729 1083 -10679
rect 1541 -10669 1601 -10357
rect 1143 -10729 1153 -10679
rect 1073 -10799 1153 -10729
rect 1073 -10859 1083 -10799
rect 1143 -10859 1153 -10799
rect 1531 -10729 1541 -10679
rect 1997 -10669 2057 -10357
rect 1601 -10729 1611 -10679
rect 1531 -10799 1611 -10729
rect 1531 -10859 1541 -10799
rect 1601 -10859 1611 -10799
rect 1987 -10729 1997 -10679
rect 2453 -10669 2513 -10357
rect 2057 -10729 2067 -10679
rect 1987 -10799 2067 -10729
rect 1987 -10859 1997 -10799
rect 2057 -10859 2067 -10799
rect 2443 -10729 2453 -10679
rect 2911 -10669 2971 -10357
rect 2513 -10729 2523 -10679
rect 2443 -10799 2523 -10729
rect 2443 -10859 2453 -10799
rect 2513 -10859 2523 -10799
rect 2901 -10729 2911 -10679
rect 3367 -10669 3427 -10357
rect 2971 -10729 2981 -10679
rect 2901 -10799 2981 -10729
rect 2901 -10859 2911 -10799
rect 2971 -10859 2981 -10799
rect 3357 -10729 3367 -10679
rect 3823 -10669 3883 -10357
rect 3427 -10729 3437 -10679
rect 3357 -10799 3437 -10729
rect 3357 -10859 3367 -10799
rect 3427 -10859 3437 -10799
rect 3813 -10729 3823 -10679
rect 4281 -10669 4341 -10357
rect 3883 -10729 3893 -10679
rect 3813 -10799 3893 -10729
rect 3813 -10859 3823 -10799
rect 3883 -10859 3893 -10799
rect 4271 -10729 4281 -10679
rect 4737 -10669 4797 -10357
rect 4341 -10729 4351 -10679
rect 4271 -10799 4351 -10729
rect 4271 -10859 4281 -10799
rect 4341 -10859 4351 -10799
rect 4727 -10729 4737 -10679
rect 5193 -10669 5253 -10357
rect 4797 -10729 4807 -10679
rect 4727 -10799 4807 -10729
rect 4727 -10859 4737 -10799
rect 4797 -10859 4807 -10799
rect 5183 -10729 5193 -10679
rect 5651 -10669 5711 -10357
rect 5253 -10729 5263 -10679
rect 5183 -10799 5263 -10729
rect 5183 -10859 5193 -10799
rect 5253 -10859 5263 -10799
rect 5641 -10729 5651 -10679
rect 6107 -10669 6167 -10357
rect 5711 -10729 5721 -10679
rect 5641 -10799 5721 -10729
rect 5641 -10859 5651 -10799
rect 5711 -10859 5721 -10799
rect 6097 -10729 6107 -10679
rect 6563 -10669 6623 -10357
rect 6167 -10729 6177 -10679
rect 6097 -10799 6177 -10729
rect 6097 -10859 6107 -10799
rect 6167 -10859 6177 -10799
rect 6553 -10729 6563 -10679
rect 7021 -10669 7081 -10357
rect 6623 -10729 6633 -10679
rect 6553 -10799 6633 -10729
rect 6553 -10859 6563 -10799
rect 6623 -10859 6633 -10799
rect 7011 -10729 7021 -10679
rect 7477 -10669 7537 -10357
rect 7081 -10729 7091 -10679
rect 7011 -10799 7091 -10729
rect 7011 -10859 7021 -10799
rect 7081 -10859 7091 -10799
rect 7467 -10729 7477 -10679
rect 7933 -10669 7993 -10357
rect 7537 -10729 7547 -10679
rect 7467 -10799 7547 -10729
rect 7467 -10859 7477 -10799
rect 7537 -10859 7547 -10799
rect 7923 -10729 7933 -10679
rect 8407 -10669 8467 -10357
rect 7993 -10729 8003 -10679
rect 7923 -10799 8003 -10729
rect 7923 -10859 7933 -10799
rect 7993 -10859 8003 -10799
rect 8397 -10729 8407 -10679
rect 8863 -10669 8923 -10357
rect 8467 -10729 8477 -10679
rect 8397 -10799 8477 -10729
rect 8397 -10859 8407 -10799
rect 8467 -10859 8477 -10799
rect 8853 -10729 8863 -10679
rect 9321 -10669 9381 -10357
rect 8923 -10729 8933 -10679
rect 8853 -10799 8933 -10729
rect 8853 -10859 8863 -10799
rect 8923 -10859 8933 -10799
rect 9311 -10729 9321 -10679
rect 9777 -10669 9837 -10357
rect 9381 -10729 9391 -10679
rect 9311 -10799 9391 -10729
rect 9311 -10859 9321 -10799
rect 9381 -10859 9391 -10799
rect 9767 -10729 9777 -10679
rect 10233 -10669 10293 -10357
rect 9837 -10729 9847 -10679
rect 9767 -10799 9847 -10729
rect 9767 -10859 9777 -10799
rect 9837 -10859 9847 -10799
rect 10223 -10729 10233 -10679
rect 10691 -10669 10751 -10357
rect 10293 -10729 10303 -10679
rect 10223 -10799 10303 -10729
rect 10223 -10859 10233 -10799
rect 10293 -10859 10303 -10799
rect 10681 -10729 10691 -10679
rect 11147 -10669 11207 -10357
rect 10751 -10729 10761 -10679
rect 10681 -10799 10761 -10729
rect 10681 -10859 10691 -10799
rect 10751 -10859 10761 -10799
rect 11137 -10729 11147 -10679
rect 11603 -10669 11663 -10357
rect 11207 -10729 11217 -10679
rect 11137 -10799 11217 -10729
rect 11137 -10859 11147 -10799
rect 11207 -10859 11217 -10799
rect 11593 -10729 11603 -10679
rect 12061 -10669 12121 -10357
rect 11663 -10729 11673 -10679
rect 11593 -10799 11673 -10729
rect 11593 -10859 11603 -10799
rect 11663 -10859 11673 -10799
rect 12051 -10729 12061 -10679
rect 12517 -10669 12577 -10357
rect 12121 -10729 12131 -10679
rect 12051 -10799 12131 -10729
rect 12051 -10859 12061 -10799
rect 12121 -10859 12131 -10799
rect 12507 -10729 12517 -10679
rect 12973 -10669 13033 -10357
rect 12577 -10729 12587 -10679
rect 12507 -10799 12587 -10729
rect 12507 -10859 12517 -10799
rect 12577 -10859 12587 -10799
rect 12963 -10729 12973 -10679
rect 13431 -10669 13491 -10357
rect 13033 -10729 13043 -10679
rect 12963 -10799 13043 -10729
rect 12963 -10859 12973 -10799
rect 13033 -10859 13043 -10799
rect 13421 -10729 13431 -10679
rect 13887 -10669 13947 -10357
rect 13491 -10729 13501 -10679
rect 13421 -10799 13501 -10729
rect 13421 -10859 13431 -10799
rect 13491 -10859 13501 -10799
rect 13877 -10729 13887 -10679
rect 14343 -10669 14403 -10357
rect 13947 -10729 13957 -10679
rect 13877 -10799 13957 -10729
rect 13877 -10859 13887 -10799
rect 13947 -10859 13957 -10799
rect 14333 -10729 14343 -10679
rect 14801 -10669 14861 -10357
rect 14403 -10729 14413 -10679
rect 14333 -10799 14413 -10729
rect 14333 -10859 14343 -10799
rect 14403 -10859 14413 -10799
rect 14791 -10729 14801 -10679
rect 15257 -10669 15317 -10357
rect 14861 -10729 14871 -10679
rect 14791 -10799 14871 -10729
rect 14791 -10859 14801 -10799
rect 14861 -10859 14871 -10799
rect 15247 -10729 15257 -10679
rect 15317 -10729 15327 -10679
rect 15247 -10799 15327 -10729
rect 15247 -10859 15257 -10799
rect 15317 -10859 15327 -10799
rect 171 -11161 231 -10859
rect 161 -11221 171 -11171
rect 627 -11161 687 -10859
rect 231 -11221 241 -11171
rect 161 -11291 241 -11221
rect 161 -11351 171 -11291
rect 231 -11351 241 -11291
rect 617 -11221 627 -11171
rect 1083 -11161 1143 -10859
rect 687 -11221 697 -11171
rect 617 -11291 697 -11221
rect 617 -11351 627 -11291
rect 687 -11351 697 -11291
rect 1073 -11221 1083 -11171
rect 1541 -11161 1601 -10859
rect 1143 -11221 1153 -11171
rect 1073 -11291 1153 -11221
rect 1073 -11351 1083 -11291
rect 1143 -11351 1153 -11291
rect 1531 -11221 1541 -11171
rect 1997 -11161 2057 -10859
rect 1601 -11221 1611 -11171
rect 1531 -11291 1611 -11221
rect 1531 -11351 1541 -11291
rect 1601 -11351 1611 -11291
rect 1987 -11221 1997 -11171
rect 2453 -11161 2513 -10859
rect 2057 -11221 2067 -11171
rect 1987 -11291 2067 -11221
rect 1987 -11351 1997 -11291
rect 2057 -11351 2067 -11291
rect 2443 -11221 2453 -11171
rect 2911 -11161 2971 -10859
rect 2513 -11221 2523 -11171
rect 2443 -11291 2523 -11221
rect 2443 -11351 2453 -11291
rect 2513 -11351 2523 -11291
rect 2901 -11221 2911 -11171
rect 3367 -11161 3427 -10859
rect 2971 -11221 2981 -11171
rect 2901 -11291 2981 -11221
rect 2901 -11351 2911 -11291
rect 2971 -11351 2981 -11291
rect 3357 -11221 3367 -11171
rect 3823 -11161 3883 -10859
rect 3427 -11221 3437 -11171
rect 3357 -11291 3437 -11221
rect 3357 -11351 3367 -11291
rect 3427 -11351 3437 -11291
rect 3813 -11221 3823 -11171
rect 4281 -11161 4341 -10859
rect 3883 -11221 3893 -11171
rect 3813 -11291 3893 -11221
rect 3813 -11351 3823 -11291
rect 3883 -11351 3893 -11291
rect 4271 -11221 4281 -11171
rect 4737 -11161 4797 -10859
rect 4341 -11221 4351 -11171
rect 4271 -11291 4351 -11221
rect 4271 -11351 4281 -11291
rect 4341 -11351 4351 -11291
rect 4727 -11221 4737 -11171
rect 5193 -11161 5253 -10859
rect 4797 -11221 4807 -11171
rect 4727 -11291 4807 -11221
rect 4727 -11351 4737 -11291
rect 4797 -11351 4807 -11291
rect 5183 -11221 5193 -11171
rect 5651 -11161 5711 -10859
rect 5253 -11221 5263 -11171
rect 5183 -11291 5263 -11221
rect 5183 -11351 5193 -11291
rect 5253 -11351 5263 -11291
rect 5641 -11221 5651 -11171
rect 6107 -11161 6167 -10859
rect 5711 -11221 5721 -11171
rect 5641 -11291 5721 -11221
rect 5641 -11351 5651 -11291
rect 5711 -11351 5721 -11291
rect 6097 -11221 6107 -11171
rect 6563 -11161 6623 -10859
rect 6167 -11221 6177 -11171
rect 6097 -11291 6177 -11221
rect 6097 -11351 6107 -11291
rect 6167 -11351 6177 -11291
rect 6553 -11221 6563 -11171
rect 7021 -11161 7081 -10859
rect 6623 -11221 6633 -11171
rect 6553 -11291 6633 -11221
rect 6553 -11351 6563 -11291
rect 6623 -11351 6633 -11291
rect 7011 -11221 7021 -11171
rect 7477 -11161 7537 -10859
rect 7081 -11221 7091 -11171
rect 7011 -11291 7091 -11221
rect 7011 -11351 7021 -11291
rect 7081 -11351 7091 -11291
rect 7467 -11221 7477 -11171
rect 7933 -11161 7993 -10859
rect 7537 -11221 7547 -11171
rect 7467 -11291 7547 -11221
rect 7467 -11351 7477 -11291
rect 7537 -11351 7547 -11291
rect 7923 -11221 7933 -11171
rect 8407 -11161 8467 -10859
rect 7993 -11221 8003 -11171
rect 7923 -11291 8003 -11221
rect 7923 -11351 7933 -11291
rect 7993 -11351 8003 -11291
rect 8397 -11221 8407 -11171
rect 8863 -11161 8923 -10859
rect 8467 -11221 8477 -11171
rect 8397 -11291 8477 -11221
rect 8397 -11351 8407 -11291
rect 8467 -11351 8477 -11291
rect 8853 -11221 8863 -11171
rect 9321 -11161 9381 -10859
rect 8923 -11221 8933 -11171
rect 8853 -11291 8933 -11221
rect 8853 -11351 8863 -11291
rect 8923 -11351 8933 -11291
rect 9311 -11221 9321 -11171
rect 9777 -11161 9837 -10859
rect 9381 -11221 9391 -11171
rect 9311 -11291 9391 -11221
rect 9311 -11351 9321 -11291
rect 9381 -11351 9391 -11291
rect 9767 -11221 9777 -11171
rect 10233 -11161 10293 -10859
rect 9837 -11221 9847 -11171
rect 9767 -11291 9847 -11221
rect 9767 -11351 9777 -11291
rect 9837 -11351 9847 -11291
rect 10223 -11221 10233 -11171
rect 10691 -11161 10751 -10859
rect 10293 -11221 10303 -11171
rect 10223 -11291 10303 -11221
rect 10223 -11351 10233 -11291
rect 10293 -11351 10303 -11291
rect 10681 -11221 10691 -11171
rect 11147 -11161 11207 -10859
rect 10751 -11221 10761 -11171
rect 10681 -11291 10761 -11221
rect 10681 -11351 10691 -11291
rect 10751 -11351 10761 -11291
rect 11137 -11221 11147 -11171
rect 11603 -11161 11663 -10859
rect 11207 -11221 11217 -11171
rect 11137 -11291 11217 -11221
rect 11137 -11351 11147 -11291
rect 11207 -11351 11217 -11291
rect 11593 -11221 11603 -11171
rect 12061 -11161 12121 -10859
rect 11663 -11221 11673 -11171
rect 11593 -11291 11673 -11221
rect 11593 -11351 11603 -11291
rect 11663 -11351 11673 -11291
rect 12051 -11221 12061 -11171
rect 12517 -11161 12577 -10859
rect 12121 -11221 12131 -11171
rect 12051 -11291 12131 -11221
rect 12051 -11351 12061 -11291
rect 12121 -11351 12131 -11291
rect 12507 -11221 12517 -11171
rect 12973 -11161 13033 -10859
rect 12577 -11221 12587 -11171
rect 12507 -11291 12587 -11221
rect 12507 -11351 12517 -11291
rect 12577 -11351 12587 -11291
rect 12963 -11221 12973 -11171
rect 13431 -11161 13491 -10859
rect 13033 -11221 13043 -11171
rect 12963 -11291 13043 -11221
rect 12963 -11351 12973 -11291
rect 13033 -11351 13043 -11291
rect 13421 -11221 13431 -11171
rect 13887 -11161 13947 -10859
rect 13491 -11221 13501 -11171
rect 13421 -11291 13501 -11221
rect 13421 -11351 13431 -11291
rect 13491 -11351 13501 -11291
rect 13877 -11221 13887 -11171
rect 14343 -11161 14403 -10859
rect 13947 -11221 13957 -11171
rect 13877 -11291 13957 -11221
rect 13877 -11351 13887 -11291
rect 13947 -11351 13957 -11291
rect 14333 -11221 14343 -11171
rect 14801 -11161 14861 -10859
rect 14403 -11221 14413 -11171
rect 14333 -11291 14413 -11221
rect 14333 -11351 14343 -11291
rect 14403 -11351 14413 -11291
rect 14791 -11221 14801 -11171
rect 15257 -11161 15317 -10859
rect 14861 -11221 14871 -11171
rect 14791 -11291 14871 -11221
rect 14791 -11351 14801 -11291
rect 14861 -11351 14871 -11291
rect 15247 -11221 15257 -11171
rect 15317 -11221 15327 -11171
rect 15247 -11291 15327 -11221
rect 15247 -11351 15257 -11291
rect 15317 -11351 15327 -11291
rect 171 -11489 231 -11351
rect 627 -11489 687 -11351
rect 1083 -11489 1143 -11351
rect 1541 -11489 1601 -11351
rect 1997 -11489 2057 -11351
rect 2453 -11489 2513 -11351
rect 2911 -11489 2971 -11351
rect 3367 -11489 3427 -11351
rect 3823 -11489 3883 -11351
rect 4281 -11489 4341 -11351
rect 4737 -11489 4797 -11351
rect 5193 -11489 5253 -11351
rect 5651 -11489 5711 -11351
rect 6107 -11489 6167 -11351
rect 6563 -11489 6623 -11351
rect 7021 -11489 7081 -11351
rect 7477 -11489 7537 -11351
rect 7933 -11489 7993 -11351
rect 8407 -11489 8467 -11351
rect 8863 -11489 8923 -11351
rect 9321 -11489 9381 -11351
rect 9777 -11489 9837 -11351
rect 10233 -11489 10293 -11351
rect 10691 -11489 10751 -11351
rect 11147 -11489 11207 -11351
rect 11603 -11489 11663 -11351
rect 12061 -11489 12121 -11351
rect 12517 -11489 12577 -11351
rect 12973 -11489 13033 -11351
rect 13431 -11489 13491 -11351
rect 13887 -11489 13947 -11351
rect 14343 -11489 14403 -11351
rect 14801 -11489 14861 -11351
rect 15257 -11489 15317 -11351
rect 170 -11491 231 -11489
rect 626 -11491 687 -11489
rect 1082 -11491 1143 -11489
rect 1540 -11491 1601 -11489
rect 1996 -11491 2057 -11489
rect 2452 -11491 2513 -11489
rect 2910 -11491 2971 -11489
rect 3366 -11491 3427 -11489
rect 3822 -11491 3883 -11489
rect 4280 -11491 4341 -11489
rect 4736 -11491 4797 -11489
rect 5192 -11491 5253 -11489
rect 5650 -11491 5711 -11489
rect 6106 -11491 6167 -11489
rect 6562 -11491 6623 -11489
rect 7020 -11491 7081 -11489
rect 7476 -11491 7537 -11489
rect 7932 -11491 7993 -11489
rect 8406 -11491 8467 -11489
rect 8862 -11491 8923 -11489
rect 9320 -11491 9381 -11489
rect 9776 -11491 9837 -11489
rect 10232 -11491 10293 -11489
rect 10690 -11491 10751 -11489
rect 11146 -11491 11207 -11489
rect 11602 -11491 11663 -11489
rect 12060 -11491 12121 -11489
rect 12516 -11491 12577 -11489
rect 12972 -11491 13033 -11489
rect 13430 -11491 13491 -11489
rect 13886 -11491 13947 -11489
rect 14342 -11491 14403 -11489
rect 14800 -11491 14861 -11489
rect 15256 -11491 15317 -11489
rect 170 -11654 230 -11491
rect 160 -11714 170 -11664
rect 626 -11654 686 -11491
rect 230 -11714 240 -11664
rect 160 -11784 240 -11714
rect 160 -11844 170 -11784
rect 230 -11844 240 -11784
rect 616 -11714 626 -11664
rect 1082 -11654 1142 -11491
rect 686 -11714 696 -11664
rect 616 -11784 696 -11714
rect 616 -11844 626 -11784
rect 686 -11844 696 -11784
rect 1072 -11714 1082 -11664
rect 1540 -11654 1600 -11491
rect 1142 -11714 1152 -11664
rect 1072 -11784 1152 -11714
rect 1072 -11844 1082 -11784
rect 1142 -11844 1152 -11784
rect 1530 -11714 1540 -11664
rect 1996 -11654 2056 -11491
rect 1600 -11714 1610 -11664
rect 1530 -11784 1610 -11714
rect 1530 -11844 1540 -11784
rect 1600 -11844 1610 -11784
rect 1986 -11714 1996 -11664
rect 2452 -11654 2512 -11491
rect 2056 -11714 2066 -11664
rect 1986 -11784 2066 -11714
rect 1986 -11844 1996 -11784
rect 2056 -11844 2066 -11784
rect 2442 -11714 2452 -11664
rect 2910 -11654 2970 -11491
rect 2512 -11714 2522 -11664
rect 2442 -11784 2522 -11714
rect 2442 -11844 2452 -11784
rect 2512 -11844 2522 -11784
rect 2900 -11714 2910 -11664
rect 3366 -11654 3426 -11491
rect 2970 -11714 2980 -11664
rect 2900 -11784 2980 -11714
rect 2900 -11844 2910 -11784
rect 2970 -11844 2980 -11784
rect 3356 -11714 3366 -11664
rect 3822 -11654 3882 -11491
rect 3426 -11714 3436 -11664
rect 3356 -11784 3436 -11714
rect 3356 -11844 3366 -11784
rect 3426 -11844 3436 -11784
rect 3812 -11714 3822 -11664
rect 4280 -11654 4340 -11491
rect 3882 -11714 3892 -11664
rect 3812 -11784 3892 -11714
rect 3812 -11844 3822 -11784
rect 3882 -11844 3892 -11784
rect 4270 -11714 4280 -11664
rect 4736 -11654 4796 -11491
rect 4340 -11714 4350 -11664
rect 4270 -11784 4350 -11714
rect 4270 -11844 4280 -11784
rect 4340 -11844 4350 -11784
rect 4726 -11714 4736 -11664
rect 5192 -11654 5252 -11491
rect 4796 -11714 4806 -11664
rect 4726 -11784 4806 -11714
rect 4726 -11844 4736 -11784
rect 4796 -11844 4806 -11784
rect 5182 -11714 5192 -11664
rect 5650 -11654 5710 -11491
rect 5252 -11714 5262 -11664
rect 5182 -11784 5262 -11714
rect 5182 -11844 5192 -11784
rect 5252 -11844 5262 -11784
rect 5640 -11714 5650 -11664
rect 6106 -11654 6166 -11491
rect 5710 -11714 5720 -11664
rect 5640 -11784 5720 -11714
rect 5640 -11844 5650 -11784
rect 5710 -11844 5720 -11784
rect 6096 -11714 6106 -11664
rect 6562 -11654 6622 -11491
rect 6166 -11714 6176 -11664
rect 6096 -11784 6176 -11714
rect 6096 -11844 6106 -11784
rect 6166 -11844 6176 -11784
rect 6552 -11714 6562 -11664
rect 7020 -11654 7080 -11491
rect 6622 -11714 6632 -11664
rect 6552 -11784 6632 -11714
rect 6552 -11844 6562 -11784
rect 6622 -11844 6632 -11784
rect 7010 -11714 7020 -11664
rect 7476 -11654 7536 -11491
rect 7080 -11714 7090 -11664
rect 7010 -11784 7090 -11714
rect 7010 -11844 7020 -11784
rect 7080 -11844 7090 -11784
rect 7466 -11714 7476 -11664
rect 7932 -11654 7992 -11491
rect 7536 -11714 7546 -11664
rect 7466 -11784 7546 -11714
rect 7466 -11844 7476 -11784
rect 7536 -11844 7546 -11784
rect 7922 -11714 7932 -11664
rect 8406 -11654 8466 -11491
rect 7992 -11714 8002 -11664
rect 7922 -11784 8002 -11714
rect 7922 -11844 7932 -11784
rect 7992 -11844 8002 -11784
rect 8396 -11714 8406 -11664
rect 8862 -11654 8922 -11491
rect 8466 -11714 8476 -11664
rect 8396 -11784 8476 -11714
rect 8396 -11844 8406 -11784
rect 8466 -11844 8476 -11784
rect 8852 -11714 8862 -11664
rect 9320 -11654 9380 -11491
rect 8922 -11714 8932 -11664
rect 8852 -11784 8932 -11714
rect 8852 -11844 8862 -11784
rect 8922 -11844 8932 -11784
rect 9310 -11714 9320 -11664
rect 9776 -11654 9836 -11491
rect 9380 -11714 9390 -11664
rect 9310 -11784 9390 -11714
rect 9310 -11844 9320 -11784
rect 9380 -11844 9390 -11784
rect 9766 -11714 9776 -11664
rect 10232 -11654 10292 -11491
rect 9836 -11714 9846 -11664
rect 9766 -11784 9846 -11714
rect 9766 -11844 9776 -11784
rect 9836 -11844 9846 -11784
rect 10222 -11714 10232 -11664
rect 10690 -11654 10750 -11491
rect 10292 -11714 10302 -11664
rect 10222 -11784 10302 -11714
rect 10222 -11844 10232 -11784
rect 10292 -11844 10302 -11784
rect 10680 -11714 10690 -11664
rect 11146 -11654 11206 -11491
rect 10750 -11714 10760 -11664
rect 10680 -11784 10760 -11714
rect 10680 -11844 10690 -11784
rect 10750 -11844 10760 -11784
rect 11136 -11714 11146 -11664
rect 11602 -11654 11662 -11491
rect 11206 -11714 11216 -11664
rect 11136 -11784 11216 -11714
rect 11136 -11844 11146 -11784
rect 11206 -11844 11216 -11784
rect 11592 -11714 11602 -11664
rect 12060 -11654 12120 -11491
rect 11662 -11714 11672 -11664
rect 11592 -11784 11672 -11714
rect 11592 -11844 11602 -11784
rect 11662 -11844 11672 -11784
rect 12050 -11714 12060 -11664
rect 12516 -11654 12576 -11491
rect 12120 -11714 12130 -11664
rect 12050 -11784 12130 -11714
rect 12050 -11844 12060 -11784
rect 12120 -11844 12130 -11784
rect 12506 -11714 12516 -11664
rect 12972 -11654 13032 -11491
rect 12576 -11714 12586 -11664
rect 12506 -11784 12586 -11714
rect 12506 -11844 12516 -11784
rect 12576 -11844 12586 -11784
rect 12962 -11714 12972 -11664
rect 13430 -11654 13490 -11491
rect 13032 -11714 13042 -11664
rect 12962 -11784 13042 -11714
rect 12962 -11844 12972 -11784
rect 13032 -11844 13042 -11784
rect 13420 -11714 13430 -11664
rect 13886 -11654 13946 -11491
rect 13490 -11714 13500 -11664
rect 13420 -11784 13500 -11714
rect 13420 -11844 13430 -11784
rect 13490 -11844 13500 -11784
rect 13876 -11714 13886 -11664
rect 14342 -11654 14402 -11491
rect 13946 -11714 13956 -11664
rect 13876 -11784 13956 -11714
rect 13876 -11844 13886 -11784
rect 13946 -11844 13956 -11784
rect 14332 -11714 14342 -11664
rect 14800 -11654 14860 -11491
rect 14402 -11714 14412 -11664
rect 14332 -11784 14412 -11714
rect 14332 -11844 14342 -11784
rect 14402 -11844 14412 -11784
rect 14790 -11714 14800 -11664
rect 15256 -11654 15316 -11491
rect 14860 -11714 14870 -11664
rect 14790 -11784 14870 -11714
rect 14790 -11844 14800 -11784
rect 14860 -11844 14870 -11784
rect 15246 -11714 15256 -11664
rect 15316 -11714 15326 -11664
rect 15246 -11784 15326 -11714
rect 15246 -11844 15256 -11784
rect 15316 -11844 15326 -11784
rect 170 -12146 230 -11844
rect 160 -12206 170 -12156
rect 626 -12146 686 -11844
rect 230 -12206 240 -12156
rect 160 -12276 240 -12206
rect 160 -12336 170 -12276
rect 230 -12336 240 -12276
rect 616 -12206 626 -12156
rect 1082 -12146 1142 -11844
rect 686 -12206 696 -12156
rect 616 -12276 696 -12206
rect 616 -12336 626 -12276
rect 686 -12336 696 -12276
rect 1072 -12206 1082 -12156
rect 1540 -12146 1600 -11844
rect 1142 -12206 1152 -12156
rect 1072 -12276 1152 -12206
rect 1072 -12336 1082 -12276
rect 1142 -12336 1152 -12276
rect 1530 -12206 1540 -12156
rect 1996 -12146 2056 -11844
rect 1600 -12206 1610 -12156
rect 1530 -12276 1610 -12206
rect 1530 -12336 1540 -12276
rect 1600 -12336 1610 -12276
rect 1986 -12206 1996 -12156
rect 2452 -12146 2512 -11844
rect 2056 -12206 2066 -12156
rect 1986 -12276 2066 -12206
rect 1986 -12336 1996 -12276
rect 2056 -12336 2066 -12276
rect 2442 -12206 2452 -12156
rect 2910 -12146 2970 -11844
rect 2512 -12206 2522 -12156
rect 2442 -12276 2522 -12206
rect 2442 -12336 2452 -12276
rect 2512 -12336 2522 -12276
rect 2900 -12206 2910 -12156
rect 3366 -12146 3426 -11844
rect 2970 -12206 2980 -12156
rect 2900 -12276 2980 -12206
rect 2900 -12336 2910 -12276
rect 2970 -12336 2980 -12276
rect 3356 -12206 3366 -12156
rect 3822 -12146 3882 -11844
rect 3426 -12206 3436 -12156
rect 3356 -12276 3436 -12206
rect 3356 -12336 3366 -12276
rect 3426 -12336 3436 -12276
rect 3812 -12206 3822 -12156
rect 4280 -12146 4340 -11844
rect 3882 -12206 3892 -12156
rect 3812 -12276 3892 -12206
rect 3812 -12336 3822 -12276
rect 3882 -12336 3892 -12276
rect 4270 -12206 4280 -12156
rect 4736 -12146 4796 -11844
rect 4340 -12206 4350 -12156
rect 4270 -12276 4350 -12206
rect 4270 -12336 4280 -12276
rect 4340 -12336 4350 -12276
rect 4726 -12206 4736 -12156
rect 5192 -12146 5252 -11844
rect 4796 -12206 4806 -12156
rect 4726 -12276 4806 -12206
rect 4726 -12336 4736 -12276
rect 4796 -12336 4806 -12276
rect 5182 -12206 5192 -12156
rect 5650 -12146 5710 -11844
rect 5252 -12206 5262 -12156
rect 5182 -12276 5262 -12206
rect 5182 -12336 5192 -12276
rect 5252 -12336 5262 -12276
rect 5640 -12206 5650 -12156
rect 6106 -12146 6166 -11844
rect 5710 -12206 5720 -12156
rect 5640 -12276 5720 -12206
rect 5640 -12336 5650 -12276
rect 5710 -12336 5720 -12276
rect 6096 -12206 6106 -12156
rect 6562 -12146 6622 -11844
rect 6166 -12206 6176 -12156
rect 6096 -12276 6176 -12206
rect 6096 -12336 6106 -12276
rect 6166 -12336 6176 -12276
rect 6552 -12206 6562 -12156
rect 7020 -12146 7080 -11844
rect 6622 -12206 6632 -12156
rect 6552 -12276 6632 -12206
rect 6552 -12336 6562 -12276
rect 6622 -12336 6632 -12276
rect 7010 -12206 7020 -12156
rect 7476 -12146 7536 -11844
rect 7080 -12206 7090 -12156
rect 7010 -12276 7090 -12206
rect 7010 -12336 7020 -12276
rect 7080 -12336 7090 -12276
rect 7466 -12206 7476 -12156
rect 7932 -12146 7992 -11844
rect 7536 -12206 7546 -12156
rect 7466 -12276 7546 -12206
rect 7466 -12336 7476 -12276
rect 7536 -12336 7546 -12276
rect 7922 -12206 7932 -12156
rect 8406 -12146 8466 -11844
rect 7992 -12206 8002 -12156
rect 7922 -12276 8002 -12206
rect 7922 -12336 7932 -12276
rect 7992 -12336 8002 -12276
rect 8396 -12206 8406 -12156
rect 8862 -12146 8922 -11844
rect 8466 -12206 8476 -12156
rect 8396 -12276 8476 -12206
rect 8396 -12336 8406 -12276
rect 8466 -12336 8476 -12276
rect 8852 -12206 8862 -12156
rect 9320 -12146 9380 -11844
rect 8922 -12206 8932 -12156
rect 8852 -12276 8932 -12206
rect 8852 -12336 8862 -12276
rect 8922 -12336 8932 -12276
rect 9310 -12206 9320 -12156
rect 9776 -12146 9836 -11844
rect 9380 -12206 9390 -12156
rect 9310 -12276 9390 -12206
rect 9310 -12336 9320 -12276
rect 9380 -12336 9390 -12276
rect 9766 -12206 9776 -12156
rect 10232 -12146 10292 -11844
rect 9836 -12206 9846 -12156
rect 9766 -12276 9846 -12206
rect 9766 -12336 9776 -12276
rect 9836 -12336 9846 -12276
rect 10222 -12206 10232 -12156
rect 10690 -12146 10750 -11844
rect 10292 -12206 10302 -12156
rect 10222 -12276 10302 -12206
rect 10222 -12336 10232 -12276
rect 10292 -12336 10302 -12276
rect 10680 -12206 10690 -12156
rect 11146 -12146 11206 -11844
rect 10750 -12206 10760 -12156
rect 10680 -12276 10760 -12206
rect 10680 -12336 10690 -12276
rect 10750 -12336 10760 -12276
rect 11136 -12206 11146 -12156
rect 11602 -12146 11662 -11844
rect 11206 -12206 11216 -12156
rect 11136 -12276 11216 -12206
rect 11136 -12336 11146 -12276
rect 11206 -12336 11216 -12276
rect 11592 -12206 11602 -12156
rect 12060 -12146 12120 -11844
rect 11662 -12206 11672 -12156
rect 11592 -12276 11672 -12206
rect 11592 -12336 11602 -12276
rect 11662 -12336 11672 -12276
rect 12050 -12206 12060 -12156
rect 12516 -12146 12576 -11844
rect 12120 -12206 12130 -12156
rect 12050 -12276 12130 -12206
rect 12050 -12336 12060 -12276
rect 12120 -12336 12130 -12276
rect 12506 -12206 12516 -12156
rect 12972 -12146 13032 -11844
rect 12576 -12206 12586 -12156
rect 12506 -12276 12586 -12206
rect 12506 -12336 12516 -12276
rect 12576 -12336 12586 -12276
rect 12962 -12206 12972 -12156
rect 13430 -12146 13490 -11844
rect 13032 -12206 13042 -12156
rect 12962 -12276 13042 -12206
rect 12962 -12336 12972 -12276
rect 13032 -12336 13042 -12276
rect 13420 -12206 13430 -12156
rect 13886 -12146 13946 -11844
rect 13490 -12206 13500 -12156
rect 13420 -12276 13500 -12206
rect 13420 -12336 13430 -12276
rect 13490 -12336 13500 -12276
rect 13876 -12206 13886 -12156
rect 14342 -12146 14402 -11844
rect 13946 -12206 13956 -12156
rect 13876 -12276 13956 -12206
rect 13876 -12336 13886 -12276
rect 13946 -12336 13956 -12276
rect 14332 -12206 14342 -12156
rect 14800 -12146 14860 -11844
rect 14402 -12206 14412 -12156
rect 14332 -12276 14412 -12206
rect 14332 -12336 14342 -12276
rect 14402 -12336 14412 -12276
rect 14790 -12206 14800 -12156
rect 15256 -12146 15316 -11844
rect 14860 -12206 14870 -12156
rect 14790 -12276 14870 -12206
rect 14790 -12336 14800 -12276
rect 14860 -12336 14870 -12276
rect 15246 -12206 15256 -12156
rect 15316 -12206 15326 -12156
rect 15246 -12276 15326 -12206
rect 15246 -12336 15256 -12276
rect 15316 -12336 15326 -12276
rect 170 -12662 230 -12336
rect 160 -12722 170 -12672
rect 626 -12662 686 -12336
rect 230 -12722 240 -12672
rect 160 -12792 240 -12722
rect 160 -12852 170 -12792
rect 230 -12852 240 -12792
rect 616 -12722 626 -12672
rect 1082 -12662 1142 -12336
rect 686 -12722 696 -12672
rect 616 -12792 696 -12722
rect 616 -12852 626 -12792
rect 686 -12852 696 -12792
rect 1072 -12722 1082 -12672
rect 1540 -12662 1600 -12336
rect 1142 -12722 1152 -12672
rect 1072 -12792 1152 -12722
rect 1072 -12852 1082 -12792
rect 1142 -12852 1152 -12792
rect 1530 -12722 1540 -12672
rect 1996 -12662 2056 -12336
rect 1600 -12722 1610 -12672
rect 1530 -12792 1610 -12722
rect 1530 -12852 1540 -12792
rect 1600 -12852 1610 -12792
rect 1986 -12722 1996 -12672
rect 2452 -12662 2512 -12336
rect 2056 -12722 2066 -12672
rect 1986 -12792 2066 -12722
rect 1986 -12852 1996 -12792
rect 2056 -12852 2066 -12792
rect 2442 -12722 2452 -12672
rect 2910 -12662 2970 -12336
rect 2512 -12722 2522 -12672
rect 2442 -12792 2522 -12722
rect 2442 -12852 2452 -12792
rect 2512 -12852 2522 -12792
rect 2900 -12722 2910 -12672
rect 3366 -12662 3426 -12336
rect 2970 -12722 2980 -12672
rect 2900 -12792 2980 -12722
rect 2900 -12852 2910 -12792
rect 2970 -12852 2980 -12792
rect 3356 -12722 3366 -12672
rect 3822 -12662 3882 -12336
rect 3426 -12722 3436 -12672
rect 3356 -12792 3436 -12722
rect 3356 -12852 3366 -12792
rect 3426 -12852 3436 -12792
rect 3812 -12722 3822 -12672
rect 4280 -12662 4340 -12336
rect 3882 -12722 3892 -12672
rect 3812 -12792 3892 -12722
rect 3812 -12852 3822 -12792
rect 3882 -12852 3892 -12792
rect 4270 -12722 4280 -12672
rect 4736 -12662 4796 -12336
rect 4340 -12722 4350 -12672
rect 4270 -12792 4350 -12722
rect 4270 -12852 4280 -12792
rect 4340 -12852 4350 -12792
rect 4726 -12722 4736 -12672
rect 5192 -12662 5252 -12336
rect 4796 -12722 4806 -12672
rect 4726 -12792 4806 -12722
rect 4726 -12852 4736 -12792
rect 4796 -12852 4806 -12792
rect 5182 -12722 5192 -12672
rect 5650 -12662 5710 -12336
rect 5252 -12722 5262 -12672
rect 5182 -12792 5262 -12722
rect 5182 -12852 5192 -12792
rect 5252 -12852 5262 -12792
rect 5640 -12722 5650 -12672
rect 6106 -12662 6166 -12336
rect 5710 -12722 5720 -12672
rect 5640 -12792 5720 -12722
rect 5640 -12852 5650 -12792
rect 5710 -12852 5720 -12792
rect 6096 -12722 6106 -12672
rect 6562 -12662 6622 -12336
rect 6166 -12722 6176 -12672
rect 6096 -12792 6176 -12722
rect 6096 -12852 6106 -12792
rect 6166 -12852 6176 -12792
rect 6552 -12722 6562 -12672
rect 7020 -12662 7080 -12336
rect 6622 -12722 6632 -12672
rect 6552 -12792 6632 -12722
rect 6552 -12852 6562 -12792
rect 6622 -12852 6632 -12792
rect 7010 -12722 7020 -12672
rect 7476 -12662 7536 -12336
rect 7080 -12722 7090 -12672
rect 7010 -12792 7090 -12722
rect 7010 -12852 7020 -12792
rect 7080 -12852 7090 -12792
rect 7466 -12722 7476 -12672
rect 7932 -12662 7992 -12336
rect 7536 -12722 7546 -12672
rect 7466 -12792 7546 -12722
rect 7466 -12852 7476 -12792
rect 7536 -12852 7546 -12792
rect 7922 -12722 7932 -12672
rect 8406 -12662 8466 -12336
rect 7992 -12722 8002 -12672
rect 7922 -12792 8002 -12722
rect 7922 -12852 7932 -12792
rect 7992 -12852 8002 -12792
rect 8396 -12722 8406 -12672
rect 8862 -12662 8922 -12336
rect 8466 -12722 8476 -12672
rect 8396 -12792 8476 -12722
rect 8396 -12852 8406 -12792
rect 8466 -12852 8476 -12792
rect 8852 -12722 8862 -12672
rect 9320 -12662 9380 -12336
rect 8922 -12722 8932 -12672
rect 8852 -12792 8932 -12722
rect 8852 -12852 8862 -12792
rect 8922 -12852 8932 -12792
rect 9310 -12722 9320 -12672
rect 9776 -12662 9836 -12336
rect 9380 -12722 9390 -12672
rect 9310 -12792 9390 -12722
rect 9310 -12852 9320 -12792
rect 9380 -12852 9390 -12792
rect 9766 -12722 9776 -12672
rect 10232 -12662 10292 -12336
rect 9836 -12722 9846 -12672
rect 9766 -12792 9846 -12722
rect 9766 -12852 9776 -12792
rect 9836 -12852 9846 -12792
rect 10222 -12722 10232 -12672
rect 10690 -12662 10750 -12336
rect 10292 -12722 10302 -12672
rect 10222 -12792 10302 -12722
rect 10222 -12852 10232 -12792
rect 10292 -12852 10302 -12792
rect 10680 -12722 10690 -12672
rect 11146 -12662 11206 -12336
rect 10750 -12722 10760 -12672
rect 10680 -12792 10760 -12722
rect 10680 -12852 10690 -12792
rect 10750 -12852 10760 -12792
rect 11136 -12722 11146 -12672
rect 11602 -12662 11662 -12336
rect 11206 -12722 11216 -12672
rect 11136 -12792 11216 -12722
rect 11136 -12852 11146 -12792
rect 11206 -12852 11216 -12792
rect 11592 -12722 11602 -12672
rect 12060 -12662 12120 -12336
rect 11662 -12722 11672 -12672
rect 11592 -12792 11672 -12722
rect 11592 -12852 11602 -12792
rect 11662 -12852 11672 -12792
rect 12050 -12722 12060 -12672
rect 12516 -12662 12576 -12336
rect 12120 -12722 12130 -12672
rect 12050 -12792 12130 -12722
rect 12050 -12852 12060 -12792
rect 12120 -12852 12130 -12792
rect 12506 -12722 12516 -12672
rect 12972 -12662 13032 -12336
rect 12576 -12722 12586 -12672
rect 12506 -12792 12586 -12722
rect 12506 -12852 12516 -12792
rect 12576 -12852 12586 -12792
rect 12962 -12722 12972 -12672
rect 13430 -12662 13490 -12336
rect 13032 -12722 13042 -12672
rect 12962 -12792 13042 -12722
rect 12962 -12852 12972 -12792
rect 13032 -12852 13042 -12792
rect 13420 -12722 13430 -12672
rect 13886 -12662 13946 -12336
rect 13490 -12722 13500 -12672
rect 13420 -12792 13500 -12722
rect 13420 -12852 13430 -12792
rect 13490 -12852 13500 -12792
rect 13876 -12722 13886 -12672
rect 14342 -12662 14402 -12336
rect 13946 -12722 13956 -12672
rect 13876 -12792 13956 -12722
rect 13876 -12852 13886 -12792
rect 13946 -12852 13956 -12792
rect 14332 -12722 14342 -12672
rect 14800 -12662 14860 -12336
rect 14402 -12722 14412 -12672
rect 14332 -12792 14412 -12722
rect 14332 -12852 14342 -12792
rect 14402 -12852 14412 -12792
rect 14790 -12722 14800 -12672
rect 15256 -12662 15316 -12336
rect 14860 -12722 14870 -12672
rect 14790 -12792 14870 -12722
rect 14790 -12852 14800 -12792
rect 14860 -12852 14870 -12792
rect 15246 -12722 15256 -12672
rect 15316 -12722 15326 -12672
rect 15246 -12792 15326 -12722
rect 15246 -12852 15256 -12792
rect 15316 -12852 15326 -12792
rect 170 -13164 230 -12852
rect 160 -13224 170 -13174
rect 626 -13164 686 -12852
rect 230 -13224 240 -13174
rect 160 -13294 240 -13224
rect 160 -13354 170 -13294
rect 230 -13354 240 -13294
rect 616 -13224 626 -13174
rect 1082 -13164 1142 -12852
rect 686 -13224 696 -13174
rect 616 -13294 696 -13224
rect 616 -13354 626 -13294
rect 686 -13354 696 -13294
rect 1072 -13224 1082 -13174
rect 1540 -13164 1600 -12852
rect 1142 -13224 1152 -13174
rect 1072 -13294 1152 -13224
rect 1072 -13354 1082 -13294
rect 1142 -13354 1152 -13294
rect 1530 -13224 1540 -13174
rect 1996 -13164 2056 -12852
rect 1600 -13224 1610 -13174
rect 1530 -13294 1610 -13224
rect 1530 -13354 1540 -13294
rect 1600 -13354 1610 -13294
rect 1986 -13224 1996 -13174
rect 2452 -13164 2512 -12852
rect 2056 -13224 2066 -13174
rect 1986 -13294 2066 -13224
rect 1986 -13354 1996 -13294
rect 2056 -13354 2066 -13294
rect 2442 -13224 2452 -13174
rect 2910 -13164 2970 -12852
rect 2512 -13224 2522 -13174
rect 2442 -13294 2522 -13224
rect 2442 -13354 2452 -13294
rect 2512 -13354 2522 -13294
rect 2900 -13224 2910 -13174
rect 3366 -13164 3426 -12852
rect 2970 -13224 2980 -13174
rect 2900 -13294 2980 -13224
rect 2900 -13354 2910 -13294
rect 2970 -13354 2980 -13294
rect 3356 -13224 3366 -13174
rect 3822 -13164 3882 -12852
rect 3426 -13224 3436 -13174
rect 3356 -13294 3436 -13224
rect 3356 -13354 3366 -13294
rect 3426 -13354 3436 -13294
rect 3812 -13224 3822 -13174
rect 4280 -13164 4340 -12852
rect 3882 -13224 3892 -13174
rect 3812 -13294 3892 -13224
rect 3812 -13354 3822 -13294
rect 3882 -13354 3892 -13294
rect 4270 -13224 4280 -13174
rect 4736 -13164 4796 -12852
rect 4340 -13224 4350 -13174
rect 4270 -13294 4350 -13224
rect 4270 -13354 4280 -13294
rect 4340 -13354 4350 -13294
rect 4726 -13224 4736 -13174
rect 5192 -13164 5252 -12852
rect 4796 -13224 4806 -13174
rect 4726 -13294 4806 -13224
rect 4726 -13354 4736 -13294
rect 4796 -13354 4806 -13294
rect 5182 -13224 5192 -13174
rect 5650 -13164 5710 -12852
rect 5252 -13224 5262 -13174
rect 5182 -13294 5262 -13224
rect 5182 -13354 5192 -13294
rect 5252 -13354 5262 -13294
rect 5640 -13224 5650 -13174
rect 6106 -13164 6166 -12852
rect 5710 -13224 5720 -13174
rect 5640 -13294 5720 -13224
rect 5640 -13354 5650 -13294
rect 5710 -13354 5720 -13294
rect 6096 -13224 6106 -13174
rect 6562 -13164 6622 -12852
rect 6166 -13224 6176 -13174
rect 6096 -13294 6176 -13224
rect 6096 -13354 6106 -13294
rect 6166 -13354 6176 -13294
rect 6552 -13224 6562 -13174
rect 7020 -13164 7080 -12852
rect 6622 -13224 6632 -13174
rect 6552 -13294 6632 -13224
rect 6552 -13354 6562 -13294
rect 6622 -13354 6632 -13294
rect 7010 -13224 7020 -13174
rect 7476 -13164 7536 -12852
rect 7080 -13224 7090 -13174
rect 7010 -13294 7090 -13224
rect 7010 -13354 7020 -13294
rect 7080 -13354 7090 -13294
rect 7466 -13224 7476 -13174
rect 7932 -13164 7992 -12852
rect 7536 -13224 7546 -13174
rect 7466 -13294 7546 -13224
rect 7466 -13354 7476 -13294
rect 7536 -13354 7546 -13294
rect 7922 -13224 7932 -13174
rect 8406 -13164 8466 -12852
rect 7992 -13224 8002 -13174
rect 7922 -13294 8002 -13224
rect 7922 -13354 7932 -13294
rect 7992 -13354 8002 -13294
rect 8396 -13224 8406 -13174
rect 8862 -13164 8922 -12852
rect 8466 -13224 8476 -13174
rect 8396 -13294 8476 -13224
rect 8396 -13354 8406 -13294
rect 8466 -13354 8476 -13294
rect 8852 -13224 8862 -13174
rect 9320 -13164 9380 -12852
rect 8922 -13224 8932 -13174
rect 8852 -13294 8932 -13224
rect 8852 -13354 8862 -13294
rect 8922 -13354 8932 -13294
rect 9310 -13224 9320 -13174
rect 9776 -13164 9836 -12852
rect 9380 -13224 9390 -13174
rect 9310 -13294 9390 -13224
rect 9310 -13354 9320 -13294
rect 9380 -13354 9390 -13294
rect 9766 -13224 9776 -13174
rect 10232 -13164 10292 -12852
rect 9836 -13224 9846 -13174
rect 9766 -13294 9846 -13224
rect 9766 -13354 9776 -13294
rect 9836 -13354 9846 -13294
rect 10222 -13224 10232 -13174
rect 10690 -13164 10750 -12852
rect 10292 -13224 10302 -13174
rect 10222 -13294 10302 -13224
rect 10222 -13354 10232 -13294
rect 10292 -13354 10302 -13294
rect 10680 -13224 10690 -13174
rect 11146 -13164 11206 -12852
rect 10750 -13224 10760 -13174
rect 10680 -13294 10760 -13224
rect 10680 -13354 10690 -13294
rect 10750 -13354 10760 -13294
rect 11136 -13224 11146 -13174
rect 11602 -13164 11662 -12852
rect 11206 -13224 11216 -13174
rect 11136 -13294 11216 -13224
rect 11136 -13354 11146 -13294
rect 11206 -13354 11216 -13294
rect 11592 -13224 11602 -13174
rect 12060 -13164 12120 -12852
rect 11662 -13224 11672 -13174
rect 11592 -13294 11672 -13224
rect 11592 -13354 11602 -13294
rect 11662 -13354 11672 -13294
rect 12050 -13224 12060 -13174
rect 12516 -13164 12576 -12852
rect 12120 -13224 12130 -13174
rect 12050 -13294 12130 -13224
rect 12050 -13354 12060 -13294
rect 12120 -13354 12130 -13294
rect 12506 -13224 12516 -13174
rect 12972 -13164 13032 -12852
rect 12576 -13224 12586 -13174
rect 12506 -13294 12586 -13224
rect 12506 -13354 12516 -13294
rect 12576 -13354 12586 -13294
rect 12962 -13224 12972 -13174
rect 13430 -13164 13490 -12852
rect 13032 -13224 13042 -13174
rect 12962 -13294 13042 -13224
rect 12962 -13354 12972 -13294
rect 13032 -13354 13042 -13294
rect 13420 -13224 13430 -13174
rect 13886 -13164 13946 -12852
rect 13490 -13224 13500 -13174
rect 13420 -13294 13500 -13224
rect 13420 -13354 13430 -13294
rect 13490 -13354 13500 -13294
rect 13876 -13224 13886 -13174
rect 14342 -13164 14402 -12852
rect 13946 -13224 13956 -13174
rect 13876 -13294 13956 -13224
rect 13876 -13354 13886 -13294
rect 13946 -13354 13956 -13294
rect 14332 -13224 14342 -13174
rect 14800 -13164 14860 -12852
rect 14402 -13224 14412 -13174
rect 14332 -13294 14412 -13224
rect 14332 -13354 14342 -13294
rect 14402 -13354 14412 -13294
rect 14790 -13224 14800 -13174
rect 15256 -13164 15316 -12852
rect 14860 -13224 14870 -13174
rect 14790 -13294 14870 -13224
rect 14790 -13354 14800 -13294
rect 14860 -13354 14870 -13294
rect 15246 -13224 15256 -13174
rect 15316 -13224 15326 -13174
rect 15246 -13294 15326 -13224
rect 15246 -13354 15256 -13294
rect 15316 -13354 15326 -13294
rect 170 -13656 230 -13354
rect 160 -13716 170 -13666
rect 626 -13656 686 -13354
rect 230 -13716 240 -13666
rect 160 -13786 240 -13716
rect 160 -13846 170 -13786
rect 230 -13846 240 -13786
rect 616 -13716 626 -13666
rect 1082 -13656 1142 -13354
rect 686 -13716 696 -13666
rect 616 -13786 696 -13716
rect 616 -13846 626 -13786
rect 686 -13846 696 -13786
rect 1072 -13716 1082 -13666
rect 1540 -13656 1600 -13354
rect 1142 -13716 1152 -13666
rect 1072 -13786 1152 -13716
rect 1072 -13846 1082 -13786
rect 1142 -13846 1152 -13786
rect 1530 -13716 1540 -13666
rect 1996 -13656 2056 -13354
rect 1600 -13716 1610 -13666
rect 1530 -13786 1610 -13716
rect 1530 -13846 1540 -13786
rect 1600 -13846 1610 -13786
rect 1986 -13716 1996 -13666
rect 2452 -13656 2512 -13354
rect 2056 -13716 2066 -13666
rect 1986 -13786 2066 -13716
rect 1986 -13846 1996 -13786
rect 2056 -13846 2066 -13786
rect 2442 -13716 2452 -13666
rect 2910 -13656 2970 -13354
rect 2512 -13716 2522 -13666
rect 2442 -13786 2522 -13716
rect 2442 -13846 2452 -13786
rect 2512 -13846 2522 -13786
rect 2900 -13716 2910 -13666
rect 3366 -13656 3426 -13354
rect 2970 -13716 2980 -13666
rect 2900 -13786 2980 -13716
rect 2900 -13846 2910 -13786
rect 2970 -13846 2980 -13786
rect 3356 -13716 3366 -13666
rect 3822 -13656 3882 -13354
rect 3426 -13716 3436 -13666
rect 3356 -13786 3436 -13716
rect 3356 -13846 3366 -13786
rect 3426 -13846 3436 -13786
rect 3812 -13716 3822 -13666
rect 4280 -13656 4340 -13354
rect 3882 -13716 3892 -13666
rect 3812 -13786 3892 -13716
rect 3812 -13846 3822 -13786
rect 3882 -13846 3892 -13786
rect 4270 -13716 4280 -13666
rect 4736 -13656 4796 -13354
rect 4340 -13716 4350 -13666
rect 4270 -13786 4350 -13716
rect 4270 -13846 4280 -13786
rect 4340 -13846 4350 -13786
rect 4726 -13716 4736 -13666
rect 5192 -13656 5252 -13354
rect 4796 -13716 4806 -13666
rect 4726 -13786 4806 -13716
rect 4726 -13846 4736 -13786
rect 4796 -13846 4806 -13786
rect 5182 -13716 5192 -13666
rect 5650 -13656 5710 -13354
rect 5252 -13716 5262 -13666
rect 5182 -13786 5262 -13716
rect 5182 -13846 5192 -13786
rect 5252 -13846 5262 -13786
rect 5640 -13716 5650 -13666
rect 6106 -13656 6166 -13354
rect 5710 -13716 5720 -13666
rect 5640 -13786 5720 -13716
rect 5640 -13846 5650 -13786
rect 5710 -13846 5720 -13786
rect 6096 -13716 6106 -13666
rect 6562 -13656 6622 -13354
rect 6166 -13716 6176 -13666
rect 6096 -13786 6176 -13716
rect 6096 -13846 6106 -13786
rect 6166 -13846 6176 -13786
rect 6552 -13716 6562 -13666
rect 7020 -13656 7080 -13354
rect 6622 -13716 6632 -13666
rect 6552 -13786 6632 -13716
rect 6552 -13846 6562 -13786
rect 6622 -13846 6632 -13786
rect 7010 -13716 7020 -13666
rect 7476 -13656 7536 -13354
rect 7080 -13716 7090 -13666
rect 7010 -13786 7090 -13716
rect 7010 -13846 7020 -13786
rect 7080 -13846 7090 -13786
rect 7466 -13716 7476 -13666
rect 7932 -13656 7992 -13354
rect 7536 -13716 7546 -13666
rect 7466 -13786 7546 -13716
rect 7466 -13846 7476 -13786
rect 7536 -13846 7546 -13786
rect 7922 -13716 7932 -13666
rect 8406 -13656 8466 -13354
rect 7992 -13716 8002 -13666
rect 7922 -13786 8002 -13716
rect 7922 -13846 7932 -13786
rect 7992 -13846 8002 -13786
rect 8396 -13716 8406 -13666
rect 8862 -13656 8922 -13354
rect 8466 -13716 8476 -13666
rect 8396 -13786 8476 -13716
rect 8396 -13846 8406 -13786
rect 8466 -13846 8476 -13786
rect 8852 -13716 8862 -13666
rect 9320 -13656 9380 -13354
rect 8922 -13716 8932 -13666
rect 8852 -13786 8932 -13716
rect 8852 -13846 8862 -13786
rect 8922 -13846 8932 -13786
rect 9310 -13716 9320 -13666
rect 9776 -13656 9836 -13354
rect 9380 -13716 9390 -13666
rect 9310 -13786 9390 -13716
rect 9310 -13846 9320 -13786
rect 9380 -13846 9390 -13786
rect 9766 -13716 9776 -13666
rect 10232 -13656 10292 -13354
rect 9836 -13716 9846 -13666
rect 9766 -13786 9846 -13716
rect 9766 -13846 9776 -13786
rect 9836 -13846 9846 -13786
rect 10222 -13716 10232 -13666
rect 10690 -13656 10750 -13354
rect 10292 -13716 10302 -13666
rect 10222 -13786 10302 -13716
rect 10222 -13846 10232 -13786
rect 10292 -13846 10302 -13786
rect 10680 -13716 10690 -13666
rect 11146 -13656 11206 -13354
rect 10750 -13716 10760 -13666
rect 10680 -13786 10760 -13716
rect 10680 -13846 10690 -13786
rect 10750 -13846 10760 -13786
rect 11136 -13716 11146 -13666
rect 11602 -13656 11662 -13354
rect 11206 -13716 11216 -13666
rect 11136 -13786 11216 -13716
rect 11136 -13846 11146 -13786
rect 11206 -13846 11216 -13786
rect 11592 -13716 11602 -13666
rect 12060 -13656 12120 -13354
rect 11662 -13716 11672 -13666
rect 11592 -13786 11672 -13716
rect 11592 -13846 11602 -13786
rect 11662 -13846 11672 -13786
rect 12050 -13716 12060 -13666
rect 12516 -13656 12576 -13354
rect 12120 -13716 12130 -13666
rect 12050 -13786 12130 -13716
rect 12050 -13846 12060 -13786
rect 12120 -13846 12130 -13786
rect 12506 -13716 12516 -13666
rect 12972 -13656 13032 -13354
rect 12576 -13716 12586 -13666
rect 12506 -13786 12586 -13716
rect 12506 -13846 12516 -13786
rect 12576 -13846 12586 -13786
rect 12962 -13716 12972 -13666
rect 13430 -13656 13490 -13354
rect 13032 -13716 13042 -13666
rect 12962 -13786 13042 -13716
rect 12962 -13846 12972 -13786
rect 13032 -13846 13042 -13786
rect 13420 -13716 13430 -13666
rect 13886 -13656 13946 -13354
rect 13490 -13716 13500 -13666
rect 13420 -13786 13500 -13716
rect 13420 -13846 13430 -13786
rect 13490 -13846 13500 -13786
rect 13876 -13716 13886 -13666
rect 14342 -13656 14402 -13354
rect 13946 -13716 13956 -13666
rect 13876 -13786 13956 -13716
rect 13876 -13846 13886 -13786
rect 13946 -13846 13956 -13786
rect 14332 -13716 14342 -13666
rect 14800 -13656 14860 -13354
rect 14402 -13716 14412 -13666
rect 14332 -13786 14412 -13716
rect 14332 -13846 14342 -13786
rect 14402 -13846 14412 -13786
rect 14790 -13716 14800 -13666
rect 15256 -13656 15316 -13354
rect 14860 -13716 14870 -13666
rect 14790 -13786 14870 -13716
rect 14790 -13846 14800 -13786
rect 14860 -13846 14870 -13786
rect 15246 -13716 15256 -13666
rect 15316 -13716 15326 -13666
rect 15246 -13786 15326 -13716
rect 15246 -13846 15256 -13786
rect 15316 -13846 15326 -13786
rect 170 -14150 230 -13846
rect 160 -14210 170 -14160
rect 626 -14150 686 -13846
rect 230 -14210 240 -14160
rect 160 -14280 240 -14210
rect 160 -14340 170 -14280
rect 230 -14340 240 -14280
rect 616 -14210 626 -14160
rect 1082 -14150 1142 -13846
rect 686 -14210 696 -14160
rect 616 -14280 696 -14210
rect 616 -14340 626 -14280
rect 686 -14340 696 -14280
rect 1072 -14210 1082 -14160
rect 1540 -14150 1600 -13846
rect 1142 -14210 1152 -14160
rect 1072 -14280 1152 -14210
rect 1072 -14340 1082 -14280
rect 1142 -14340 1152 -14280
rect 1530 -14210 1540 -14160
rect 1996 -14150 2056 -13846
rect 1600 -14210 1610 -14160
rect 1530 -14280 1610 -14210
rect 1530 -14340 1540 -14280
rect 1600 -14340 1610 -14280
rect 1986 -14210 1996 -14160
rect 2452 -14150 2512 -13846
rect 2056 -14210 2066 -14160
rect 1986 -14280 2066 -14210
rect 1986 -14340 1996 -14280
rect 2056 -14340 2066 -14280
rect 2442 -14210 2452 -14160
rect 2910 -14150 2970 -13846
rect 2512 -14210 2522 -14160
rect 2442 -14280 2522 -14210
rect 2442 -14340 2452 -14280
rect 2512 -14340 2522 -14280
rect 2900 -14210 2910 -14160
rect 3366 -14150 3426 -13846
rect 2970 -14210 2980 -14160
rect 2900 -14280 2980 -14210
rect 2900 -14340 2910 -14280
rect 2970 -14340 2980 -14280
rect 3356 -14210 3366 -14160
rect 3822 -14150 3882 -13846
rect 3426 -14210 3436 -14160
rect 3356 -14280 3436 -14210
rect 3356 -14340 3366 -14280
rect 3426 -14340 3436 -14280
rect 3812 -14210 3822 -14160
rect 4280 -14150 4340 -13846
rect 3882 -14210 3892 -14160
rect 3812 -14280 3892 -14210
rect 3812 -14340 3822 -14280
rect 3882 -14340 3892 -14280
rect 4270 -14210 4280 -14160
rect 4736 -14150 4796 -13846
rect 4340 -14210 4350 -14160
rect 4270 -14280 4350 -14210
rect 4270 -14340 4280 -14280
rect 4340 -14340 4350 -14280
rect 4726 -14210 4736 -14160
rect 5192 -14150 5252 -13846
rect 4796 -14210 4806 -14160
rect 4726 -14280 4806 -14210
rect 4726 -14340 4736 -14280
rect 4796 -14340 4806 -14280
rect 5182 -14210 5192 -14160
rect 5650 -14150 5710 -13846
rect 5252 -14210 5262 -14160
rect 5182 -14280 5262 -14210
rect 5182 -14340 5192 -14280
rect 5252 -14340 5262 -14280
rect 5640 -14210 5650 -14160
rect 6106 -14150 6166 -13846
rect 5710 -14210 5720 -14160
rect 5640 -14280 5720 -14210
rect 5640 -14340 5650 -14280
rect 5710 -14340 5720 -14280
rect 6096 -14210 6106 -14160
rect 6562 -14150 6622 -13846
rect 6166 -14210 6176 -14160
rect 6096 -14280 6176 -14210
rect 6096 -14340 6106 -14280
rect 6166 -14340 6176 -14280
rect 6552 -14210 6562 -14160
rect 7020 -14150 7080 -13846
rect 6622 -14210 6632 -14160
rect 6552 -14280 6632 -14210
rect 6552 -14340 6562 -14280
rect 6622 -14340 6632 -14280
rect 7010 -14210 7020 -14160
rect 7476 -14150 7536 -13846
rect 7080 -14210 7090 -14160
rect 7010 -14280 7090 -14210
rect 7010 -14340 7020 -14280
rect 7080 -14340 7090 -14280
rect 7466 -14210 7476 -14160
rect 7932 -14150 7992 -13846
rect 7536 -14210 7546 -14160
rect 7466 -14280 7546 -14210
rect 7466 -14340 7476 -14280
rect 7536 -14340 7546 -14280
rect 7922 -14210 7932 -14160
rect 8406 -14150 8466 -13846
rect 7992 -14210 8002 -14160
rect 7922 -14280 8002 -14210
rect 7922 -14340 7932 -14280
rect 7992 -14340 8002 -14280
rect 8396 -14210 8406 -14160
rect 8862 -14150 8922 -13846
rect 8466 -14210 8476 -14160
rect 8396 -14280 8476 -14210
rect 8396 -14340 8406 -14280
rect 8466 -14340 8476 -14280
rect 8852 -14210 8862 -14160
rect 9320 -14150 9380 -13846
rect 8922 -14210 8932 -14160
rect 8852 -14280 8932 -14210
rect 8852 -14340 8862 -14280
rect 8922 -14340 8932 -14280
rect 9310 -14210 9320 -14160
rect 9776 -14150 9836 -13846
rect 9380 -14210 9390 -14160
rect 9310 -14280 9390 -14210
rect 9310 -14340 9320 -14280
rect 9380 -14340 9390 -14280
rect 9766 -14210 9776 -14160
rect 10232 -14150 10292 -13846
rect 9836 -14210 9846 -14160
rect 9766 -14280 9846 -14210
rect 9766 -14340 9776 -14280
rect 9836 -14340 9846 -14280
rect 10222 -14210 10232 -14160
rect 10690 -14150 10750 -13846
rect 10292 -14210 10302 -14160
rect 10222 -14280 10302 -14210
rect 10222 -14340 10232 -14280
rect 10292 -14340 10302 -14280
rect 10680 -14210 10690 -14160
rect 11146 -14150 11206 -13846
rect 10750 -14210 10760 -14160
rect 10680 -14280 10760 -14210
rect 10680 -14340 10690 -14280
rect 10750 -14340 10760 -14280
rect 11136 -14210 11146 -14160
rect 11602 -14150 11662 -13846
rect 11206 -14210 11216 -14160
rect 11136 -14280 11216 -14210
rect 11136 -14340 11146 -14280
rect 11206 -14340 11216 -14280
rect 11592 -14210 11602 -14160
rect 12060 -14150 12120 -13846
rect 11662 -14210 11672 -14160
rect 11592 -14280 11672 -14210
rect 11592 -14340 11602 -14280
rect 11662 -14340 11672 -14280
rect 12050 -14210 12060 -14160
rect 12516 -14150 12576 -13846
rect 12120 -14210 12130 -14160
rect 12050 -14280 12130 -14210
rect 12050 -14340 12060 -14280
rect 12120 -14340 12130 -14280
rect 12506 -14210 12516 -14160
rect 12972 -14150 13032 -13846
rect 12576 -14210 12586 -14160
rect 12506 -14280 12586 -14210
rect 12506 -14340 12516 -14280
rect 12576 -14340 12586 -14280
rect 12962 -14210 12972 -14160
rect 13430 -14150 13490 -13846
rect 13032 -14210 13042 -14160
rect 12962 -14280 13042 -14210
rect 12962 -14340 12972 -14280
rect 13032 -14340 13042 -14280
rect 13420 -14210 13430 -14160
rect 13886 -14150 13946 -13846
rect 13490 -14210 13500 -14160
rect 13420 -14280 13500 -14210
rect 13420 -14340 13430 -14280
rect 13490 -14340 13500 -14280
rect 13876 -14210 13886 -14160
rect 14342 -14150 14402 -13846
rect 13946 -14210 13956 -14160
rect 13876 -14280 13956 -14210
rect 13876 -14340 13886 -14280
rect 13946 -14340 13956 -14280
rect 14332 -14210 14342 -14160
rect 14800 -14150 14860 -13846
rect 14402 -14210 14412 -14160
rect 14332 -14280 14412 -14210
rect 14332 -14340 14342 -14280
rect 14402 -14340 14412 -14280
rect 14790 -14210 14800 -14160
rect 15256 -14150 15316 -13846
rect 14860 -14210 14870 -14160
rect 14790 -14280 14870 -14210
rect 14790 -14340 14800 -14280
rect 14860 -14340 14870 -14280
rect 15246 -14210 15256 -14160
rect 15316 -14210 15326 -14160
rect 15246 -14280 15326 -14210
rect 15246 -14340 15256 -14280
rect 15316 -14340 15326 -14280
rect 170 -14652 230 -14340
rect 160 -14712 170 -14662
rect 626 -14652 686 -14340
rect 230 -14712 240 -14662
rect 160 -14782 240 -14712
rect 160 -14842 170 -14782
rect 230 -14842 240 -14782
rect 616 -14712 626 -14662
rect 1082 -14652 1142 -14340
rect 686 -14712 696 -14662
rect 616 -14782 696 -14712
rect 616 -14842 626 -14782
rect 686 -14842 696 -14782
rect 1072 -14712 1082 -14662
rect 1540 -14652 1600 -14340
rect 1142 -14712 1152 -14662
rect 1072 -14782 1152 -14712
rect 1072 -14842 1082 -14782
rect 1142 -14842 1152 -14782
rect 1530 -14712 1540 -14662
rect 1996 -14652 2056 -14340
rect 1600 -14712 1610 -14662
rect 1530 -14782 1610 -14712
rect 1530 -14842 1540 -14782
rect 1600 -14842 1610 -14782
rect 1986 -14712 1996 -14662
rect 2452 -14652 2512 -14340
rect 2056 -14712 2066 -14662
rect 1986 -14782 2066 -14712
rect 1986 -14842 1996 -14782
rect 2056 -14842 2066 -14782
rect 2442 -14712 2452 -14662
rect 2910 -14652 2970 -14340
rect 2512 -14712 2522 -14662
rect 2442 -14782 2522 -14712
rect 2442 -14842 2452 -14782
rect 2512 -14842 2522 -14782
rect 2900 -14712 2910 -14662
rect 3366 -14652 3426 -14340
rect 2970 -14712 2980 -14662
rect 2900 -14782 2980 -14712
rect 2900 -14842 2910 -14782
rect 2970 -14842 2980 -14782
rect 3356 -14712 3366 -14662
rect 3822 -14652 3882 -14340
rect 3426 -14712 3436 -14662
rect 3356 -14782 3436 -14712
rect 3356 -14842 3366 -14782
rect 3426 -14842 3436 -14782
rect 3812 -14712 3822 -14662
rect 4280 -14652 4340 -14340
rect 3882 -14712 3892 -14662
rect 3812 -14782 3892 -14712
rect 3812 -14842 3822 -14782
rect 3882 -14842 3892 -14782
rect 4270 -14712 4280 -14662
rect 4736 -14652 4796 -14340
rect 4340 -14712 4350 -14662
rect 4270 -14782 4350 -14712
rect 4270 -14842 4280 -14782
rect 4340 -14842 4350 -14782
rect 4726 -14712 4736 -14662
rect 5192 -14652 5252 -14340
rect 4796 -14712 4806 -14662
rect 4726 -14782 4806 -14712
rect 4726 -14842 4736 -14782
rect 4796 -14842 4806 -14782
rect 5182 -14712 5192 -14662
rect 5650 -14652 5710 -14340
rect 5252 -14712 5262 -14662
rect 5182 -14782 5262 -14712
rect 5182 -14842 5192 -14782
rect 5252 -14842 5262 -14782
rect 5640 -14712 5650 -14662
rect 6106 -14652 6166 -14340
rect 5710 -14712 5720 -14662
rect 5640 -14782 5720 -14712
rect 5640 -14842 5650 -14782
rect 5710 -14842 5720 -14782
rect 6096 -14712 6106 -14662
rect 6562 -14652 6622 -14340
rect 6166 -14712 6176 -14662
rect 6096 -14782 6176 -14712
rect 6096 -14842 6106 -14782
rect 6166 -14842 6176 -14782
rect 6552 -14712 6562 -14662
rect 7020 -14652 7080 -14340
rect 6622 -14712 6632 -14662
rect 6552 -14782 6632 -14712
rect 6552 -14842 6562 -14782
rect 6622 -14842 6632 -14782
rect 7010 -14712 7020 -14662
rect 7476 -14652 7536 -14340
rect 7080 -14712 7090 -14662
rect 7010 -14782 7090 -14712
rect 7010 -14842 7020 -14782
rect 7080 -14842 7090 -14782
rect 7466 -14712 7476 -14662
rect 7932 -14652 7992 -14340
rect 7536 -14712 7546 -14662
rect 7466 -14782 7546 -14712
rect 7466 -14842 7476 -14782
rect 7536 -14842 7546 -14782
rect 7922 -14712 7932 -14662
rect 8406 -14652 8466 -14340
rect 7992 -14712 8002 -14662
rect 7922 -14782 8002 -14712
rect 7922 -14842 7932 -14782
rect 7992 -14842 8002 -14782
rect 8396 -14712 8406 -14662
rect 8862 -14652 8922 -14340
rect 8466 -14712 8476 -14662
rect 8396 -14782 8476 -14712
rect 8396 -14842 8406 -14782
rect 8466 -14842 8476 -14782
rect 8852 -14712 8862 -14662
rect 9320 -14652 9380 -14340
rect 8922 -14712 8932 -14662
rect 8852 -14782 8932 -14712
rect 8852 -14842 8862 -14782
rect 8922 -14842 8932 -14782
rect 9310 -14712 9320 -14662
rect 9776 -14652 9836 -14340
rect 9380 -14712 9390 -14662
rect 9310 -14782 9390 -14712
rect 9310 -14842 9320 -14782
rect 9380 -14842 9390 -14782
rect 9766 -14712 9776 -14662
rect 10232 -14652 10292 -14340
rect 9836 -14712 9846 -14662
rect 9766 -14782 9846 -14712
rect 9766 -14842 9776 -14782
rect 9836 -14842 9846 -14782
rect 10222 -14712 10232 -14662
rect 10690 -14652 10750 -14340
rect 10292 -14712 10302 -14662
rect 10222 -14782 10302 -14712
rect 10222 -14842 10232 -14782
rect 10292 -14842 10302 -14782
rect 10680 -14712 10690 -14662
rect 11146 -14652 11206 -14340
rect 10750 -14712 10760 -14662
rect 10680 -14782 10760 -14712
rect 10680 -14842 10690 -14782
rect 10750 -14842 10760 -14782
rect 11136 -14712 11146 -14662
rect 11602 -14652 11662 -14340
rect 11206 -14712 11216 -14662
rect 11136 -14782 11216 -14712
rect 11136 -14842 11146 -14782
rect 11206 -14842 11216 -14782
rect 11592 -14712 11602 -14662
rect 12060 -14652 12120 -14340
rect 11662 -14712 11672 -14662
rect 11592 -14782 11672 -14712
rect 11592 -14842 11602 -14782
rect 11662 -14842 11672 -14782
rect 12050 -14712 12060 -14662
rect 12516 -14652 12576 -14340
rect 12120 -14712 12130 -14662
rect 12050 -14782 12130 -14712
rect 12050 -14842 12060 -14782
rect 12120 -14842 12130 -14782
rect 12506 -14712 12516 -14662
rect 12972 -14652 13032 -14340
rect 12576 -14712 12586 -14662
rect 12506 -14782 12586 -14712
rect 12506 -14842 12516 -14782
rect 12576 -14842 12586 -14782
rect 12962 -14712 12972 -14662
rect 13430 -14652 13490 -14340
rect 13032 -14712 13042 -14662
rect 12962 -14782 13042 -14712
rect 12962 -14842 12972 -14782
rect 13032 -14842 13042 -14782
rect 13420 -14712 13430 -14662
rect 13886 -14652 13946 -14340
rect 13490 -14712 13500 -14662
rect 13420 -14782 13500 -14712
rect 13420 -14842 13430 -14782
rect 13490 -14842 13500 -14782
rect 13876 -14712 13886 -14662
rect 14342 -14652 14402 -14340
rect 13946 -14712 13956 -14662
rect 13876 -14782 13956 -14712
rect 13876 -14842 13886 -14782
rect 13946 -14842 13956 -14782
rect 14332 -14712 14342 -14662
rect 14800 -14652 14860 -14340
rect 14402 -14712 14412 -14662
rect 14332 -14782 14412 -14712
rect 14332 -14842 14342 -14782
rect 14402 -14842 14412 -14782
rect 14790 -14712 14800 -14662
rect 15256 -14652 15316 -14340
rect 14860 -14712 14870 -14662
rect 14790 -14782 14870 -14712
rect 14790 -14842 14800 -14782
rect 14860 -14842 14870 -14782
rect 15246 -14712 15256 -14662
rect 15316 -14712 15326 -14662
rect 15246 -14782 15326 -14712
rect 15246 -14842 15256 -14782
rect 15316 -14842 15326 -14782
rect 170 -15144 230 -14842
rect 160 -15204 170 -15154
rect 626 -15144 686 -14842
rect 230 -15204 240 -15154
rect 160 -15274 240 -15204
rect 160 -15334 170 -15274
rect 230 -15334 240 -15274
rect 616 -15204 626 -15154
rect 1082 -15144 1142 -14842
rect 686 -15204 696 -15154
rect 616 -15274 696 -15204
rect 616 -15334 626 -15274
rect 686 -15334 696 -15274
rect 1072 -15204 1082 -15154
rect 1540 -15144 1600 -14842
rect 1142 -15204 1152 -15154
rect 1072 -15274 1152 -15204
rect 1072 -15334 1082 -15274
rect 1142 -15334 1152 -15274
rect 1530 -15204 1540 -15154
rect 1996 -15144 2056 -14842
rect 1600 -15204 1610 -15154
rect 1530 -15274 1610 -15204
rect 1530 -15334 1540 -15274
rect 1600 -15334 1610 -15274
rect 1986 -15204 1996 -15154
rect 2452 -15144 2512 -14842
rect 2056 -15204 2066 -15154
rect 1986 -15274 2066 -15204
rect 1986 -15334 1996 -15274
rect 2056 -15334 2066 -15274
rect 2442 -15204 2452 -15154
rect 2910 -15144 2970 -14842
rect 2512 -15204 2522 -15154
rect 2442 -15274 2522 -15204
rect 2442 -15334 2452 -15274
rect 2512 -15334 2522 -15274
rect 2900 -15204 2910 -15154
rect 3366 -15144 3426 -14842
rect 2970 -15204 2980 -15154
rect 2900 -15274 2980 -15204
rect 2900 -15334 2910 -15274
rect 2970 -15334 2980 -15274
rect 3356 -15204 3366 -15154
rect 3822 -15144 3882 -14842
rect 3426 -15204 3436 -15154
rect 3356 -15274 3436 -15204
rect 3356 -15334 3366 -15274
rect 3426 -15334 3436 -15274
rect 3812 -15204 3822 -15154
rect 4280 -15144 4340 -14842
rect 3882 -15204 3892 -15154
rect 3812 -15274 3892 -15204
rect 3812 -15334 3822 -15274
rect 3882 -15334 3892 -15274
rect 4270 -15204 4280 -15154
rect 4736 -15144 4796 -14842
rect 4340 -15204 4350 -15154
rect 4270 -15274 4350 -15204
rect 4270 -15334 4280 -15274
rect 4340 -15334 4350 -15274
rect 4726 -15204 4736 -15154
rect 5192 -15144 5252 -14842
rect 4796 -15204 4806 -15154
rect 4726 -15274 4806 -15204
rect 4726 -15334 4736 -15274
rect 4796 -15334 4806 -15274
rect 5182 -15204 5192 -15154
rect 5650 -15144 5710 -14842
rect 5252 -15204 5262 -15154
rect 5182 -15274 5262 -15204
rect 5182 -15334 5192 -15274
rect 5252 -15334 5262 -15274
rect 5640 -15204 5650 -15154
rect 6106 -15144 6166 -14842
rect 5710 -15204 5720 -15154
rect 5640 -15274 5720 -15204
rect 5640 -15334 5650 -15274
rect 5710 -15334 5720 -15274
rect 6096 -15204 6106 -15154
rect 6562 -15144 6622 -14842
rect 6166 -15204 6176 -15154
rect 6096 -15274 6176 -15204
rect 6096 -15334 6106 -15274
rect 6166 -15334 6176 -15274
rect 6552 -15204 6562 -15154
rect 7020 -15144 7080 -14842
rect 6622 -15204 6632 -15154
rect 6552 -15274 6632 -15204
rect 6552 -15334 6562 -15274
rect 6622 -15334 6632 -15274
rect 7010 -15204 7020 -15154
rect 7476 -15144 7536 -14842
rect 7080 -15204 7090 -15154
rect 7010 -15274 7090 -15204
rect 7010 -15334 7020 -15274
rect 7080 -15334 7090 -15274
rect 7466 -15204 7476 -15154
rect 7932 -15144 7992 -14842
rect 7536 -15204 7546 -15154
rect 7466 -15274 7546 -15204
rect 7466 -15334 7476 -15274
rect 7536 -15334 7546 -15274
rect 7922 -15204 7932 -15154
rect 8406 -15144 8466 -14842
rect 7992 -15204 8002 -15154
rect 7922 -15274 8002 -15204
rect 7922 -15334 7932 -15274
rect 7992 -15334 8002 -15274
rect 8396 -15204 8406 -15154
rect 8862 -15144 8922 -14842
rect 8466 -15204 8476 -15154
rect 8396 -15274 8476 -15204
rect 8396 -15334 8406 -15274
rect 8466 -15334 8476 -15274
rect 8852 -15204 8862 -15154
rect 9320 -15144 9380 -14842
rect 8922 -15204 8932 -15154
rect 8852 -15274 8932 -15204
rect 8852 -15334 8862 -15274
rect 8922 -15334 8932 -15274
rect 9310 -15204 9320 -15154
rect 9776 -15144 9836 -14842
rect 9380 -15204 9390 -15154
rect 9310 -15274 9390 -15204
rect 9310 -15334 9320 -15274
rect 9380 -15334 9390 -15274
rect 9766 -15204 9776 -15154
rect 10232 -15144 10292 -14842
rect 9836 -15204 9846 -15154
rect 9766 -15274 9846 -15204
rect 9766 -15334 9776 -15274
rect 9836 -15334 9846 -15274
rect 10222 -15204 10232 -15154
rect 10690 -15144 10750 -14842
rect 10292 -15204 10302 -15154
rect 10222 -15274 10302 -15204
rect 10222 -15334 10232 -15274
rect 10292 -15334 10302 -15274
rect 10680 -15204 10690 -15154
rect 11146 -15144 11206 -14842
rect 10750 -15204 10760 -15154
rect 10680 -15274 10760 -15204
rect 10680 -15334 10690 -15274
rect 10750 -15334 10760 -15274
rect 11136 -15204 11146 -15154
rect 11602 -15144 11662 -14842
rect 11206 -15204 11216 -15154
rect 11136 -15274 11216 -15204
rect 11136 -15334 11146 -15274
rect 11206 -15334 11216 -15274
rect 11592 -15204 11602 -15154
rect 12060 -15144 12120 -14842
rect 11662 -15204 11672 -15154
rect 11592 -15274 11672 -15204
rect 11592 -15334 11602 -15274
rect 11662 -15334 11672 -15274
rect 12050 -15204 12060 -15154
rect 12516 -15144 12576 -14842
rect 12120 -15204 12130 -15154
rect 12050 -15274 12130 -15204
rect 12050 -15334 12060 -15274
rect 12120 -15334 12130 -15274
rect 12506 -15204 12516 -15154
rect 12972 -15144 13032 -14842
rect 12576 -15204 12586 -15154
rect 12506 -15274 12586 -15204
rect 12506 -15334 12516 -15274
rect 12576 -15334 12586 -15274
rect 12962 -15204 12972 -15154
rect 13430 -15144 13490 -14842
rect 13032 -15204 13042 -15154
rect 12962 -15274 13042 -15204
rect 12962 -15334 12972 -15274
rect 13032 -15334 13042 -15274
rect 13420 -15204 13430 -15154
rect 13886 -15144 13946 -14842
rect 13490 -15204 13500 -15154
rect 13420 -15274 13500 -15204
rect 13420 -15334 13430 -15274
rect 13490 -15334 13500 -15274
rect 13876 -15204 13886 -15154
rect 14342 -15144 14402 -14842
rect 13946 -15204 13956 -15154
rect 13876 -15274 13956 -15204
rect 13876 -15334 13886 -15274
rect 13946 -15334 13956 -15274
rect 14332 -15204 14342 -15154
rect 14800 -15144 14860 -14842
rect 14402 -15204 14412 -15154
rect 14332 -15274 14412 -15204
rect 14332 -15334 14342 -15274
rect 14402 -15334 14412 -15274
rect 14790 -15204 14800 -15154
rect 15256 -15144 15316 -14842
rect 14860 -15204 14870 -15154
rect 14790 -15274 14870 -15204
rect 14790 -15334 14800 -15274
rect 14860 -15334 14870 -15274
rect 15246 -15204 15256 -15154
rect 15316 -15204 15326 -15154
rect 15246 -15274 15326 -15204
rect 15246 -15334 15256 -15274
rect 15316 -15334 15326 -15274
rect 170 -15660 230 -15334
rect 160 -15720 170 -15670
rect 626 -15660 686 -15334
rect 230 -15720 240 -15670
rect 160 -15790 240 -15720
rect 160 -15850 170 -15790
rect 230 -15850 240 -15790
rect 616 -15720 626 -15670
rect 1082 -15660 1142 -15334
rect 686 -15720 696 -15670
rect 616 -15790 696 -15720
rect 616 -15850 626 -15790
rect 686 -15850 696 -15790
rect 1072 -15720 1082 -15670
rect 1540 -15660 1600 -15334
rect 1142 -15720 1152 -15670
rect 1072 -15790 1152 -15720
rect 1072 -15850 1082 -15790
rect 1142 -15850 1152 -15790
rect 1530 -15720 1540 -15670
rect 1996 -15660 2056 -15334
rect 1600 -15720 1610 -15670
rect 1530 -15790 1610 -15720
rect 1530 -15850 1540 -15790
rect 1600 -15850 1610 -15790
rect 1986 -15720 1996 -15670
rect 2452 -15660 2512 -15334
rect 2056 -15720 2066 -15670
rect 1986 -15790 2066 -15720
rect 1986 -15850 1996 -15790
rect 2056 -15850 2066 -15790
rect 2442 -15720 2452 -15670
rect 2910 -15660 2970 -15334
rect 2512 -15720 2522 -15670
rect 2442 -15790 2522 -15720
rect 2442 -15850 2452 -15790
rect 2512 -15850 2522 -15790
rect 2900 -15720 2910 -15670
rect 3366 -15660 3426 -15334
rect 2970 -15720 2980 -15670
rect 2900 -15790 2980 -15720
rect 2900 -15850 2910 -15790
rect 2970 -15850 2980 -15790
rect 3356 -15720 3366 -15670
rect 3822 -15660 3882 -15334
rect 3426 -15720 3436 -15670
rect 3356 -15790 3436 -15720
rect 3356 -15850 3366 -15790
rect 3426 -15850 3436 -15790
rect 3812 -15720 3822 -15670
rect 4280 -15660 4340 -15334
rect 3882 -15720 3892 -15670
rect 3812 -15790 3892 -15720
rect 3812 -15850 3822 -15790
rect 3882 -15850 3892 -15790
rect 4270 -15720 4280 -15670
rect 4736 -15660 4796 -15334
rect 4340 -15720 4350 -15670
rect 4270 -15790 4350 -15720
rect 4270 -15850 4280 -15790
rect 4340 -15850 4350 -15790
rect 4726 -15720 4736 -15670
rect 5192 -15660 5252 -15334
rect 4796 -15720 4806 -15670
rect 4726 -15790 4806 -15720
rect 4726 -15850 4736 -15790
rect 4796 -15850 4806 -15790
rect 5182 -15720 5192 -15670
rect 5650 -15660 5710 -15334
rect 5252 -15720 5262 -15670
rect 5182 -15790 5262 -15720
rect 5182 -15850 5192 -15790
rect 5252 -15850 5262 -15790
rect 5640 -15720 5650 -15670
rect 6106 -15660 6166 -15334
rect 5710 -15720 5720 -15670
rect 5640 -15790 5720 -15720
rect 5640 -15850 5650 -15790
rect 5710 -15850 5720 -15790
rect 6096 -15720 6106 -15670
rect 6562 -15660 6622 -15334
rect 6166 -15720 6176 -15670
rect 6096 -15790 6176 -15720
rect 6096 -15850 6106 -15790
rect 6166 -15850 6176 -15790
rect 6552 -15720 6562 -15670
rect 7020 -15660 7080 -15334
rect 6622 -15720 6632 -15670
rect 6552 -15790 6632 -15720
rect 6552 -15850 6562 -15790
rect 6622 -15850 6632 -15790
rect 7010 -15720 7020 -15670
rect 7476 -15660 7536 -15334
rect 7080 -15720 7090 -15670
rect 7010 -15790 7090 -15720
rect 7010 -15850 7020 -15790
rect 7080 -15850 7090 -15790
rect 7466 -15720 7476 -15670
rect 7932 -15660 7992 -15334
rect 7536 -15720 7546 -15670
rect 7466 -15790 7546 -15720
rect 7466 -15850 7476 -15790
rect 7536 -15850 7546 -15790
rect 7922 -15720 7932 -15670
rect 8406 -15660 8466 -15334
rect 7992 -15720 8002 -15670
rect 7922 -15790 8002 -15720
rect 7922 -15850 7932 -15790
rect 7992 -15850 8002 -15790
rect 8396 -15720 8406 -15670
rect 8862 -15660 8922 -15334
rect 8466 -15720 8476 -15670
rect 8396 -15790 8476 -15720
rect 8396 -15850 8406 -15790
rect 8466 -15850 8476 -15790
rect 8852 -15720 8862 -15670
rect 9320 -15660 9380 -15334
rect 8922 -15720 8932 -15670
rect 8852 -15790 8932 -15720
rect 8852 -15850 8862 -15790
rect 8922 -15850 8932 -15790
rect 9310 -15720 9320 -15670
rect 9776 -15660 9836 -15334
rect 9380 -15720 9390 -15670
rect 9310 -15790 9390 -15720
rect 9310 -15850 9320 -15790
rect 9380 -15850 9390 -15790
rect 9766 -15720 9776 -15670
rect 10232 -15660 10292 -15334
rect 9836 -15720 9846 -15670
rect 9766 -15790 9846 -15720
rect 9766 -15850 9776 -15790
rect 9836 -15850 9846 -15790
rect 10222 -15720 10232 -15670
rect 10690 -15660 10750 -15334
rect 10292 -15720 10302 -15670
rect 10222 -15790 10302 -15720
rect 10222 -15850 10232 -15790
rect 10292 -15850 10302 -15790
rect 10680 -15720 10690 -15670
rect 11146 -15660 11206 -15334
rect 10750 -15720 10760 -15670
rect 10680 -15790 10760 -15720
rect 10680 -15850 10690 -15790
rect 10750 -15850 10760 -15790
rect 11136 -15720 11146 -15670
rect 11602 -15660 11662 -15334
rect 11206 -15720 11216 -15670
rect 11136 -15790 11216 -15720
rect 11136 -15850 11146 -15790
rect 11206 -15850 11216 -15790
rect 11592 -15720 11602 -15670
rect 12060 -15660 12120 -15334
rect 11662 -15720 11672 -15670
rect 11592 -15790 11672 -15720
rect 11592 -15850 11602 -15790
rect 11662 -15850 11672 -15790
rect 12050 -15720 12060 -15670
rect 12516 -15660 12576 -15334
rect 12120 -15720 12130 -15670
rect 12050 -15790 12130 -15720
rect 12050 -15850 12060 -15790
rect 12120 -15850 12130 -15790
rect 12506 -15720 12516 -15670
rect 12972 -15660 13032 -15334
rect 12576 -15720 12586 -15670
rect 12506 -15790 12586 -15720
rect 12506 -15850 12516 -15790
rect 12576 -15850 12586 -15790
rect 12962 -15720 12972 -15670
rect 13430 -15660 13490 -15334
rect 13032 -15720 13042 -15670
rect 12962 -15790 13042 -15720
rect 12962 -15850 12972 -15790
rect 13032 -15850 13042 -15790
rect 13420 -15720 13430 -15670
rect 13886 -15660 13946 -15334
rect 13490 -15720 13500 -15670
rect 13420 -15790 13500 -15720
rect 13420 -15850 13430 -15790
rect 13490 -15850 13500 -15790
rect 13876 -15720 13886 -15670
rect 14342 -15660 14402 -15334
rect 13946 -15720 13956 -15670
rect 13876 -15790 13956 -15720
rect 13876 -15850 13886 -15790
rect 13946 -15850 13956 -15790
rect 14332 -15720 14342 -15670
rect 14800 -15660 14860 -15334
rect 14402 -15720 14412 -15670
rect 14332 -15790 14412 -15720
rect 14332 -15850 14342 -15790
rect 14402 -15850 14412 -15790
rect 14790 -15720 14800 -15670
rect 15256 -15660 15316 -15334
rect 14860 -15720 14870 -15670
rect 14790 -15790 14870 -15720
rect 14790 -15850 14800 -15790
rect 14860 -15850 14870 -15790
rect 15246 -15720 15256 -15670
rect 15316 -15720 15326 -15670
rect 15246 -15790 15326 -15720
rect 15246 -15850 15256 -15790
rect 15316 -15850 15326 -15790
rect 170 -16162 230 -15850
rect 160 -16222 170 -16172
rect 626 -16162 686 -15850
rect 230 -16222 240 -16172
rect 160 -16292 240 -16222
rect 160 -16352 170 -16292
rect 230 -16352 240 -16292
rect 616 -16222 626 -16172
rect 1082 -16162 1142 -15850
rect 686 -16222 696 -16172
rect 616 -16292 696 -16222
rect 616 -16352 626 -16292
rect 686 -16352 696 -16292
rect 1072 -16222 1082 -16172
rect 1540 -16162 1600 -15850
rect 1142 -16222 1152 -16172
rect 1072 -16292 1152 -16222
rect 1072 -16352 1082 -16292
rect 1142 -16352 1152 -16292
rect 1530 -16222 1540 -16172
rect 1996 -16162 2056 -15850
rect 1600 -16222 1610 -16172
rect 1530 -16292 1610 -16222
rect 1530 -16352 1540 -16292
rect 1600 -16352 1610 -16292
rect 1986 -16222 1996 -16172
rect 2452 -16162 2512 -15850
rect 2056 -16222 2066 -16172
rect 1986 -16292 2066 -16222
rect 1986 -16352 1996 -16292
rect 2056 -16352 2066 -16292
rect 2442 -16222 2452 -16172
rect 2910 -16162 2970 -15850
rect 2512 -16222 2522 -16172
rect 2442 -16292 2522 -16222
rect 2442 -16352 2452 -16292
rect 2512 -16352 2522 -16292
rect 2900 -16222 2910 -16172
rect 3366 -16162 3426 -15850
rect 2970 -16222 2980 -16172
rect 2900 -16292 2980 -16222
rect 2900 -16352 2910 -16292
rect 2970 -16352 2980 -16292
rect 3356 -16222 3366 -16172
rect 3822 -16162 3882 -15850
rect 3426 -16222 3436 -16172
rect 3356 -16292 3436 -16222
rect 3356 -16352 3366 -16292
rect 3426 -16352 3436 -16292
rect 3812 -16222 3822 -16172
rect 4280 -16162 4340 -15850
rect 3882 -16222 3892 -16172
rect 3812 -16292 3892 -16222
rect 3812 -16352 3822 -16292
rect 3882 -16352 3892 -16292
rect 4270 -16222 4280 -16172
rect 4736 -16162 4796 -15850
rect 4340 -16222 4350 -16172
rect 4270 -16292 4350 -16222
rect 4270 -16352 4280 -16292
rect 4340 -16352 4350 -16292
rect 4726 -16222 4736 -16172
rect 5192 -16162 5252 -15850
rect 4796 -16222 4806 -16172
rect 4726 -16292 4806 -16222
rect 4726 -16352 4736 -16292
rect 4796 -16352 4806 -16292
rect 5182 -16222 5192 -16172
rect 5650 -16162 5710 -15850
rect 5252 -16222 5262 -16172
rect 5182 -16292 5262 -16222
rect 5182 -16352 5192 -16292
rect 5252 -16352 5262 -16292
rect 5640 -16222 5650 -16172
rect 6106 -16162 6166 -15850
rect 5710 -16222 5720 -16172
rect 5640 -16292 5720 -16222
rect 5640 -16352 5650 -16292
rect 5710 -16352 5720 -16292
rect 6096 -16222 6106 -16172
rect 6562 -16162 6622 -15850
rect 6166 -16222 6176 -16172
rect 6096 -16292 6176 -16222
rect 6096 -16352 6106 -16292
rect 6166 -16352 6176 -16292
rect 6552 -16222 6562 -16172
rect 7020 -16162 7080 -15850
rect 6622 -16222 6632 -16172
rect 6552 -16292 6632 -16222
rect 6552 -16352 6562 -16292
rect 6622 -16352 6632 -16292
rect 7010 -16222 7020 -16172
rect 7476 -16162 7536 -15850
rect 7080 -16222 7090 -16172
rect 7010 -16292 7090 -16222
rect 7010 -16352 7020 -16292
rect 7080 -16352 7090 -16292
rect 7466 -16222 7476 -16172
rect 7932 -16162 7992 -15850
rect 7536 -16222 7546 -16172
rect 7466 -16292 7546 -16222
rect 7466 -16352 7476 -16292
rect 7536 -16352 7546 -16292
rect 7922 -16222 7932 -16172
rect 8406 -16162 8466 -15850
rect 7992 -16222 8002 -16172
rect 7922 -16292 8002 -16222
rect 7922 -16352 7932 -16292
rect 7992 -16352 8002 -16292
rect 8396 -16222 8406 -16172
rect 8862 -16162 8922 -15850
rect 8466 -16222 8476 -16172
rect 8396 -16292 8476 -16222
rect 8396 -16352 8406 -16292
rect 8466 -16352 8476 -16292
rect 8852 -16222 8862 -16172
rect 9320 -16162 9380 -15850
rect 8922 -16222 8932 -16172
rect 8852 -16292 8932 -16222
rect 8852 -16352 8862 -16292
rect 8922 -16352 8932 -16292
rect 9310 -16222 9320 -16172
rect 9776 -16162 9836 -15850
rect 9380 -16222 9390 -16172
rect 9310 -16292 9390 -16222
rect 9310 -16352 9320 -16292
rect 9380 -16352 9390 -16292
rect 9766 -16222 9776 -16172
rect 10232 -16162 10292 -15850
rect 9836 -16222 9846 -16172
rect 9766 -16292 9846 -16222
rect 9766 -16352 9776 -16292
rect 9836 -16352 9846 -16292
rect 10222 -16222 10232 -16172
rect 10690 -16162 10750 -15850
rect 10292 -16222 10302 -16172
rect 10222 -16292 10302 -16222
rect 10222 -16352 10232 -16292
rect 10292 -16352 10302 -16292
rect 10680 -16222 10690 -16172
rect 11146 -16162 11206 -15850
rect 10750 -16222 10760 -16172
rect 10680 -16292 10760 -16222
rect 10680 -16352 10690 -16292
rect 10750 -16352 10760 -16292
rect 11136 -16222 11146 -16172
rect 11602 -16162 11662 -15850
rect 11206 -16222 11216 -16172
rect 11136 -16292 11216 -16222
rect 11136 -16352 11146 -16292
rect 11206 -16352 11216 -16292
rect 11592 -16222 11602 -16172
rect 12060 -16162 12120 -15850
rect 11662 -16222 11672 -16172
rect 11592 -16292 11672 -16222
rect 11592 -16352 11602 -16292
rect 11662 -16352 11672 -16292
rect 12050 -16222 12060 -16172
rect 12516 -16162 12576 -15850
rect 12120 -16222 12130 -16172
rect 12050 -16292 12130 -16222
rect 12050 -16352 12060 -16292
rect 12120 -16352 12130 -16292
rect 12506 -16222 12516 -16172
rect 12972 -16162 13032 -15850
rect 12576 -16222 12586 -16172
rect 12506 -16292 12586 -16222
rect 12506 -16352 12516 -16292
rect 12576 -16352 12586 -16292
rect 12962 -16222 12972 -16172
rect 13430 -16162 13490 -15850
rect 13032 -16222 13042 -16172
rect 12962 -16292 13042 -16222
rect 12962 -16352 12972 -16292
rect 13032 -16352 13042 -16292
rect 13420 -16222 13430 -16172
rect 13886 -16162 13946 -15850
rect 13490 -16222 13500 -16172
rect 13420 -16292 13500 -16222
rect 13420 -16352 13430 -16292
rect 13490 -16352 13500 -16292
rect 13876 -16222 13886 -16172
rect 14342 -16162 14402 -15850
rect 13946 -16222 13956 -16172
rect 13876 -16292 13956 -16222
rect 13876 -16352 13886 -16292
rect 13946 -16352 13956 -16292
rect 14332 -16222 14342 -16172
rect 14800 -16162 14860 -15850
rect 14402 -16222 14412 -16172
rect 14332 -16292 14412 -16222
rect 14332 -16352 14342 -16292
rect 14402 -16352 14412 -16292
rect 14790 -16222 14800 -16172
rect 15256 -16162 15316 -15850
rect 14860 -16222 14870 -16172
rect 14790 -16292 14870 -16222
rect 14790 -16352 14800 -16292
rect 14860 -16352 14870 -16292
rect 15246 -16222 15256 -16172
rect 15316 -16222 15326 -16172
rect 15246 -16292 15326 -16222
rect 15246 -16352 15256 -16292
rect 15316 -16352 15326 -16292
rect 170 -16654 230 -16352
rect 160 -16714 170 -16664
rect 626 -16654 686 -16352
rect 230 -16714 240 -16664
rect 160 -16784 240 -16714
rect 160 -16844 170 -16784
rect 230 -16844 240 -16784
rect 616 -16714 626 -16664
rect 1082 -16654 1142 -16352
rect 686 -16714 696 -16664
rect 616 -16784 696 -16714
rect 616 -16844 626 -16784
rect 686 -16844 696 -16784
rect 1072 -16714 1082 -16664
rect 1540 -16654 1600 -16352
rect 1142 -16714 1152 -16664
rect 1072 -16784 1152 -16714
rect 1072 -16844 1082 -16784
rect 1142 -16844 1152 -16784
rect 1530 -16714 1540 -16664
rect 1996 -16654 2056 -16352
rect 1600 -16714 1610 -16664
rect 1530 -16784 1610 -16714
rect 1530 -16844 1540 -16784
rect 1600 -16844 1610 -16784
rect 1986 -16714 1996 -16664
rect 2452 -16654 2512 -16352
rect 2056 -16714 2066 -16664
rect 1986 -16784 2066 -16714
rect 1986 -16844 1996 -16784
rect 2056 -16844 2066 -16784
rect 2442 -16714 2452 -16664
rect 2910 -16654 2970 -16352
rect 2512 -16714 2522 -16664
rect 2442 -16784 2522 -16714
rect 2442 -16844 2452 -16784
rect 2512 -16844 2522 -16784
rect 2900 -16714 2910 -16664
rect 3366 -16654 3426 -16352
rect 2970 -16714 2980 -16664
rect 2900 -16784 2980 -16714
rect 2900 -16844 2910 -16784
rect 2970 -16844 2980 -16784
rect 3356 -16714 3366 -16664
rect 3822 -16654 3882 -16352
rect 3426 -16714 3436 -16664
rect 3356 -16784 3436 -16714
rect 3356 -16844 3366 -16784
rect 3426 -16844 3436 -16784
rect 3812 -16714 3822 -16664
rect 4280 -16654 4340 -16352
rect 3882 -16714 3892 -16664
rect 3812 -16784 3892 -16714
rect 3812 -16844 3822 -16784
rect 3882 -16844 3892 -16784
rect 4270 -16714 4280 -16664
rect 4736 -16654 4796 -16352
rect 4340 -16714 4350 -16664
rect 4270 -16784 4350 -16714
rect 4270 -16844 4280 -16784
rect 4340 -16844 4350 -16784
rect 4726 -16714 4736 -16664
rect 5192 -16654 5252 -16352
rect 4796 -16714 4806 -16664
rect 4726 -16784 4806 -16714
rect 4726 -16844 4736 -16784
rect 4796 -16844 4806 -16784
rect 5182 -16714 5192 -16664
rect 5650 -16654 5710 -16352
rect 5252 -16714 5262 -16664
rect 5182 -16784 5262 -16714
rect 5182 -16844 5192 -16784
rect 5252 -16844 5262 -16784
rect 5640 -16714 5650 -16664
rect 6106 -16654 6166 -16352
rect 5710 -16714 5720 -16664
rect 5640 -16784 5720 -16714
rect 5640 -16844 5650 -16784
rect 5710 -16844 5720 -16784
rect 6096 -16714 6106 -16664
rect 6562 -16654 6622 -16352
rect 6166 -16714 6176 -16664
rect 6096 -16784 6176 -16714
rect 6096 -16844 6106 -16784
rect 6166 -16844 6176 -16784
rect 6552 -16714 6562 -16664
rect 7020 -16654 7080 -16352
rect 6622 -16714 6632 -16664
rect 6552 -16784 6632 -16714
rect 6552 -16844 6562 -16784
rect 6622 -16844 6632 -16784
rect 7010 -16714 7020 -16664
rect 7476 -16654 7536 -16352
rect 7080 -16714 7090 -16664
rect 7010 -16784 7090 -16714
rect 7010 -16844 7020 -16784
rect 7080 -16844 7090 -16784
rect 7466 -16714 7476 -16664
rect 7932 -16654 7992 -16352
rect 7536 -16714 7546 -16664
rect 7466 -16784 7546 -16714
rect 7466 -16844 7476 -16784
rect 7536 -16844 7546 -16784
rect 7922 -16714 7932 -16664
rect 8406 -16654 8466 -16352
rect 7992 -16714 8002 -16664
rect 7922 -16784 8002 -16714
rect 7922 -16844 7932 -16784
rect 7992 -16844 8002 -16784
rect 8396 -16714 8406 -16664
rect 8862 -16654 8922 -16352
rect 8466 -16714 8476 -16664
rect 8396 -16784 8476 -16714
rect 8396 -16844 8406 -16784
rect 8466 -16844 8476 -16784
rect 8852 -16714 8862 -16664
rect 9320 -16654 9380 -16352
rect 8922 -16714 8932 -16664
rect 8852 -16784 8932 -16714
rect 8852 -16844 8862 -16784
rect 8922 -16844 8932 -16784
rect 9310 -16714 9320 -16664
rect 9776 -16654 9836 -16352
rect 9380 -16714 9390 -16664
rect 9310 -16784 9390 -16714
rect 9310 -16844 9320 -16784
rect 9380 -16844 9390 -16784
rect 9766 -16714 9776 -16664
rect 10232 -16654 10292 -16352
rect 9836 -16714 9846 -16664
rect 9766 -16784 9846 -16714
rect 9766 -16844 9776 -16784
rect 9836 -16844 9846 -16784
rect 10222 -16714 10232 -16664
rect 10690 -16654 10750 -16352
rect 10292 -16714 10302 -16664
rect 10222 -16784 10302 -16714
rect 10222 -16844 10232 -16784
rect 10292 -16844 10302 -16784
rect 10680 -16714 10690 -16664
rect 11146 -16654 11206 -16352
rect 10750 -16714 10760 -16664
rect 10680 -16784 10760 -16714
rect 10680 -16844 10690 -16784
rect 10750 -16844 10760 -16784
rect 11136 -16714 11146 -16664
rect 11602 -16654 11662 -16352
rect 11206 -16714 11216 -16664
rect 11136 -16784 11216 -16714
rect 11136 -16844 11146 -16784
rect 11206 -16844 11216 -16784
rect 11592 -16714 11602 -16664
rect 12060 -16654 12120 -16352
rect 11662 -16714 11672 -16664
rect 11592 -16784 11672 -16714
rect 11592 -16844 11602 -16784
rect 11662 -16844 11672 -16784
rect 12050 -16714 12060 -16664
rect 12516 -16654 12576 -16352
rect 12120 -16714 12130 -16664
rect 12050 -16784 12130 -16714
rect 12050 -16844 12060 -16784
rect 12120 -16844 12130 -16784
rect 12506 -16714 12516 -16664
rect 12972 -16654 13032 -16352
rect 12576 -16714 12586 -16664
rect 12506 -16784 12586 -16714
rect 12506 -16844 12516 -16784
rect 12576 -16844 12586 -16784
rect 12962 -16714 12972 -16664
rect 13430 -16654 13490 -16352
rect 13032 -16714 13042 -16664
rect 12962 -16784 13042 -16714
rect 12962 -16844 12972 -16784
rect 13032 -16844 13042 -16784
rect 13420 -16714 13430 -16664
rect 13886 -16654 13946 -16352
rect 13490 -16714 13500 -16664
rect 13420 -16784 13500 -16714
rect 13420 -16844 13430 -16784
rect 13490 -16844 13500 -16784
rect 13876 -16714 13886 -16664
rect 14342 -16654 14402 -16352
rect 13946 -16714 13956 -16664
rect 13876 -16784 13956 -16714
rect 13876 -16844 13886 -16784
rect 13946 -16844 13956 -16784
rect 14332 -16714 14342 -16664
rect 14800 -16654 14860 -16352
rect 14402 -16714 14412 -16664
rect 14332 -16784 14412 -16714
rect 14332 -16844 14342 -16784
rect 14402 -16844 14412 -16784
rect 14790 -16714 14800 -16664
rect 15256 -16654 15316 -16352
rect 14860 -16714 14870 -16664
rect 14790 -16784 14870 -16714
rect 14790 -16844 14800 -16784
rect 14860 -16844 14870 -16784
rect 15246 -16714 15256 -16664
rect 15316 -16714 15326 -16664
rect 15246 -16784 15326 -16714
rect 15246 -16844 15256 -16784
rect 15316 -16844 15326 -16784
rect 170 -16980 230 -16844
rect 626 -16980 686 -16844
rect 1082 -16980 1142 -16844
rect 1540 -16980 1600 -16844
rect 1996 -16980 2056 -16844
rect 2452 -16980 2512 -16844
rect 2910 -16980 2970 -16844
rect 3366 -16980 3426 -16844
rect 3822 -16980 3882 -16844
rect 4280 -16980 4340 -16844
rect 4736 -16980 4796 -16844
rect 5192 -16980 5252 -16844
rect 5650 -16980 5710 -16844
rect 6106 -16980 6166 -16844
rect 6562 -16980 6622 -16844
rect 7020 -16980 7080 -16844
rect 7476 -16980 7536 -16844
rect 7932 -16980 7992 -16844
rect 8406 -16980 8466 -16844
rect 8862 -16980 8922 -16844
rect 9320 -16980 9380 -16844
rect 9776 -16980 9836 -16844
rect 10232 -16980 10292 -16844
rect 10690 -16980 10750 -16844
rect 11146 -16980 11206 -16844
rect 11602 -16980 11662 -16844
rect 12060 -16980 12120 -16844
rect 12516 -16980 12576 -16844
rect 12972 -16980 13032 -16844
rect 13430 -16980 13490 -16844
rect 13886 -16980 13946 -16844
rect 14342 -16980 14402 -16844
rect 14800 -16980 14860 -16844
rect 15256 -16980 15316 -16844
rect 170 -16984 231 -16980
rect 626 -16984 687 -16980
rect 1082 -16984 1143 -16980
rect 1540 -16984 1601 -16980
rect 1996 -16984 2057 -16980
rect 2452 -16984 2513 -16980
rect 2910 -16984 2971 -16980
rect 3366 -16984 3427 -16980
rect 3822 -16984 3883 -16980
rect 4280 -16984 4341 -16980
rect 4736 -16984 4797 -16980
rect 5192 -16984 5253 -16980
rect 5650 -16984 5711 -16980
rect 6106 -16984 6167 -16980
rect 6562 -16984 6623 -16980
rect 7020 -16984 7081 -16980
rect 7476 -16984 7537 -16980
rect 7932 -16984 7993 -16980
rect 8406 -16984 8467 -16980
rect 8862 -16984 8923 -16980
rect 9320 -16984 9381 -16980
rect 9776 -16984 9837 -16980
rect 10232 -16984 10293 -16980
rect 10690 -16984 10751 -16980
rect 11146 -16984 11207 -16980
rect 11602 -16984 11663 -16980
rect 12060 -16984 12121 -16980
rect 12516 -16984 12577 -16980
rect 12972 -16984 13033 -16980
rect 13430 -16984 13491 -16980
rect 13886 -16984 13947 -16980
rect 14342 -16984 14403 -16980
rect 14800 -16984 14861 -16980
rect 15256 -16984 15317 -16980
rect 171 -17151 231 -16984
rect 161 -17211 171 -17161
rect 627 -17151 687 -16984
rect 231 -17211 241 -17161
rect 161 -17281 241 -17211
rect 161 -17341 171 -17281
rect 231 -17341 241 -17281
rect 617 -17211 627 -17161
rect 1083 -17151 1143 -16984
rect 687 -17211 697 -17161
rect 617 -17281 697 -17211
rect 617 -17341 627 -17281
rect 687 -17341 697 -17281
rect 1073 -17211 1083 -17161
rect 1541 -17151 1601 -16984
rect 1143 -17211 1153 -17161
rect 1073 -17281 1153 -17211
rect 1073 -17341 1083 -17281
rect 1143 -17341 1153 -17281
rect 1531 -17211 1541 -17161
rect 1997 -17151 2057 -16984
rect 1601 -17211 1611 -17161
rect 1531 -17281 1611 -17211
rect 1531 -17341 1541 -17281
rect 1601 -17341 1611 -17281
rect 1987 -17211 1997 -17161
rect 2453 -17151 2513 -16984
rect 2057 -17211 2067 -17161
rect 1987 -17281 2067 -17211
rect 1987 -17341 1997 -17281
rect 2057 -17341 2067 -17281
rect 2443 -17211 2453 -17161
rect 2911 -17151 2971 -16984
rect 2513 -17211 2523 -17161
rect 2443 -17281 2523 -17211
rect 2443 -17341 2453 -17281
rect 2513 -17341 2523 -17281
rect 2901 -17211 2911 -17161
rect 3367 -17151 3427 -16984
rect 2971 -17211 2981 -17161
rect 2901 -17281 2981 -17211
rect 2901 -17341 2911 -17281
rect 2971 -17341 2981 -17281
rect 3357 -17211 3367 -17161
rect 3823 -17151 3883 -16984
rect 3427 -17211 3437 -17161
rect 3357 -17281 3437 -17211
rect 3357 -17341 3367 -17281
rect 3427 -17341 3437 -17281
rect 3813 -17211 3823 -17161
rect 4281 -17151 4341 -16984
rect 3883 -17211 3893 -17161
rect 3813 -17281 3893 -17211
rect 3813 -17341 3823 -17281
rect 3883 -17341 3893 -17281
rect 4271 -17211 4281 -17161
rect 4737 -17151 4797 -16984
rect 4341 -17211 4351 -17161
rect 4271 -17281 4351 -17211
rect 4271 -17341 4281 -17281
rect 4341 -17341 4351 -17281
rect 4727 -17211 4737 -17161
rect 5193 -17151 5253 -16984
rect 4797 -17211 4807 -17161
rect 4727 -17281 4807 -17211
rect 4727 -17341 4737 -17281
rect 4797 -17341 4807 -17281
rect 5183 -17211 5193 -17161
rect 5651 -17151 5711 -16984
rect 5253 -17211 5263 -17161
rect 5183 -17281 5263 -17211
rect 5183 -17341 5193 -17281
rect 5253 -17341 5263 -17281
rect 5641 -17211 5651 -17161
rect 6107 -17151 6167 -16984
rect 5711 -17211 5721 -17161
rect 5641 -17281 5721 -17211
rect 5641 -17341 5651 -17281
rect 5711 -17341 5721 -17281
rect 6097 -17211 6107 -17161
rect 6563 -17151 6623 -16984
rect 6167 -17211 6177 -17161
rect 6097 -17281 6177 -17211
rect 6097 -17341 6107 -17281
rect 6167 -17341 6177 -17281
rect 6553 -17211 6563 -17161
rect 7021 -17151 7081 -16984
rect 6623 -17211 6633 -17161
rect 6553 -17281 6633 -17211
rect 6553 -17341 6563 -17281
rect 6623 -17341 6633 -17281
rect 7011 -17211 7021 -17161
rect 7477 -17151 7537 -16984
rect 7081 -17211 7091 -17161
rect 7011 -17281 7091 -17211
rect 7011 -17341 7021 -17281
rect 7081 -17341 7091 -17281
rect 7467 -17211 7477 -17161
rect 7933 -17151 7993 -16984
rect 7537 -17211 7547 -17161
rect 7467 -17281 7547 -17211
rect 7467 -17341 7477 -17281
rect 7537 -17341 7547 -17281
rect 7923 -17211 7933 -17161
rect 8407 -17151 8467 -16984
rect 7993 -17211 8003 -17161
rect 7923 -17281 8003 -17211
rect 7923 -17341 7933 -17281
rect 7993 -17341 8003 -17281
rect 8397 -17211 8407 -17161
rect 8863 -17151 8923 -16984
rect 8467 -17211 8477 -17161
rect 8397 -17281 8477 -17211
rect 8397 -17341 8407 -17281
rect 8467 -17341 8477 -17281
rect 8853 -17211 8863 -17161
rect 9321 -17151 9381 -16984
rect 8923 -17211 8933 -17161
rect 8853 -17281 8933 -17211
rect 8853 -17341 8863 -17281
rect 8923 -17341 8933 -17281
rect 9311 -17211 9321 -17161
rect 9777 -17151 9837 -16984
rect 9381 -17211 9391 -17161
rect 9311 -17281 9391 -17211
rect 9311 -17341 9321 -17281
rect 9381 -17341 9391 -17281
rect 9767 -17211 9777 -17161
rect 10233 -17151 10293 -16984
rect 9837 -17211 9847 -17161
rect 9767 -17281 9847 -17211
rect 9767 -17341 9777 -17281
rect 9837 -17341 9847 -17281
rect 10223 -17211 10233 -17161
rect 10691 -17151 10751 -16984
rect 10293 -17211 10303 -17161
rect 10223 -17281 10303 -17211
rect 10223 -17341 10233 -17281
rect 10293 -17341 10303 -17281
rect 10681 -17211 10691 -17161
rect 11147 -17151 11207 -16984
rect 10751 -17211 10761 -17161
rect 10681 -17281 10761 -17211
rect 10681 -17341 10691 -17281
rect 10751 -17341 10761 -17281
rect 11137 -17211 11147 -17161
rect 11603 -17151 11663 -16984
rect 11207 -17211 11217 -17161
rect 11137 -17281 11217 -17211
rect 11137 -17341 11147 -17281
rect 11207 -17341 11217 -17281
rect 11593 -17211 11603 -17161
rect 12061 -17151 12121 -16984
rect 11663 -17211 11673 -17161
rect 11593 -17281 11673 -17211
rect 11593 -17341 11603 -17281
rect 11663 -17341 11673 -17281
rect 12051 -17211 12061 -17161
rect 12517 -17151 12577 -16984
rect 12121 -17211 12131 -17161
rect 12051 -17281 12131 -17211
rect 12051 -17341 12061 -17281
rect 12121 -17341 12131 -17281
rect 12507 -17211 12517 -17161
rect 12973 -17151 13033 -16984
rect 12577 -17211 12587 -17161
rect 12507 -17281 12587 -17211
rect 12507 -17341 12517 -17281
rect 12577 -17341 12587 -17281
rect 12963 -17211 12973 -17161
rect 13431 -17151 13491 -16984
rect 13033 -17211 13043 -17161
rect 12963 -17281 13043 -17211
rect 12963 -17341 12973 -17281
rect 13033 -17341 13043 -17281
rect 13421 -17211 13431 -17161
rect 13887 -17151 13947 -16984
rect 13491 -17211 13501 -17161
rect 13421 -17281 13501 -17211
rect 13421 -17341 13431 -17281
rect 13491 -17341 13501 -17281
rect 13877 -17211 13887 -17161
rect 14343 -17151 14403 -16984
rect 13947 -17211 13957 -17161
rect 13877 -17281 13957 -17211
rect 13877 -17341 13887 -17281
rect 13947 -17341 13957 -17281
rect 14333 -17211 14343 -17161
rect 14801 -17151 14861 -16984
rect 14403 -17211 14413 -17161
rect 14333 -17281 14413 -17211
rect 14333 -17341 14343 -17281
rect 14403 -17341 14413 -17281
rect 14791 -17211 14801 -17161
rect 15257 -17151 15317 -16984
rect 14861 -17211 14871 -17161
rect 14791 -17281 14871 -17211
rect 14791 -17341 14801 -17281
rect 14861 -17341 14871 -17281
rect 15247 -17211 15257 -17161
rect 15317 -17211 15327 -17161
rect 15247 -17281 15327 -17211
rect 15247 -17341 15257 -17281
rect 15317 -17341 15327 -17281
rect 171 -17643 231 -17341
rect 161 -17703 171 -17653
rect 627 -17643 687 -17341
rect 231 -17703 241 -17653
rect 161 -17773 241 -17703
rect 161 -17833 171 -17773
rect 231 -17833 241 -17773
rect 617 -17703 627 -17653
rect 1083 -17643 1143 -17341
rect 687 -17703 697 -17653
rect 617 -17773 697 -17703
rect 617 -17833 627 -17773
rect 687 -17833 697 -17773
rect 1073 -17703 1083 -17653
rect 1541 -17643 1601 -17341
rect 1143 -17703 1153 -17653
rect 1073 -17773 1153 -17703
rect 1073 -17833 1083 -17773
rect 1143 -17833 1153 -17773
rect 1531 -17703 1541 -17653
rect 1997 -17643 2057 -17341
rect 1601 -17703 1611 -17653
rect 1531 -17773 1611 -17703
rect 1531 -17833 1541 -17773
rect 1601 -17833 1611 -17773
rect 1987 -17703 1997 -17653
rect 2453 -17643 2513 -17341
rect 2057 -17703 2067 -17653
rect 1987 -17773 2067 -17703
rect 1987 -17833 1997 -17773
rect 2057 -17833 2067 -17773
rect 2443 -17703 2453 -17653
rect 2911 -17643 2971 -17341
rect 2513 -17703 2523 -17653
rect 2443 -17773 2523 -17703
rect 2443 -17833 2453 -17773
rect 2513 -17833 2523 -17773
rect 2901 -17703 2911 -17653
rect 3367 -17643 3427 -17341
rect 2971 -17703 2981 -17653
rect 2901 -17773 2981 -17703
rect 2901 -17833 2911 -17773
rect 2971 -17833 2981 -17773
rect 3357 -17703 3367 -17653
rect 3823 -17643 3883 -17341
rect 3427 -17703 3437 -17653
rect 3357 -17773 3437 -17703
rect 3357 -17833 3367 -17773
rect 3427 -17833 3437 -17773
rect 3813 -17703 3823 -17653
rect 4281 -17643 4341 -17341
rect 3883 -17703 3893 -17653
rect 3813 -17773 3893 -17703
rect 3813 -17833 3823 -17773
rect 3883 -17833 3893 -17773
rect 4271 -17703 4281 -17653
rect 4737 -17643 4797 -17341
rect 4341 -17703 4351 -17653
rect 4271 -17773 4351 -17703
rect 4271 -17833 4281 -17773
rect 4341 -17833 4351 -17773
rect 4727 -17703 4737 -17653
rect 5193 -17643 5253 -17341
rect 4797 -17703 4807 -17653
rect 4727 -17773 4807 -17703
rect 4727 -17833 4737 -17773
rect 4797 -17833 4807 -17773
rect 5183 -17703 5193 -17653
rect 5651 -17643 5711 -17341
rect 5253 -17703 5263 -17653
rect 5183 -17773 5263 -17703
rect 5183 -17833 5193 -17773
rect 5253 -17833 5263 -17773
rect 5641 -17703 5651 -17653
rect 6107 -17643 6167 -17341
rect 5711 -17703 5721 -17653
rect 5641 -17773 5721 -17703
rect 5641 -17833 5651 -17773
rect 5711 -17833 5721 -17773
rect 6097 -17703 6107 -17653
rect 6563 -17643 6623 -17341
rect 6167 -17703 6177 -17653
rect 6097 -17773 6177 -17703
rect 6097 -17833 6107 -17773
rect 6167 -17833 6177 -17773
rect 6553 -17703 6563 -17653
rect 7021 -17643 7081 -17341
rect 6623 -17703 6633 -17653
rect 6553 -17773 6633 -17703
rect 6553 -17833 6563 -17773
rect 6623 -17833 6633 -17773
rect 7011 -17703 7021 -17653
rect 7477 -17643 7537 -17341
rect 7081 -17703 7091 -17653
rect 7011 -17773 7091 -17703
rect 7011 -17833 7021 -17773
rect 7081 -17833 7091 -17773
rect 7467 -17703 7477 -17653
rect 7933 -17643 7993 -17341
rect 7537 -17703 7547 -17653
rect 7467 -17773 7547 -17703
rect 7467 -17833 7477 -17773
rect 7537 -17833 7547 -17773
rect 7923 -17703 7933 -17653
rect 8407 -17643 8467 -17341
rect 7993 -17703 8003 -17653
rect 7923 -17773 8003 -17703
rect 7923 -17833 7933 -17773
rect 7993 -17833 8003 -17773
rect 8397 -17703 8407 -17653
rect 8863 -17643 8923 -17341
rect 8467 -17703 8477 -17653
rect 8397 -17773 8477 -17703
rect 8397 -17833 8407 -17773
rect 8467 -17833 8477 -17773
rect 8853 -17703 8863 -17653
rect 9321 -17643 9381 -17341
rect 8923 -17703 8933 -17653
rect 8853 -17773 8933 -17703
rect 8853 -17833 8863 -17773
rect 8923 -17833 8933 -17773
rect 9311 -17703 9321 -17653
rect 9777 -17643 9837 -17341
rect 9381 -17703 9391 -17653
rect 9311 -17773 9391 -17703
rect 9311 -17833 9321 -17773
rect 9381 -17833 9391 -17773
rect 9767 -17703 9777 -17653
rect 10233 -17643 10293 -17341
rect 9837 -17703 9847 -17653
rect 9767 -17773 9847 -17703
rect 9767 -17833 9777 -17773
rect 9837 -17833 9847 -17773
rect 10223 -17703 10233 -17653
rect 10691 -17643 10751 -17341
rect 10293 -17703 10303 -17653
rect 10223 -17773 10303 -17703
rect 10223 -17833 10233 -17773
rect 10293 -17833 10303 -17773
rect 10681 -17703 10691 -17653
rect 11147 -17643 11207 -17341
rect 10751 -17703 10761 -17653
rect 10681 -17773 10761 -17703
rect 10681 -17833 10691 -17773
rect 10751 -17833 10761 -17773
rect 11137 -17703 11147 -17653
rect 11603 -17643 11663 -17341
rect 11207 -17703 11217 -17653
rect 11137 -17773 11217 -17703
rect 11137 -17833 11147 -17773
rect 11207 -17833 11217 -17773
rect 11593 -17703 11603 -17653
rect 12061 -17643 12121 -17341
rect 11663 -17703 11673 -17653
rect 11593 -17773 11673 -17703
rect 11593 -17833 11603 -17773
rect 11663 -17833 11673 -17773
rect 12051 -17703 12061 -17653
rect 12517 -17643 12577 -17341
rect 12121 -17703 12131 -17653
rect 12051 -17773 12131 -17703
rect 12051 -17833 12061 -17773
rect 12121 -17833 12131 -17773
rect 12507 -17703 12517 -17653
rect 12973 -17643 13033 -17341
rect 12577 -17703 12587 -17653
rect 12507 -17773 12587 -17703
rect 12507 -17833 12517 -17773
rect 12577 -17833 12587 -17773
rect 12963 -17703 12973 -17653
rect 13431 -17643 13491 -17341
rect 13033 -17703 13043 -17653
rect 12963 -17773 13043 -17703
rect 12963 -17833 12973 -17773
rect 13033 -17833 13043 -17773
rect 13421 -17703 13431 -17653
rect 13887 -17643 13947 -17341
rect 13491 -17703 13501 -17653
rect 13421 -17773 13501 -17703
rect 13421 -17833 13431 -17773
rect 13491 -17833 13501 -17773
rect 13877 -17703 13887 -17653
rect 14343 -17643 14403 -17341
rect 13947 -17703 13957 -17653
rect 13877 -17773 13957 -17703
rect 13877 -17833 13887 -17773
rect 13947 -17833 13957 -17773
rect 14333 -17703 14343 -17653
rect 14801 -17643 14861 -17341
rect 14403 -17703 14413 -17653
rect 14333 -17773 14413 -17703
rect 14333 -17833 14343 -17773
rect 14403 -17833 14413 -17773
rect 14791 -17703 14801 -17653
rect 15257 -17643 15317 -17341
rect 14861 -17703 14871 -17653
rect 14791 -17773 14871 -17703
rect 14791 -17833 14801 -17773
rect 14861 -17833 14871 -17773
rect 15247 -17703 15257 -17653
rect 15317 -17703 15327 -17653
rect 15247 -17773 15327 -17703
rect 15247 -17833 15257 -17773
rect 15317 -17833 15327 -17773
rect 171 -18159 231 -17833
rect 161 -18219 171 -18169
rect 627 -18159 687 -17833
rect 231 -18219 241 -18169
rect 161 -18289 241 -18219
rect 161 -18349 171 -18289
rect 231 -18349 241 -18289
rect 617 -18219 627 -18169
rect 1083 -18159 1143 -17833
rect 687 -18219 697 -18169
rect 617 -18289 697 -18219
rect 617 -18349 627 -18289
rect 687 -18349 697 -18289
rect 1073 -18219 1083 -18169
rect 1541 -18159 1601 -17833
rect 1143 -18219 1153 -18169
rect 1073 -18289 1153 -18219
rect 1073 -18349 1083 -18289
rect 1143 -18349 1153 -18289
rect 1531 -18219 1541 -18169
rect 1997 -18159 2057 -17833
rect 1601 -18219 1611 -18169
rect 1531 -18289 1611 -18219
rect 1531 -18349 1541 -18289
rect 1601 -18349 1611 -18289
rect 1987 -18219 1997 -18169
rect 2453 -18159 2513 -17833
rect 2057 -18219 2067 -18169
rect 1987 -18289 2067 -18219
rect 1987 -18349 1997 -18289
rect 2057 -18349 2067 -18289
rect 2443 -18219 2453 -18169
rect 2911 -18159 2971 -17833
rect 2513 -18219 2523 -18169
rect 2443 -18289 2523 -18219
rect 2443 -18349 2453 -18289
rect 2513 -18349 2523 -18289
rect 2901 -18219 2911 -18169
rect 3367 -18159 3427 -17833
rect 2971 -18219 2981 -18169
rect 2901 -18289 2981 -18219
rect 2901 -18349 2911 -18289
rect 2971 -18349 2981 -18289
rect 3357 -18219 3367 -18169
rect 3823 -18159 3883 -17833
rect 3427 -18219 3437 -18169
rect 3357 -18289 3437 -18219
rect 3357 -18349 3367 -18289
rect 3427 -18349 3437 -18289
rect 3813 -18219 3823 -18169
rect 4281 -18159 4341 -17833
rect 3883 -18219 3893 -18169
rect 3813 -18289 3893 -18219
rect 3813 -18349 3823 -18289
rect 3883 -18349 3893 -18289
rect 4271 -18219 4281 -18169
rect 4737 -18159 4797 -17833
rect 4341 -18219 4351 -18169
rect 4271 -18289 4351 -18219
rect 4271 -18349 4281 -18289
rect 4341 -18349 4351 -18289
rect 4727 -18219 4737 -18169
rect 5193 -18159 5253 -17833
rect 4797 -18219 4807 -18169
rect 4727 -18289 4807 -18219
rect 4727 -18349 4737 -18289
rect 4797 -18349 4807 -18289
rect 5183 -18219 5193 -18169
rect 5651 -18159 5711 -17833
rect 5253 -18219 5263 -18169
rect 5183 -18289 5263 -18219
rect 5183 -18349 5193 -18289
rect 5253 -18349 5263 -18289
rect 5641 -18219 5651 -18169
rect 6107 -18159 6167 -17833
rect 5711 -18219 5721 -18169
rect 5641 -18289 5721 -18219
rect 5641 -18349 5651 -18289
rect 5711 -18349 5721 -18289
rect 6097 -18219 6107 -18169
rect 6563 -18159 6623 -17833
rect 6167 -18219 6177 -18169
rect 6097 -18289 6177 -18219
rect 6097 -18349 6107 -18289
rect 6167 -18349 6177 -18289
rect 6553 -18219 6563 -18169
rect 7021 -18159 7081 -17833
rect 6623 -18219 6633 -18169
rect 6553 -18289 6633 -18219
rect 6553 -18349 6563 -18289
rect 6623 -18349 6633 -18289
rect 7011 -18219 7021 -18169
rect 7477 -18159 7537 -17833
rect 7081 -18219 7091 -18169
rect 7011 -18289 7091 -18219
rect 7011 -18349 7021 -18289
rect 7081 -18349 7091 -18289
rect 7467 -18219 7477 -18169
rect 7933 -18159 7993 -17833
rect 7537 -18219 7547 -18169
rect 7467 -18289 7547 -18219
rect 7467 -18349 7477 -18289
rect 7537 -18349 7547 -18289
rect 7923 -18219 7933 -18169
rect 8407 -18159 8467 -17833
rect 7993 -18219 8003 -18169
rect 7923 -18289 8003 -18219
rect 7923 -18349 7933 -18289
rect 7993 -18349 8003 -18289
rect 8397 -18219 8407 -18169
rect 8863 -18159 8923 -17833
rect 8467 -18219 8477 -18169
rect 8397 -18289 8477 -18219
rect 8397 -18349 8407 -18289
rect 8467 -18349 8477 -18289
rect 8853 -18219 8863 -18169
rect 9321 -18159 9381 -17833
rect 8923 -18219 8933 -18169
rect 8853 -18289 8933 -18219
rect 8853 -18349 8863 -18289
rect 8923 -18349 8933 -18289
rect 9311 -18219 9321 -18169
rect 9777 -18159 9837 -17833
rect 9381 -18219 9391 -18169
rect 9311 -18289 9391 -18219
rect 9311 -18349 9321 -18289
rect 9381 -18349 9391 -18289
rect 9767 -18219 9777 -18169
rect 10233 -18159 10293 -17833
rect 9837 -18219 9847 -18169
rect 9767 -18289 9847 -18219
rect 9767 -18349 9777 -18289
rect 9837 -18349 9847 -18289
rect 10223 -18219 10233 -18169
rect 10691 -18159 10751 -17833
rect 10293 -18219 10303 -18169
rect 10223 -18289 10303 -18219
rect 10223 -18349 10233 -18289
rect 10293 -18349 10303 -18289
rect 10681 -18219 10691 -18169
rect 11147 -18159 11207 -17833
rect 10751 -18219 10761 -18169
rect 10681 -18289 10761 -18219
rect 10681 -18349 10691 -18289
rect 10751 -18349 10761 -18289
rect 11137 -18219 11147 -18169
rect 11603 -18159 11663 -17833
rect 11207 -18219 11217 -18169
rect 11137 -18289 11217 -18219
rect 11137 -18349 11147 -18289
rect 11207 -18349 11217 -18289
rect 11593 -18219 11603 -18169
rect 12061 -18159 12121 -17833
rect 11663 -18219 11673 -18169
rect 11593 -18289 11673 -18219
rect 11593 -18349 11603 -18289
rect 11663 -18349 11673 -18289
rect 12051 -18219 12061 -18169
rect 12517 -18159 12577 -17833
rect 12121 -18219 12131 -18169
rect 12051 -18289 12131 -18219
rect 12051 -18349 12061 -18289
rect 12121 -18349 12131 -18289
rect 12507 -18219 12517 -18169
rect 12973 -18159 13033 -17833
rect 12577 -18219 12587 -18169
rect 12507 -18289 12587 -18219
rect 12507 -18349 12517 -18289
rect 12577 -18349 12587 -18289
rect 12963 -18219 12973 -18169
rect 13431 -18159 13491 -17833
rect 13033 -18219 13043 -18169
rect 12963 -18289 13043 -18219
rect 12963 -18349 12973 -18289
rect 13033 -18349 13043 -18289
rect 13421 -18219 13431 -18169
rect 13887 -18159 13947 -17833
rect 13491 -18219 13501 -18169
rect 13421 -18289 13501 -18219
rect 13421 -18349 13431 -18289
rect 13491 -18349 13501 -18289
rect 13877 -18219 13887 -18169
rect 14343 -18159 14403 -17833
rect 13947 -18219 13957 -18169
rect 13877 -18289 13957 -18219
rect 13877 -18349 13887 -18289
rect 13947 -18349 13957 -18289
rect 14333 -18219 14343 -18169
rect 14801 -18159 14861 -17833
rect 14403 -18219 14413 -18169
rect 14333 -18289 14413 -18219
rect 14333 -18349 14343 -18289
rect 14403 -18349 14413 -18289
rect 14791 -18219 14801 -18169
rect 15257 -18159 15317 -17833
rect 14861 -18219 14871 -18169
rect 14791 -18289 14871 -18219
rect 14791 -18349 14801 -18289
rect 14861 -18349 14871 -18289
rect 15247 -18219 15257 -18169
rect 15317 -18219 15327 -18169
rect 15247 -18289 15327 -18219
rect 15247 -18349 15257 -18289
rect 15317 -18349 15327 -18289
rect 171 -18661 231 -18349
rect 161 -18721 171 -18671
rect 627 -18661 687 -18349
rect 231 -18721 241 -18671
rect 161 -18791 241 -18721
rect 161 -18851 171 -18791
rect 231 -18851 241 -18791
rect 617 -18721 627 -18671
rect 1083 -18661 1143 -18349
rect 687 -18721 697 -18671
rect 617 -18791 697 -18721
rect 617 -18851 627 -18791
rect 687 -18851 697 -18791
rect 1073 -18721 1083 -18671
rect 1541 -18661 1601 -18349
rect 1143 -18721 1153 -18671
rect 1073 -18791 1153 -18721
rect 1073 -18851 1083 -18791
rect 1143 -18851 1153 -18791
rect 1531 -18721 1541 -18671
rect 1997 -18661 2057 -18349
rect 1601 -18721 1611 -18671
rect 1531 -18791 1611 -18721
rect 1531 -18851 1541 -18791
rect 1601 -18851 1611 -18791
rect 1987 -18721 1997 -18671
rect 2453 -18661 2513 -18349
rect 2057 -18721 2067 -18671
rect 1987 -18791 2067 -18721
rect 1987 -18851 1997 -18791
rect 2057 -18851 2067 -18791
rect 2443 -18721 2453 -18671
rect 2911 -18661 2971 -18349
rect 2513 -18721 2523 -18671
rect 2443 -18791 2523 -18721
rect 2443 -18851 2453 -18791
rect 2513 -18851 2523 -18791
rect 2901 -18721 2911 -18671
rect 3367 -18661 3427 -18349
rect 2971 -18721 2981 -18671
rect 2901 -18791 2981 -18721
rect 2901 -18851 2911 -18791
rect 2971 -18851 2981 -18791
rect 3357 -18721 3367 -18671
rect 3823 -18661 3883 -18349
rect 3427 -18721 3437 -18671
rect 3357 -18791 3437 -18721
rect 3357 -18851 3367 -18791
rect 3427 -18851 3437 -18791
rect 3813 -18721 3823 -18671
rect 4281 -18661 4341 -18349
rect 3883 -18721 3893 -18671
rect 3813 -18791 3893 -18721
rect 3813 -18851 3823 -18791
rect 3883 -18851 3893 -18791
rect 4271 -18721 4281 -18671
rect 4737 -18661 4797 -18349
rect 4341 -18721 4351 -18671
rect 4271 -18791 4351 -18721
rect 4271 -18851 4281 -18791
rect 4341 -18851 4351 -18791
rect 4727 -18721 4737 -18671
rect 5193 -18661 5253 -18349
rect 4797 -18721 4807 -18671
rect 4727 -18791 4807 -18721
rect 4727 -18851 4737 -18791
rect 4797 -18851 4807 -18791
rect 5183 -18721 5193 -18671
rect 5651 -18661 5711 -18349
rect 5253 -18721 5263 -18671
rect 5183 -18791 5263 -18721
rect 5183 -18851 5193 -18791
rect 5253 -18851 5263 -18791
rect 5641 -18721 5651 -18671
rect 6107 -18661 6167 -18349
rect 5711 -18721 5721 -18671
rect 5641 -18791 5721 -18721
rect 5641 -18851 5651 -18791
rect 5711 -18851 5721 -18791
rect 6097 -18721 6107 -18671
rect 6563 -18661 6623 -18349
rect 6167 -18721 6177 -18671
rect 6097 -18791 6177 -18721
rect 6097 -18851 6107 -18791
rect 6167 -18851 6177 -18791
rect 6553 -18721 6563 -18671
rect 7021 -18661 7081 -18349
rect 6623 -18721 6633 -18671
rect 6553 -18791 6633 -18721
rect 6553 -18851 6563 -18791
rect 6623 -18851 6633 -18791
rect 7011 -18721 7021 -18671
rect 7477 -18661 7537 -18349
rect 7081 -18721 7091 -18671
rect 7011 -18791 7091 -18721
rect 7011 -18851 7021 -18791
rect 7081 -18851 7091 -18791
rect 7467 -18721 7477 -18671
rect 7933 -18661 7993 -18349
rect 7537 -18721 7547 -18671
rect 7467 -18791 7547 -18721
rect 7467 -18851 7477 -18791
rect 7537 -18851 7547 -18791
rect 7923 -18721 7933 -18671
rect 8407 -18661 8467 -18349
rect 7993 -18721 8003 -18671
rect 7923 -18791 8003 -18721
rect 7923 -18851 7933 -18791
rect 7993 -18851 8003 -18791
rect 8397 -18721 8407 -18671
rect 8863 -18661 8923 -18349
rect 8467 -18721 8477 -18671
rect 8397 -18791 8477 -18721
rect 8397 -18851 8407 -18791
rect 8467 -18851 8477 -18791
rect 8853 -18721 8863 -18671
rect 9321 -18661 9381 -18349
rect 8923 -18721 8933 -18671
rect 8853 -18791 8933 -18721
rect 8853 -18851 8863 -18791
rect 8923 -18851 8933 -18791
rect 9311 -18721 9321 -18671
rect 9777 -18661 9837 -18349
rect 9381 -18721 9391 -18671
rect 9311 -18791 9391 -18721
rect 9311 -18851 9321 -18791
rect 9381 -18851 9391 -18791
rect 9767 -18721 9777 -18671
rect 10233 -18661 10293 -18349
rect 9837 -18721 9847 -18671
rect 9767 -18791 9847 -18721
rect 9767 -18851 9777 -18791
rect 9837 -18851 9847 -18791
rect 10223 -18721 10233 -18671
rect 10691 -18661 10751 -18349
rect 10293 -18721 10303 -18671
rect 10223 -18791 10303 -18721
rect 10223 -18851 10233 -18791
rect 10293 -18851 10303 -18791
rect 10681 -18721 10691 -18671
rect 11147 -18661 11207 -18349
rect 10751 -18721 10761 -18671
rect 10681 -18791 10761 -18721
rect 10681 -18851 10691 -18791
rect 10751 -18851 10761 -18791
rect 11137 -18721 11147 -18671
rect 11603 -18661 11663 -18349
rect 11207 -18721 11217 -18671
rect 11137 -18791 11217 -18721
rect 11137 -18851 11147 -18791
rect 11207 -18851 11217 -18791
rect 11593 -18721 11603 -18671
rect 12061 -18661 12121 -18349
rect 11663 -18721 11673 -18671
rect 11593 -18791 11673 -18721
rect 11593 -18851 11603 -18791
rect 11663 -18851 11673 -18791
rect 12051 -18721 12061 -18671
rect 12517 -18661 12577 -18349
rect 12121 -18721 12131 -18671
rect 12051 -18791 12131 -18721
rect 12051 -18851 12061 -18791
rect 12121 -18851 12131 -18791
rect 12507 -18721 12517 -18671
rect 12973 -18661 13033 -18349
rect 12577 -18721 12587 -18671
rect 12507 -18791 12587 -18721
rect 12507 -18851 12517 -18791
rect 12577 -18851 12587 -18791
rect 12963 -18721 12973 -18671
rect 13431 -18661 13491 -18349
rect 13033 -18721 13043 -18671
rect 12963 -18791 13043 -18721
rect 12963 -18851 12973 -18791
rect 13033 -18851 13043 -18791
rect 13421 -18721 13431 -18671
rect 13887 -18661 13947 -18349
rect 13491 -18721 13501 -18671
rect 13421 -18791 13501 -18721
rect 13421 -18851 13431 -18791
rect 13491 -18851 13501 -18791
rect 13877 -18721 13887 -18671
rect 14343 -18661 14403 -18349
rect 13947 -18721 13957 -18671
rect 13877 -18791 13957 -18721
rect 13877 -18851 13887 -18791
rect 13947 -18851 13957 -18791
rect 14333 -18721 14343 -18671
rect 14801 -18661 14861 -18349
rect 14403 -18721 14413 -18671
rect 14333 -18791 14413 -18721
rect 14333 -18851 14343 -18791
rect 14403 -18851 14413 -18791
rect 14791 -18721 14801 -18671
rect 15257 -18661 15317 -18349
rect 14861 -18721 14871 -18671
rect 14791 -18791 14871 -18721
rect 14791 -18851 14801 -18791
rect 14861 -18851 14871 -18791
rect 15247 -18721 15257 -18671
rect 15317 -18721 15327 -18671
rect 15247 -18791 15327 -18721
rect 15247 -18851 15257 -18791
rect 15317 -18851 15327 -18791
rect 171 -19153 231 -18851
rect 161 -19213 171 -19163
rect 627 -19153 687 -18851
rect 231 -19213 241 -19163
rect 161 -19283 241 -19213
rect 161 -19343 171 -19283
rect 231 -19343 241 -19283
rect 617 -19213 627 -19163
rect 1083 -19153 1143 -18851
rect 687 -19213 697 -19163
rect 617 -19283 697 -19213
rect 617 -19343 627 -19283
rect 687 -19343 697 -19283
rect 1073 -19213 1083 -19163
rect 1541 -19153 1601 -18851
rect 1143 -19213 1153 -19163
rect 1073 -19283 1153 -19213
rect 1073 -19343 1083 -19283
rect 1143 -19343 1153 -19283
rect 1531 -19213 1541 -19163
rect 1997 -19153 2057 -18851
rect 1601 -19213 1611 -19163
rect 1531 -19283 1611 -19213
rect 1531 -19343 1541 -19283
rect 1601 -19343 1611 -19283
rect 1987 -19213 1997 -19163
rect 2453 -19153 2513 -18851
rect 2057 -19213 2067 -19163
rect 1987 -19283 2067 -19213
rect 1987 -19343 1997 -19283
rect 2057 -19343 2067 -19283
rect 2443 -19213 2453 -19163
rect 2911 -19153 2971 -18851
rect 2513 -19213 2523 -19163
rect 2443 -19283 2523 -19213
rect 2443 -19343 2453 -19283
rect 2513 -19343 2523 -19283
rect 2901 -19213 2911 -19163
rect 3367 -19153 3427 -18851
rect 2971 -19213 2981 -19163
rect 2901 -19283 2981 -19213
rect 2901 -19343 2911 -19283
rect 2971 -19343 2981 -19283
rect 3357 -19213 3367 -19163
rect 3823 -19153 3883 -18851
rect 3427 -19213 3437 -19163
rect 3357 -19283 3437 -19213
rect 3357 -19343 3367 -19283
rect 3427 -19343 3437 -19283
rect 3813 -19213 3823 -19163
rect 4281 -19153 4341 -18851
rect 3883 -19213 3893 -19163
rect 3813 -19283 3893 -19213
rect 3813 -19343 3823 -19283
rect 3883 -19343 3893 -19283
rect 4271 -19213 4281 -19163
rect 4737 -19153 4797 -18851
rect 4341 -19213 4351 -19163
rect 4271 -19283 4351 -19213
rect 4271 -19343 4281 -19283
rect 4341 -19343 4351 -19283
rect 4727 -19213 4737 -19163
rect 5193 -19153 5253 -18851
rect 4797 -19213 4807 -19163
rect 4727 -19283 4807 -19213
rect 4727 -19343 4737 -19283
rect 4797 -19343 4807 -19283
rect 5183 -19213 5193 -19163
rect 5651 -19153 5711 -18851
rect 5253 -19213 5263 -19163
rect 5183 -19283 5263 -19213
rect 5183 -19343 5193 -19283
rect 5253 -19343 5263 -19283
rect 5641 -19213 5651 -19163
rect 6107 -19153 6167 -18851
rect 5711 -19213 5721 -19163
rect 5641 -19283 5721 -19213
rect 5641 -19343 5651 -19283
rect 5711 -19343 5721 -19283
rect 6097 -19213 6107 -19163
rect 6563 -19153 6623 -18851
rect 6167 -19213 6177 -19163
rect 6097 -19283 6177 -19213
rect 6097 -19343 6107 -19283
rect 6167 -19343 6177 -19283
rect 6553 -19213 6563 -19163
rect 7021 -19153 7081 -18851
rect 6623 -19213 6633 -19163
rect 6553 -19283 6633 -19213
rect 6553 -19343 6563 -19283
rect 6623 -19343 6633 -19283
rect 7011 -19213 7021 -19163
rect 7477 -19153 7537 -18851
rect 7081 -19213 7091 -19163
rect 7011 -19283 7091 -19213
rect 7011 -19343 7021 -19283
rect 7081 -19343 7091 -19283
rect 7467 -19213 7477 -19163
rect 7933 -19153 7993 -18851
rect 7537 -19213 7547 -19163
rect 7467 -19283 7547 -19213
rect 7467 -19343 7477 -19283
rect 7537 -19343 7547 -19283
rect 7923 -19213 7933 -19163
rect 8407 -19153 8467 -18851
rect 7993 -19213 8003 -19163
rect 7923 -19283 8003 -19213
rect 7923 -19343 7933 -19283
rect 7993 -19343 8003 -19283
rect 8397 -19213 8407 -19163
rect 8863 -19153 8923 -18851
rect 8467 -19213 8477 -19163
rect 8397 -19283 8477 -19213
rect 8397 -19343 8407 -19283
rect 8467 -19343 8477 -19283
rect 8853 -19213 8863 -19163
rect 9321 -19153 9381 -18851
rect 8923 -19213 8933 -19163
rect 8853 -19283 8933 -19213
rect 8853 -19343 8863 -19283
rect 8923 -19343 8933 -19283
rect 9311 -19213 9321 -19163
rect 9777 -19153 9837 -18851
rect 9381 -19213 9391 -19163
rect 9311 -19283 9391 -19213
rect 9311 -19343 9321 -19283
rect 9381 -19343 9391 -19283
rect 9767 -19213 9777 -19163
rect 10233 -19153 10293 -18851
rect 9837 -19213 9847 -19163
rect 9767 -19283 9847 -19213
rect 9767 -19343 9777 -19283
rect 9837 -19343 9847 -19283
rect 10223 -19213 10233 -19163
rect 10691 -19153 10751 -18851
rect 10293 -19213 10303 -19163
rect 10223 -19283 10303 -19213
rect 10223 -19343 10233 -19283
rect 10293 -19343 10303 -19283
rect 10681 -19213 10691 -19163
rect 11147 -19153 11207 -18851
rect 10751 -19213 10761 -19163
rect 10681 -19283 10761 -19213
rect 10681 -19343 10691 -19283
rect 10751 -19343 10761 -19283
rect 11137 -19213 11147 -19163
rect 11603 -19153 11663 -18851
rect 11207 -19213 11217 -19163
rect 11137 -19283 11217 -19213
rect 11137 -19343 11147 -19283
rect 11207 -19343 11217 -19283
rect 11593 -19213 11603 -19163
rect 12061 -19153 12121 -18851
rect 11663 -19213 11673 -19163
rect 11593 -19283 11673 -19213
rect 11593 -19343 11603 -19283
rect 11663 -19343 11673 -19283
rect 12051 -19213 12061 -19163
rect 12517 -19153 12577 -18851
rect 12121 -19213 12131 -19163
rect 12051 -19283 12131 -19213
rect 12051 -19343 12061 -19283
rect 12121 -19343 12131 -19283
rect 12507 -19213 12517 -19163
rect 12973 -19153 13033 -18851
rect 12577 -19213 12587 -19163
rect 12507 -19283 12587 -19213
rect 12507 -19343 12517 -19283
rect 12577 -19343 12587 -19283
rect 12963 -19213 12973 -19163
rect 13431 -19153 13491 -18851
rect 13033 -19213 13043 -19163
rect 12963 -19283 13043 -19213
rect 12963 -19343 12973 -19283
rect 13033 -19343 13043 -19283
rect 13421 -19213 13431 -19163
rect 13887 -19153 13947 -18851
rect 13491 -19213 13501 -19163
rect 13421 -19283 13501 -19213
rect 13421 -19343 13431 -19283
rect 13491 -19343 13501 -19283
rect 13877 -19213 13887 -19163
rect 14343 -19153 14403 -18851
rect 13947 -19213 13957 -19163
rect 13877 -19283 13957 -19213
rect 13877 -19343 13887 -19283
rect 13947 -19343 13957 -19283
rect 14333 -19213 14343 -19163
rect 14801 -19153 14861 -18851
rect 14403 -19213 14413 -19163
rect 14333 -19283 14413 -19213
rect 14333 -19343 14343 -19283
rect 14403 -19343 14413 -19283
rect 14791 -19213 14801 -19163
rect 15257 -19153 15317 -18851
rect 14861 -19213 14871 -19163
rect 14791 -19283 14871 -19213
rect 14791 -19343 14801 -19283
rect 14861 -19343 14871 -19283
rect 15247 -19213 15257 -19163
rect 15317 -19213 15327 -19163
rect 15247 -19283 15327 -19213
rect 15247 -19343 15257 -19283
rect 15317 -19343 15327 -19283
rect 171 -19647 231 -19343
rect 161 -19707 171 -19657
rect 627 -19647 687 -19343
rect 231 -19707 241 -19657
rect 161 -19777 241 -19707
rect 161 -19837 171 -19777
rect 231 -19837 241 -19777
rect 617 -19707 627 -19657
rect 1083 -19647 1143 -19343
rect 687 -19707 697 -19657
rect 617 -19777 697 -19707
rect 617 -19837 627 -19777
rect 687 -19837 697 -19777
rect 1073 -19707 1083 -19657
rect 1541 -19647 1601 -19343
rect 1143 -19707 1153 -19657
rect 1073 -19777 1153 -19707
rect 1073 -19837 1083 -19777
rect 1143 -19837 1153 -19777
rect 1531 -19707 1541 -19657
rect 1997 -19647 2057 -19343
rect 1601 -19707 1611 -19657
rect 1531 -19777 1611 -19707
rect 1531 -19837 1541 -19777
rect 1601 -19837 1611 -19777
rect 1987 -19707 1997 -19657
rect 2453 -19647 2513 -19343
rect 2057 -19707 2067 -19657
rect 1987 -19777 2067 -19707
rect 1987 -19837 1997 -19777
rect 2057 -19837 2067 -19777
rect 2443 -19707 2453 -19657
rect 2911 -19647 2971 -19343
rect 2513 -19707 2523 -19657
rect 2443 -19777 2523 -19707
rect 2443 -19837 2453 -19777
rect 2513 -19837 2523 -19777
rect 2901 -19707 2911 -19657
rect 3367 -19647 3427 -19343
rect 2971 -19707 2981 -19657
rect 2901 -19777 2981 -19707
rect 2901 -19837 2911 -19777
rect 2971 -19837 2981 -19777
rect 3357 -19707 3367 -19657
rect 3823 -19647 3883 -19343
rect 3427 -19707 3437 -19657
rect 3357 -19777 3437 -19707
rect 3357 -19837 3367 -19777
rect 3427 -19837 3437 -19777
rect 3813 -19707 3823 -19657
rect 4281 -19647 4341 -19343
rect 3883 -19707 3893 -19657
rect 3813 -19777 3893 -19707
rect 3813 -19837 3823 -19777
rect 3883 -19837 3893 -19777
rect 4271 -19707 4281 -19657
rect 4737 -19647 4797 -19343
rect 4341 -19707 4351 -19657
rect 4271 -19777 4351 -19707
rect 4271 -19837 4281 -19777
rect 4341 -19837 4351 -19777
rect 4727 -19707 4737 -19657
rect 5193 -19647 5253 -19343
rect 4797 -19707 4807 -19657
rect 4727 -19777 4807 -19707
rect 4727 -19837 4737 -19777
rect 4797 -19837 4807 -19777
rect 5183 -19707 5193 -19657
rect 5651 -19647 5711 -19343
rect 5253 -19707 5263 -19657
rect 5183 -19777 5263 -19707
rect 5183 -19837 5193 -19777
rect 5253 -19837 5263 -19777
rect 5641 -19707 5651 -19657
rect 6107 -19647 6167 -19343
rect 5711 -19707 5721 -19657
rect 5641 -19777 5721 -19707
rect 5641 -19837 5651 -19777
rect 5711 -19837 5721 -19777
rect 6097 -19707 6107 -19657
rect 6563 -19647 6623 -19343
rect 6167 -19707 6177 -19657
rect 6097 -19777 6177 -19707
rect 6097 -19837 6107 -19777
rect 6167 -19837 6177 -19777
rect 6553 -19707 6563 -19657
rect 7021 -19647 7081 -19343
rect 6623 -19707 6633 -19657
rect 6553 -19777 6633 -19707
rect 6553 -19837 6563 -19777
rect 6623 -19837 6633 -19777
rect 7011 -19707 7021 -19657
rect 7477 -19647 7537 -19343
rect 7081 -19707 7091 -19657
rect 7011 -19777 7091 -19707
rect 7011 -19837 7021 -19777
rect 7081 -19837 7091 -19777
rect 7467 -19707 7477 -19657
rect 7933 -19647 7993 -19343
rect 7537 -19707 7547 -19657
rect 7467 -19777 7547 -19707
rect 7467 -19837 7477 -19777
rect 7537 -19837 7547 -19777
rect 7923 -19707 7933 -19657
rect 8407 -19647 8467 -19343
rect 7993 -19707 8003 -19657
rect 7923 -19777 8003 -19707
rect 7923 -19837 7933 -19777
rect 7993 -19837 8003 -19777
rect 8397 -19707 8407 -19657
rect 8863 -19647 8923 -19343
rect 8467 -19707 8477 -19657
rect 8397 -19777 8477 -19707
rect 8397 -19837 8407 -19777
rect 8467 -19837 8477 -19777
rect 8853 -19707 8863 -19657
rect 9321 -19647 9381 -19343
rect 8923 -19707 8933 -19657
rect 8853 -19777 8933 -19707
rect 8853 -19837 8863 -19777
rect 8923 -19837 8933 -19777
rect 9311 -19707 9321 -19657
rect 9777 -19647 9837 -19343
rect 9381 -19707 9391 -19657
rect 9311 -19777 9391 -19707
rect 9311 -19837 9321 -19777
rect 9381 -19837 9391 -19777
rect 9767 -19707 9777 -19657
rect 10233 -19647 10293 -19343
rect 9837 -19707 9847 -19657
rect 9767 -19777 9847 -19707
rect 9767 -19837 9777 -19777
rect 9837 -19837 9847 -19777
rect 10223 -19707 10233 -19657
rect 10691 -19647 10751 -19343
rect 10293 -19707 10303 -19657
rect 10223 -19777 10303 -19707
rect 10223 -19837 10233 -19777
rect 10293 -19837 10303 -19777
rect 10681 -19707 10691 -19657
rect 11147 -19647 11207 -19343
rect 10751 -19707 10761 -19657
rect 10681 -19777 10761 -19707
rect 10681 -19837 10691 -19777
rect 10751 -19837 10761 -19777
rect 11137 -19707 11147 -19657
rect 11603 -19647 11663 -19343
rect 11207 -19707 11217 -19657
rect 11137 -19777 11217 -19707
rect 11137 -19837 11147 -19777
rect 11207 -19837 11217 -19777
rect 11593 -19707 11603 -19657
rect 12061 -19647 12121 -19343
rect 11663 -19707 11673 -19657
rect 11593 -19777 11673 -19707
rect 11593 -19837 11603 -19777
rect 11663 -19837 11673 -19777
rect 12051 -19707 12061 -19657
rect 12517 -19647 12577 -19343
rect 12121 -19707 12131 -19657
rect 12051 -19777 12131 -19707
rect 12051 -19837 12061 -19777
rect 12121 -19837 12131 -19777
rect 12507 -19707 12517 -19657
rect 12973 -19647 13033 -19343
rect 12577 -19707 12587 -19657
rect 12507 -19777 12587 -19707
rect 12507 -19837 12517 -19777
rect 12577 -19837 12587 -19777
rect 12963 -19707 12973 -19657
rect 13431 -19647 13491 -19343
rect 13033 -19707 13043 -19657
rect 12963 -19777 13043 -19707
rect 12963 -19837 12973 -19777
rect 13033 -19837 13043 -19777
rect 13421 -19707 13431 -19657
rect 13887 -19647 13947 -19343
rect 13491 -19707 13501 -19657
rect 13421 -19777 13501 -19707
rect 13421 -19837 13431 -19777
rect 13491 -19837 13501 -19777
rect 13877 -19707 13887 -19657
rect 14343 -19647 14403 -19343
rect 13947 -19707 13957 -19657
rect 13877 -19777 13957 -19707
rect 13877 -19837 13887 -19777
rect 13947 -19837 13957 -19777
rect 14333 -19707 14343 -19657
rect 14801 -19647 14861 -19343
rect 14403 -19707 14413 -19657
rect 14333 -19777 14413 -19707
rect 14333 -19837 14343 -19777
rect 14403 -19837 14413 -19777
rect 14791 -19707 14801 -19657
rect 15257 -19647 15317 -19343
rect 14861 -19707 14871 -19657
rect 14791 -19777 14871 -19707
rect 14791 -19837 14801 -19777
rect 14861 -19837 14871 -19777
rect 15247 -19707 15257 -19657
rect 15317 -19707 15327 -19657
rect 15247 -19777 15327 -19707
rect 15247 -19837 15257 -19777
rect 15317 -19837 15327 -19777
rect 171 -20149 231 -19837
rect 161 -20209 171 -20159
rect 627 -20149 687 -19837
rect 231 -20209 241 -20159
rect 161 -20279 241 -20209
rect 161 -20339 171 -20279
rect 231 -20339 241 -20279
rect 617 -20209 627 -20159
rect 1083 -20149 1143 -19837
rect 687 -20209 697 -20159
rect 617 -20279 697 -20209
rect 617 -20339 627 -20279
rect 687 -20339 697 -20279
rect 1073 -20209 1083 -20159
rect 1541 -20149 1601 -19837
rect 1143 -20209 1153 -20159
rect 1073 -20279 1153 -20209
rect 1073 -20339 1083 -20279
rect 1143 -20339 1153 -20279
rect 1531 -20209 1541 -20159
rect 1997 -20149 2057 -19837
rect 1601 -20209 1611 -20159
rect 1531 -20279 1611 -20209
rect 1531 -20339 1541 -20279
rect 1601 -20339 1611 -20279
rect 1987 -20209 1997 -20159
rect 2453 -20149 2513 -19837
rect 2057 -20209 2067 -20159
rect 1987 -20279 2067 -20209
rect 1987 -20339 1997 -20279
rect 2057 -20339 2067 -20279
rect 2443 -20209 2453 -20159
rect 2911 -20149 2971 -19837
rect 2513 -20209 2523 -20159
rect 2443 -20279 2523 -20209
rect 2443 -20339 2453 -20279
rect 2513 -20339 2523 -20279
rect 2901 -20209 2911 -20159
rect 3367 -20149 3427 -19837
rect 2971 -20209 2981 -20159
rect 2901 -20279 2981 -20209
rect 2901 -20339 2911 -20279
rect 2971 -20339 2981 -20279
rect 3357 -20209 3367 -20159
rect 3823 -20149 3883 -19837
rect 3427 -20209 3437 -20159
rect 3357 -20279 3437 -20209
rect 3357 -20339 3367 -20279
rect 3427 -20339 3437 -20279
rect 3813 -20209 3823 -20159
rect 4281 -20149 4341 -19837
rect 3883 -20209 3893 -20159
rect 3813 -20279 3893 -20209
rect 3813 -20339 3823 -20279
rect 3883 -20339 3893 -20279
rect 4271 -20209 4281 -20159
rect 4737 -20149 4797 -19837
rect 4341 -20209 4351 -20159
rect 4271 -20279 4351 -20209
rect 4271 -20339 4281 -20279
rect 4341 -20339 4351 -20279
rect 4727 -20209 4737 -20159
rect 5193 -20149 5253 -19837
rect 4797 -20209 4807 -20159
rect 4727 -20279 4807 -20209
rect 4727 -20339 4737 -20279
rect 4797 -20339 4807 -20279
rect 5183 -20209 5193 -20159
rect 5651 -20149 5711 -19837
rect 5253 -20209 5263 -20159
rect 5183 -20279 5263 -20209
rect 5183 -20339 5193 -20279
rect 5253 -20339 5263 -20279
rect 5641 -20209 5651 -20159
rect 6107 -20149 6167 -19837
rect 5711 -20209 5721 -20159
rect 5641 -20279 5721 -20209
rect 5641 -20339 5651 -20279
rect 5711 -20339 5721 -20279
rect 6097 -20209 6107 -20159
rect 6563 -20149 6623 -19837
rect 6167 -20209 6177 -20159
rect 6097 -20279 6177 -20209
rect 6097 -20339 6107 -20279
rect 6167 -20339 6177 -20279
rect 6553 -20209 6563 -20159
rect 7021 -20149 7081 -19837
rect 6623 -20209 6633 -20159
rect 6553 -20279 6633 -20209
rect 6553 -20339 6563 -20279
rect 6623 -20339 6633 -20279
rect 7011 -20209 7021 -20159
rect 7477 -20149 7537 -19837
rect 7081 -20209 7091 -20159
rect 7011 -20279 7091 -20209
rect 7011 -20339 7021 -20279
rect 7081 -20339 7091 -20279
rect 7467 -20209 7477 -20159
rect 7933 -20149 7993 -19837
rect 7537 -20209 7547 -20159
rect 7467 -20279 7547 -20209
rect 7467 -20339 7477 -20279
rect 7537 -20339 7547 -20279
rect 7923 -20209 7933 -20159
rect 8407 -20149 8467 -19837
rect 7993 -20209 8003 -20159
rect 7923 -20279 8003 -20209
rect 7923 -20339 7933 -20279
rect 7993 -20339 8003 -20279
rect 8397 -20209 8407 -20159
rect 8863 -20149 8923 -19837
rect 8467 -20209 8477 -20159
rect 8397 -20279 8477 -20209
rect 8397 -20339 8407 -20279
rect 8467 -20339 8477 -20279
rect 8853 -20209 8863 -20159
rect 9321 -20149 9381 -19837
rect 8923 -20209 8933 -20159
rect 8853 -20279 8933 -20209
rect 8853 -20339 8863 -20279
rect 8923 -20339 8933 -20279
rect 9311 -20209 9321 -20159
rect 9777 -20149 9837 -19837
rect 9381 -20209 9391 -20159
rect 9311 -20279 9391 -20209
rect 9311 -20339 9321 -20279
rect 9381 -20339 9391 -20279
rect 9767 -20209 9777 -20159
rect 10233 -20149 10293 -19837
rect 9837 -20209 9847 -20159
rect 9767 -20279 9847 -20209
rect 9767 -20339 9777 -20279
rect 9837 -20339 9847 -20279
rect 10223 -20209 10233 -20159
rect 10691 -20149 10751 -19837
rect 10293 -20209 10303 -20159
rect 10223 -20279 10303 -20209
rect 10223 -20339 10233 -20279
rect 10293 -20339 10303 -20279
rect 10681 -20209 10691 -20159
rect 11147 -20149 11207 -19837
rect 10751 -20209 10761 -20159
rect 10681 -20279 10761 -20209
rect 10681 -20339 10691 -20279
rect 10751 -20339 10761 -20279
rect 11137 -20209 11147 -20159
rect 11603 -20149 11663 -19837
rect 11207 -20209 11217 -20159
rect 11137 -20279 11217 -20209
rect 11137 -20339 11147 -20279
rect 11207 -20339 11217 -20279
rect 11593 -20209 11603 -20159
rect 12061 -20149 12121 -19837
rect 11663 -20209 11673 -20159
rect 11593 -20279 11673 -20209
rect 11593 -20339 11603 -20279
rect 11663 -20339 11673 -20279
rect 12051 -20209 12061 -20159
rect 12517 -20149 12577 -19837
rect 12121 -20209 12131 -20159
rect 12051 -20279 12131 -20209
rect 12051 -20339 12061 -20279
rect 12121 -20339 12131 -20279
rect 12507 -20209 12517 -20159
rect 12973 -20149 13033 -19837
rect 12577 -20209 12587 -20159
rect 12507 -20279 12587 -20209
rect 12507 -20339 12517 -20279
rect 12577 -20339 12587 -20279
rect 12963 -20209 12973 -20159
rect 13431 -20149 13491 -19837
rect 13033 -20209 13043 -20159
rect 12963 -20279 13043 -20209
rect 12963 -20339 12973 -20279
rect 13033 -20339 13043 -20279
rect 13421 -20209 13431 -20159
rect 13887 -20149 13947 -19837
rect 13491 -20209 13501 -20159
rect 13421 -20279 13501 -20209
rect 13421 -20339 13431 -20279
rect 13491 -20339 13501 -20279
rect 13877 -20209 13887 -20159
rect 14343 -20149 14403 -19837
rect 13947 -20209 13957 -20159
rect 13877 -20279 13957 -20209
rect 13877 -20339 13887 -20279
rect 13947 -20339 13957 -20279
rect 14333 -20209 14343 -20159
rect 14801 -20149 14861 -19837
rect 14403 -20209 14413 -20159
rect 14333 -20279 14413 -20209
rect 14333 -20339 14343 -20279
rect 14403 -20339 14413 -20279
rect 14791 -20209 14801 -20159
rect 15257 -20149 15317 -19837
rect 14861 -20209 14871 -20159
rect 14791 -20279 14871 -20209
rect 14791 -20339 14801 -20279
rect 14861 -20339 14871 -20279
rect 15247 -20209 15257 -20159
rect 15317 -20209 15327 -20159
rect 15247 -20279 15327 -20209
rect 15247 -20339 15257 -20279
rect 15317 -20339 15327 -20279
rect 171 -20641 231 -20339
rect 161 -20701 171 -20651
rect 627 -20641 687 -20339
rect 231 -20701 241 -20651
rect 161 -20771 241 -20701
rect 161 -20831 171 -20771
rect 231 -20831 241 -20771
rect 617 -20701 627 -20651
rect 1083 -20641 1143 -20339
rect 687 -20701 697 -20651
rect 617 -20771 697 -20701
rect 617 -20831 627 -20771
rect 687 -20831 697 -20771
rect 1073 -20701 1083 -20651
rect 1541 -20641 1601 -20339
rect 1143 -20701 1153 -20651
rect 1073 -20771 1153 -20701
rect 1073 -20831 1083 -20771
rect 1143 -20831 1153 -20771
rect 1531 -20701 1541 -20651
rect 1997 -20641 2057 -20339
rect 1601 -20701 1611 -20651
rect 1531 -20771 1611 -20701
rect 1531 -20831 1541 -20771
rect 1601 -20831 1611 -20771
rect 1987 -20701 1997 -20651
rect 2453 -20641 2513 -20339
rect 2057 -20701 2067 -20651
rect 1987 -20771 2067 -20701
rect 1987 -20831 1997 -20771
rect 2057 -20831 2067 -20771
rect 2443 -20701 2453 -20651
rect 2911 -20641 2971 -20339
rect 2513 -20701 2523 -20651
rect 2443 -20771 2523 -20701
rect 2443 -20831 2453 -20771
rect 2513 -20831 2523 -20771
rect 2901 -20701 2911 -20651
rect 3367 -20641 3427 -20339
rect 2971 -20701 2981 -20651
rect 2901 -20771 2981 -20701
rect 2901 -20831 2911 -20771
rect 2971 -20831 2981 -20771
rect 3357 -20701 3367 -20651
rect 3823 -20641 3883 -20339
rect 3427 -20701 3437 -20651
rect 3357 -20771 3437 -20701
rect 3357 -20831 3367 -20771
rect 3427 -20831 3437 -20771
rect 3813 -20701 3823 -20651
rect 4281 -20641 4341 -20339
rect 3883 -20701 3893 -20651
rect 3813 -20771 3893 -20701
rect 3813 -20831 3823 -20771
rect 3883 -20831 3893 -20771
rect 4271 -20701 4281 -20651
rect 4737 -20641 4797 -20339
rect 4341 -20701 4351 -20651
rect 4271 -20771 4351 -20701
rect 4271 -20831 4281 -20771
rect 4341 -20831 4351 -20771
rect 4727 -20701 4737 -20651
rect 5193 -20641 5253 -20339
rect 4797 -20701 4807 -20651
rect 4727 -20771 4807 -20701
rect 4727 -20831 4737 -20771
rect 4797 -20831 4807 -20771
rect 5183 -20701 5193 -20651
rect 5651 -20641 5711 -20339
rect 5253 -20701 5263 -20651
rect 5183 -20771 5263 -20701
rect 5183 -20831 5193 -20771
rect 5253 -20831 5263 -20771
rect 5641 -20701 5651 -20651
rect 6107 -20641 6167 -20339
rect 5711 -20701 5721 -20651
rect 5641 -20771 5721 -20701
rect 5641 -20831 5651 -20771
rect 5711 -20831 5721 -20771
rect 6097 -20701 6107 -20651
rect 6563 -20641 6623 -20339
rect 6167 -20701 6177 -20651
rect 6097 -20771 6177 -20701
rect 6097 -20831 6107 -20771
rect 6167 -20831 6177 -20771
rect 6553 -20701 6563 -20651
rect 7021 -20641 7081 -20339
rect 6623 -20701 6633 -20651
rect 6553 -20771 6633 -20701
rect 6553 -20831 6563 -20771
rect 6623 -20831 6633 -20771
rect 7011 -20701 7021 -20651
rect 7477 -20641 7537 -20339
rect 7081 -20701 7091 -20651
rect 7011 -20771 7091 -20701
rect 7011 -20831 7021 -20771
rect 7081 -20831 7091 -20771
rect 7467 -20701 7477 -20651
rect 7933 -20641 7993 -20339
rect 7537 -20701 7547 -20651
rect 7467 -20771 7547 -20701
rect 7467 -20831 7477 -20771
rect 7537 -20831 7547 -20771
rect 7923 -20701 7933 -20651
rect 8407 -20641 8467 -20339
rect 7993 -20701 8003 -20651
rect 7923 -20771 8003 -20701
rect 7923 -20831 7933 -20771
rect 7993 -20831 8003 -20771
rect 8397 -20701 8407 -20651
rect 8863 -20641 8923 -20339
rect 8467 -20701 8477 -20651
rect 8397 -20771 8477 -20701
rect 8397 -20831 8407 -20771
rect 8467 -20831 8477 -20771
rect 8853 -20701 8863 -20651
rect 9321 -20641 9381 -20339
rect 8923 -20701 8933 -20651
rect 8853 -20771 8933 -20701
rect 8853 -20831 8863 -20771
rect 8923 -20831 8933 -20771
rect 9311 -20701 9321 -20651
rect 9777 -20641 9837 -20339
rect 9381 -20701 9391 -20651
rect 9311 -20771 9391 -20701
rect 9311 -20831 9321 -20771
rect 9381 -20831 9391 -20771
rect 9767 -20701 9777 -20651
rect 10233 -20641 10293 -20339
rect 9837 -20701 9847 -20651
rect 9767 -20771 9847 -20701
rect 9767 -20831 9777 -20771
rect 9837 -20831 9847 -20771
rect 10223 -20701 10233 -20651
rect 10691 -20641 10751 -20339
rect 10293 -20701 10303 -20651
rect 10223 -20771 10303 -20701
rect 10223 -20831 10233 -20771
rect 10293 -20831 10303 -20771
rect 10681 -20701 10691 -20651
rect 11147 -20641 11207 -20339
rect 10751 -20701 10761 -20651
rect 10681 -20771 10761 -20701
rect 10681 -20831 10691 -20771
rect 10751 -20831 10761 -20771
rect 11137 -20701 11147 -20651
rect 11603 -20641 11663 -20339
rect 11207 -20701 11217 -20651
rect 11137 -20771 11217 -20701
rect 11137 -20831 11147 -20771
rect 11207 -20831 11217 -20771
rect 11593 -20701 11603 -20651
rect 12061 -20641 12121 -20339
rect 11663 -20701 11673 -20651
rect 11593 -20771 11673 -20701
rect 11593 -20831 11603 -20771
rect 11663 -20831 11673 -20771
rect 12051 -20701 12061 -20651
rect 12517 -20641 12577 -20339
rect 12121 -20701 12131 -20651
rect 12051 -20771 12131 -20701
rect 12051 -20831 12061 -20771
rect 12121 -20831 12131 -20771
rect 12507 -20701 12517 -20651
rect 12973 -20641 13033 -20339
rect 12577 -20701 12587 -20651
rect 12507 -20771 12587 -20701
rect 12507 -20831 12517 -20771
rect 12577 -20831 12587 -20771
rect 12963 -20701 12973 -20651
rect 13431 -20641 13491 -20339
rect 13033 -20701 13043 -20651
rect 12963 -20771 13043 -20701
rect 12963 -20831 12973 -20771
rect 13033 -20831 13043 -20771
rect 13421 -20701 13431 -20651
rect 13887 -20641 13947 -20339
rect 13491 -20701 13501 -20651
rect 13421 -20771 13501 -20701
rect 13421 -20831 13431 -20771
rect 13491 -20831 13501 -20771
rect 13877 -20701 13887 -20651
rect 14343 -20641 14403 -20339
rect 13947 -20701 13957 -20651
rect 13877 -20771 13957 -20701
rect 13877 -20831 13887 -20771
rect 13947 -20831 13957 -20771
rect 14333 -20701 14343 -20651
rect 14801 -20641 14861 -20339
rect 14403 -20701 14413 -20651
rect 14333 -20771 14413 -20701
rect 14333 -20831 14343 -20771
rect 14403 -20831 14413 -20771
rect 14791 -20701 14801 -20651
rect 15257 -20641 15317 -20339
rect 14861 -20701 14871 -20651
rect 14791 -20771 14871 -20701
rect 14791 -20831 14801 -20771
rect 14861 -20831 14871 -20771
rect 15247 -20701 15257 -20651
rect 15317 -20701 15327 -20651
rect 15247 -20771 15327 -20701
rect 15247 -20831 15257 -20771
rect 15317 -20831 15327 -20771
rect 171 -21157 231 -20831
rect 161 -21217 171 -21167
rect 627 -21157 687 -20831
rect 231 -21217 241 -21167
rect 161 -21287 241 -21217
rect 161 -21347 171 -21287
rect 231 -21347 241 -21287
rect 617 -21217 627 -21167
rect 1083 -21157 1143 -20831
rect 687 -21217 697 -21167
rect 617 -21287 697 -21217
rect 617 -21347 627 -21287
rect 687 -21347 697 -21287
rect 1073 -21217 1083 -21167
rect 1541 -21157 1601 -20831
rect 1143 -21217 1153 -21167
rect 1073 -21287 1153 -21217
rect 1073 -21347 1083 -21287
rect 1143 -21347 1153 -21287
rect 1531 -21217 1541 -21167
rect 1997 -21157 2057 -20831
rect 1601 -21217 1611 -21167
rect 1531 -21287 1611 -21217
rect 1531 -21347 1541 -21287
rect 1601 -21347 1611 -21287
rect 1987 -21217 1997 -21167
rect 2453 -21157 2513 -20831
rect 2057 -21217 2067 -21167
rect 1987 -21287 2067 -21217
rect 1987 -21347 1997 -21287
rect 2057 -21347 2067 -21287
rect 2443 -21217 2453 -21167
rect 2911 -21157 2971 -20831
rect 2513 -21217 2523 -21167
rect 2443 -21287 2523 -21217
rect 2443 -21347 2453 -21287
rect 2513 -21347 2523 -21287
rect 2901 -21217 2911 -21167
rect 3367 -21157 3427 -20831
rect 2971 -21217 2981 -21167
rect 2901 -21287 2981 -21217
rect 2901 -21347 2911 -21287
rect 2971 -21347 2981 -21287
rect 3357 -21217 3367 -21167
rect 3823 -21157 3883 -20831
rect 3427 -21217 3437 -21167
rect 3357 -21287 3437 -21217
rect 3357 -21347 3367 -21287
rect 3427 -21347 3437 -21287
rect 3813 -21217 3823 -21167
rect 4281 -21157 4341 -20831
rect 3883 -21217 3893 -21167
rect 3813 -21287 3893 -21217
rect 3813 -21347 3823 -21287
rect 3883 -21347 3893 -21287
rect 4271 -21217 4281 -21167
rect 4737 -21157 4797 -20831
rect 4341 -21217 4351 -21167
rect 4271 -21287 4351 -21217
rect 4271 -21347 4281 -21287
rect 4341 -21347 4351 -21287
rect 4727 -21217 4737 -21167
rect 5193 -21157 5253 -20831
rect 4797 -21217 4807 -21167
rect 4727 -21287 4807 -21217
rect 4727 -21347 4737 -21287
rect 4797 -21347 4807 -21287
rect 5183 -21217 5193 -21167
rect 5651 -21157 5711 -20831
rect 5253 -21217 5263 -21167
rect 5183 -21287 5263 -21217
rect 5183 -21347 5193 -21287
rect 5253 -21347 5263 -21287
rect 5641 -21217 5651 -21167
rect 6107 -21157 6167 -20831
rect 5711 -21217 5721 -21167
rect 5641 -21287 5721 -21217
rect 5641 -21347 5651 -21287
rect 5711 -21347 5721 -21287
rect 6097 -21217 6107 -21167
rect 6563 -21157 6623 -20831
rect 6167 -21217 6177 -21167
rect 6097 -21287 6177 -21217
rect 6097 -21347 6107 -21287
rect 6167 -21347 6177 -21287
rect 6553 -21217 6563 -21167
rect 7021 -21157 7081 -20831
rect 6623 -21217 6633 -21167
rect 6553 -21287 6633 -21217
rect 6553 -21347 6563 -21287
rect 6623 -21347 6633 -21287
rect 7011 -21217 7021 -21167
rect 7477 -21157 7537 -20831
rect 7081 -21217 7091 -21167
rect 7011 -21287 7091 -21217
rect 7011 -21347 7021 -21287
rect 7081 -21347 7091 -21287
rect 7467 -21217 7477 -21167
rect 7933 -21157 7993 -20831
rect 7537 -21217 7547 -21167
rect 7467 -21287 7547 -21217
rect 7467 -21347 7477 -21287
rect 7537 -21347 7547 -21287
rect 7923 -21217 7933 -21167
rect 8407 -21157 8467 -20831
rect 7993 -21217 8003 -21167
rect 7923 -21287 8003 -21217
rect 7923 -21347 7933 -21287
rect 7993 -21347 8003 -21287
rect 8397 -21217 8407 -21167
rect 8863 -21157 8923 -20831
rect 8467 -21217 8477 -21167
rect 8397 -21287 8477 -21217
rect 8397 -21347 8407 -21287
rect 8467 -21347 8477 -21287
rect 8853 -21217 8863 -21167
rect 9321 -21157 9381 -20831
rect 8923 -21217 8933 -21167
rect 8853 -21287 8933 -21217
rect 8853 -21347 8863 -21287
rect 8923 -21347 8933 -21287
rect 9311 -21217 9321 -21167
rect 9777 -21157 9837 -20831
rect 9381 -21217 9391 -21167
rect 9311 -21287 9391 -21217
rect 9311 -21347 9321 -21287
rect 9381 -21347 9391 -21287
rect 9767 -21217 9777 -21167
rect 10233 -21157 10293 -20831
rect 9837 -21217 9847 -21167
rect 9767 -21287 9847 -21217
rect 9767 -21347 9777 -21287
rect 9837 -21347 9847 -21287
rect 10223 -21217 10233 -21167
rect 10691 -21157 10751 -20831
rect 10293 -21217 10303 -21167
rect 10223 -21287 10303 -21217
rect 10223 -21347 10233 -21287
rect 10293 -21347 10303 -21287
rect 10681 -21217 10691 -21167
rect 11147 -21157 11207 -20831
rect 10751 -21217 10761 -21167
rect 10681 -21287 10761 -21217
rect 10681 -21347 10691 -21287
rect 10751 -21347 10761 -21287
rect 11137 -21217 11147 -21167
rect 11603 -21157 11663 -20831
rect 11207 -21217 11217 -21167
rect 11137 -21287 11217 -21217
rect 11137 -21347 11147 -21287
rect 11207 -21347 11217 -21287
rect 11593 -21217 11603 -21167
rect 12061 -21157 12121 -20831
rect 11663 -21217 11673 -21167
rect 11593 -21287 11673 -21217
rect 11593 -21347 11603 -21287
rect 11663 -21347 11673 -21287
rect 12051 -21217 12061 -21167
rect 12517 -21157 12577 -20831
rect 12121 -21217 12131 -21167
rect 12051 -21287 12131 -21217
rect 12051 -21347 12061 -21287
rect 12121 -21347 12131 -21287
rect 12507 -21217 12517 -21167
rect 12973 -21157 13033 -20831
rect 12577 -21217 12587 -21167
rect 12507 -21287 12587 -21217
rect 12507 -21347 12517 -21287
rect 12577 -21347 12587 -21287
rect 12963 -21217 12973 -21167
rect 13431 -21157 13491 -20831
rect 13033 -21217 13043 -21167
rect 12963 -21287 13043 -21217
rect 12963 -21347 12973 -21287
rect 13033 -21347 13043 -21287
rect 13421 -21217 13431 -21167
rect 13887 -21157 13947 -20831
rect 13491 -21217 13501 -21167
rect 13421 -21287 13501 -21217
rect 13421 -21347 13431 -21287
rect 13491 -21347 13501 -21287
rect 13877 -21217 13887 -21167
rect 14343 -21157 14403 -20831
rect 13947 -21217 13957 -21167
rect 13877 -21287 13957 -21217
rect 13877 -21347 13887 -21287
rect 13947 -21347 13957 -21287
rect 14333 -21217 14343 -21167
rect 14801 -21157 14861 -20831
rect 14403 -21217 14413 -21167
rect 14333 -21287 14413 -21217
rect 14333 -21347 14343 -21287
rect 14403 -21347 14413 -21287
rect 14791 -21217 14801 -21167
rect 15257 -21157 15317 -20831
rect 14861 -21217 14871 -21167
rect 14791 -21287 14871 -21217
rect 14791 -21347 14801 -21287
rect 14861 -21347 14871 -21287
rect 15247 -21217 15257 -21167
rect 15317 -21217 15327 -21167
rect 15247 -21287 15327 -21217
rect 15247 -21347 15257 -21287
rect 15317 -21347 15327 -21287
rect 171 -21659 231 -21347
rect 161 -21719 171 -21669
rect 627 -21659 687 -21347
rect 231 -21719 241 -21669
rect 161 -21789 241 -21719
rect 161 -21849 171 -21789
rect 231 -21849 241 -21789
rect 617 -21719 627 -21669
rect 1083 -21659 1143 -21347
rect 687 -21719 697 -21669
rect 617 -21789 697 -21719
rect 617 -21849 627 -21789
rect 687 -21849 697 -21789
rect 1073 -21719 1083 -21669
rect 1541 -21659 1601 -21347
rect 1143 -21719 1153 -21669
rect 1073 -21789 1153 -21719
rect 1073 -21849 1083 -21789
rect 1143 -21849 1153 -21789
rect 1531 -21719 1541 -21669
rect 1997 -21659 2057 -21347
rect 1601 -21719 1611 -21669
rect 1531 -21789 1611 -21719
rect 1531 -21849 1541 -21789
rect 1601 -21849 1611 -21789
rect 1987 -21719 1997 -21669
rect 2453 -21659 2513 -21347
rect 2057 -21719 2067 -21669
rect 1987 -21789 2067 -21719
rect 1987 -21849 1997 -21789
rect 2057 -21849 2067 -21789
rect 2443 -21719 2453 -21669
rect 2911 -21659 2971 -21347
rect 2513 -21719 2523 -21669
rect 2443 -21789 2523 -21719
rect 2443 -21849 2453 -21789
rect 2513 -21849 2523 -21789
rect 2901 -21719 2911 -21669
rect 3367 -21659 3427 -21347
rect 2971 -21719 2981 -21669
rect 2901 -21789 2981 -21719
rect 2901 -21849 2911 -21789
rect 2971 -21849 2981 -21789
rect 3357 -21719 3367 -21669
rect 3823 -21659 3883 -21347
rect 3427 -21719 3437 -21669
rect 3357 -21789 3437 -21719
rect 3357 -21849 3367 -21789
rect 3427 -21849 3437 -21789
rect 3813 -21719 3823 -21669
rect 4281 -21659 4341 -21347
rect 3883 -21719 3893 -21669
rect 3813 -21789 3893 -21719
rect 3813 -21849 3823 -21789
rect 3883 -21849 3893 -21789
rect 4271 -21719 4281 -21669
rect 4737 -21659 4797 -21347
rect 4341 -21719 4351 -21669
rect 4271 -21789 4351 -21719
rect 4271 -21849 4281 -21789
rect 4341 -21849 4351 -21789
rect 4727 -21719 4737 -21669
rect 5193 -21659 5253 -21347
rect 4797 -21719 4807 -21669
rect 4727 -21789 4807 -21719
rect 4727 -21849 4737 -21789
rect 4797 -21849 4807 -21789
rect 5183 -21719 5193 -21669
rect 5651 -21659 5711 -21347
rect 5253 -21719 5263 -21669
rect 5183 -21789 5263 -21719
rect 5183 -21849 5193 -21789
rect 5253 -21849 5263 -21789
rect 5641 -21719 5651 -21669
rect 6107 -21659 6167 -21347
rect 5711 -21719 5721 -21669
rect 5641 -21789 5721 -21719
rect 5641 -21849 5651 -21789
rect 5711 -21849 5721 -21789
rect 6097 -21719 6107 -21669
rect 6563 -21659 6623 -21347
rect 6167 -21719 6177 -21669
rect 6097 -21789 6177 -21719
rect 6097 -21849 6107 -21789
rect 6167 -21849 6177 -21789
rect 6553 -21719 6563 -21669
rect 7021 -21659 7081 -21347
rect 6623 -21719 6633 -21669
rect 6553 -21789 6633 -21719
rect 6553 -21849 6563 -21789
rect 6623 -21849 6633 -21789
rect 7011 -21719 7021 -21669
rect 7477 -21659 7537 -21347
rect 7081 -21719 7091 -21669
rect 7011 -21789 7091 -21719
rect 7011 -21849 7021 -21789
rect 7081 -21849 7091 -21789
rect 7467 -21719 7477 -21669
rect 7933 -21659 7993 -21347
rect 7537 -21719 7547 -21669
rect 7467 -21789 7547 -21719
rect 7467 -21849 7477 -21789
rect 7537 -21849 7547 -21789
rect 7923 -21719 7933 -21669
rect 8407 -21659 8467 -21347
rect 7993 -21719 8003 -21669
rect 7923 -21789 8003 -21719
rect 7923 -21849 7933 -21789
rect 7993 -21849 8003 -21789
rect 8397 -21719 8407 -21669
rect 8863 -21659 8923 -21347
rect 8467 -21719 8477 -21669
rect 8397 -21789 8477 -21719
rect 8397 -21849 8407 -21789
rect 8467 -21849 8477 -21789
rect 8853 -21719 8863 -21669
rect 9321 -21659 9381 -21347
rect 8923 -21719 8933 -21669
rect 8853 -21789 8933 -21719
rect 8853 -21849 8863 -21789
rect 8923 -21849 8933 -21789
rect 9311 -21719 9321 -21669
rect 9777 -21659 9837 -21347
rect 9381 -21719 9391 -21669
rect 9311 -21789 9391 -21719
rect 9311 -21849 9321 -21789
rect 9381 -21849 9391 -21789
rect 9767 -21719 9777 -21669
rect 10233 -21659 10293 -21347
rect 9837 -21719 9847 -21669
rect 9767 -21789 9847 -21719
rect 9767 -21849 9777 -21789
rect 9837 -21849 9847 -21789
rect 10223 -21719 10233 -21669
rect 10691 -21659 10751 -21347
rect 10293 -21719 10303 -21669
rect 10223 -21789 10303 -21719
rect 10223 -21849 10233 -21789
rect 10293 -21849 10303 -21789
rect 10681 -21719 10691 -21669
rect 11147 -21659 11207 -21347
rect 10751 -21719 10761 -21669
rect 10681 -21789 10761 -21719
rect 10681 -21849 10691 -21789
rect 10751 -21849 10761 -21789
rect 11137 -21719 11147 -21669
rect 11603 -21659 11663 -21347
rect 11207 -21719 11217 -21669
rect 11137 -21789 11217 -21719
rect 11137 -21849 11147 -21789
rect 11207 -21849 11217 -21789
rect 11593 -21719 11603 -21669
rect 12061 -21659 12121 -21347
rect 11663 -21719 11673 -21669
rect 11593 -21789 11673 -21719
rect 11593 -21849 11603 -21789
rect 11663 -21849 11673 -21789
rect 12051 -21719 12061 -21669
rect 12517 -21659 12577 -21347
rect 12121 -21719 12131 -21669
rect 12051 -21789 12131 -21719
rect 12051 -21849 12061 -21789
rect 12121 -21849 12131 -21789
rect 12507 -21719 12517 -21669
rect 12973 -21659 13033 -21347
rect 12577 -21719 12587 -21669
rect 12507 -21789 12587 -21719
rect 12507 -21849 12517 -21789
rect 12577 -21849 12587 -21789
rect 12963 -21719 12973 -21669
rect 13431 -21659 13491 -21347
rect 13033 -21719 13043 -21669
rect 12963 -21789 13043 -21719
rect 12963 -21849 12973 -21789
rect 13033 -21849 13043 -21789
rect 13421 -21719 13431 -21669
rect 13887 -21659 13947 -21347
rect 13491 -21719 13501 -21669
rect 13421 -21789 13501 -21719
rect 13421 -21849 13431 -21789
rect 13491 -21849 13501 -21789
rect 13877 -21719 13887 -21669
rect 14343 -21659 14403 -21347
rect 13947 -21719 13957 -21669
rect 13877 -21789 13957 -21719
rect 13877 -21849 13887 -21789
rect 13947 -21849 13957 -21789
rect 14333 -21719 14343 -21669
rect 14801 -21659 14861 -21347
rect 14403 -21719 14413 -21669
rect 14333 -21789 14413 -21719
rect 14333 -21849 14343 -21789
rect 14403 -21849 14413 -21789
rect 14791 -21719 14801 -21669
rect 15257 -21659 15317 -21347
rect 14861 -21719 14871 -21669
rect 14791 -21789 14871 -21719
rect 14791 -21849 14801 -21789
rect 14861 -21849 14871 -21789
rect 15247 -21719 15257 -21669
rect 15317 -21719 15327 -21669
rect 15247 -21789 15327 -21719
rect 15247 -21849 15257 -21789
rect 15317 -21849 15327 -21789
rect 171 -22151 231 -21849
rect 161 -22211 171 -22161
rect 627 -22151 687 -21849
rect 231 -22211 241 -22161
rect 161 -22281 241 -22211
rect 161 -22341 171 -22281
rect 231 -22341 241 -22281
rect 617 -22211 627 -22161
rect 1083 -22151 1143 -21849
rect 687 -22211 697 -22161
rect 617 -22281 697 -22211
rect 617 -22341 627 -22281
rect 687 -22341 697 -22281
rect 1073 -22211 1083 -22161
rect 1541 -22151 1601 -21849
rect 1143 -22211 1153 -22161
rect 1073 -22281 1153 -22211
rect 1073 -22341 1083 -22281
rect 1143 -22341 1153 -22281
rect 1531 -22211 1541 -22161
rect 1997 -22151 2057 -21849
rect 1601 -22211 1611 -22161
rect 1531 -22281 1611 -22211
rect 1531 -22341 1541 -22281
rect 1601 -22341 1611 -22281
rect 1987 -22211 1997 -22161
rect 2453 -22151 2513 -21849
rect 2057 -22211 2067 -22161
rect 1987 -22281 2067 -22211
rect 1987 -22341 1997 -22281
rect 2057 -22341 2067 -22281
rect 2443 -22211 2453 -22161
rect 2911 -22151 2971 -21849
rect 2513 -22211 2523 -22161
rect 2443 -22281 2523 -22211
rect 2443 -22341 2453 -22281
rect 2513 -22341 2523 -22281
rect 2901 -22211 2911 -22161
rect 3367 -22151 3427 -21849
rect 2971 -22211 2981 -22161
rect 2901 -22281 2981 -22211
rect 2901 -22341 2911 -22281
rect 2971 -22341 2981 -22281
rect 3357 -22211 3367 -22161
rect 3823 -22151 3883 -21849
rect 3427 -22211 3437 -22161
rect 3357 -22281 3437 -22211
rect 3357 -22341 3367 -22281
rect 3427 -22341 3437 -22281
rect 3813 -22211 3823 -22161
rect 4281 -22151 4341 -21849
rect 3883 -22211 3893 -22161
rect 3813 -22281 3893 -22211
rect 3813 -22341 3823 -22281
rect 3883 -22341 3893 -22281
rect 4271 -22211 4281 -22161
rect 4737 -22151 4797 -21849
rect 4341 -22211 4351 -22161
rect 4271 -22281 4351 -22211
rect 4271 -22341 4281 -22281
rect 4341 -22341 4351 -22281
rect 4727 -22211 4737 -22161
rect 5193 -22151 5253 -21849
rect 4797 -22211 4807 -22161
rect 4727 -22281 4807 -22211
rect 4727 -22341 4737 -22281
rect 4797 -22341 4807 -22281
rect 5183 -22211 5193 -22161
rect 5651 -22151 5711 -21849
rect 5253 -22211 5263 -22161
rect 5183 -22281 5263 -22211
rect 5183 -22341 5193 -22281
rect 5253 -22341 5263 -22281
rect 5641 -22211 5651 -22161
rect 6107 -22151 6167 -21849
rect 5711 -22211 5721 -22161
rect 5641 -22281 5721 -22211
rect 5641 -22341 5651 -22281
rect 5711 -22341 5721 -22281
rect 6097 -22211 6107 -22161
rect 6563 -22151 6623 -21849
rect 6167 -22211 6177 -22161
rect 6097 -22281 6177 -22211
rect 6097 -22341 6107 -22281
rect 6167 -22341 6177 -22281
rect 6553 -22211 6563 -22161
rect 7021 -22151 7081 -21849
rect 6623 -22211 6633 -22161
rect 6553 -22281 6633 -22211
rect 6553 -22341 6563 -22281
rect 6623 -22341 6633 -22281
rect 7011 -22211 7021 -22161
rect 7477 -22151 7537 -21849
rect 7081 -22211 7091 -22161
rect 7011 -22281 7091 -22211
rect 7011 -22341 7021 -22281
rect 7081 -22341 7091 -22281
rect 7467 -22211 7477 -22161
rect 7933 -22151 7993 -21849
rect 7537 -22211 7547 -22161
rect 7467 -22281 7547 -22211
rect 7467 -22341 7477 -22281
rect 7537 -22341 7547 -22281
rect 7923 -22211 7933 -22161
rect 8407 -22151 8467 -21849
rect 7993 -22211 8003 -22161
rect 7923 -22281 8003 -22211
rect 7923 -22341 7933 -22281
rect 7993 -22341 8003 -22281
rect 8397 -22211 8407 -22161
rect 8863 -22151 8923 -21849
rect 8467 -22211 8477 -22161
rect 8397 -22281 8477 -22211
rect 8397 -22341 8407 -22281
rect 8467 -22341 8477 -22281
rect 8853 -22211 8863 -22161
rect 9321 -22151 9381 -21849
rect 8923 -22211 8933 -22161
rect 8853 -22281 8933 -22211
rect 8853 -22341 8863 -22281
rect 8923 -22341 8933 -22281
rect 9311 -22211 9321 -22161
rect 9777 -22151 9837 -21849
rect 9381 -22211 9391 -22161
rect 9311 -22281 9391 -22211
rect 9311 -22341 9321 -22281
rect 9381 -22341 9391 -22281
rect 9767 -22211 9777 -22161
rect 10233 -22151 10293 -21849
rect 9837 -22211 9847 -22161
rect 9767 -22281 9847 -22211
rect 9767 -22341 9777 -22281
rect 9837 -22341 9847 -22281
rect 10223 -22211 10233 -22161
rect 10691 -22151 10751 -21849
rect 10293 -22211 10303 -22161
rect 10223 -22281 10303 -22211
rect 10223 -22341 10233 -22281
rect 10293 -22341 10303 -22281
rect 10681 -22211 10691 -22161
rect 11147 -22151 11207 -21849
rect 10751 -22211 10761 -22161
rect 10681 -22281 10761 -22211
rect 10681 -22341 10691 -22281
rect 10751 -22341 10761 -22281
rect 11137 -22211 11147 -22161
rect 11603 -22151 11663 -21849
rect 11207 -22211 11217 -22161
rect 11137 -22281 11217 -22211
rect 11137 -22341 11147 -22281
rect 11207 -22341 11217 -22281
rect 11593 -22211 11603 -22161
rect 12061 -22151 12121 -21849
rect 11663 -22211 11673 -22161
rect 11593 -22281 11673 -22211
rect 11593 -22341 11603 -22281
rect 11663 -22341 11673 -22281
rect 12051 -22211 12061 -22161
rect 12517 -22151 12577 -21849
rect 12121 -22211 12131 -22161
rect 12051 -22281 12131 -22211
rect 12051 -22341 12061 -22281
rect 12121 -22341 12131 -22281
rect 12507 -22211 12517 -22161
rect 12973 -22151 13033 -21849
rect 12577 -22211 12587 -22161
rect 12507 -22281 12587 -22211
rect 12507 -22341 12517 -22281
rect 12577 -22341 12587 -22281
rect 12963 -22211 12973 -22161
rect 13431 -22151 13491 -21849
rect 13033 -22211 13043 -22161
rect 12963 -22281 13043 -22211
rect 12963 -22341 12973 -22281
rect 13033 -22341 13043 -22281
rect 13421 -22211 13431 -22161
rect 13887 -22151 13947 -21849
rect 13491 -22211 13501 -22161
rect 13421 -22281 13501 -22211
rect 13421 -22341 13431 -22281
rect 13491 -22341 13501 -22281
rect 13877 -22211 13887 -22161
rect 14343 -22151 14403 -21849
rect 13947 -22211 13957 -22161
rect 13877 -22281 13957 -22211
rect 13877 -22341 13887 -22281
rect 13947 -22341 13957 -22281
rect 14333 -22211 14343 -22161
rect 14801 -22151 14861 -21849
rect 14403 -22211 14413 -22161
rect 14333 -22281 14413 -22211
rect 14333 -22341 14343 -22281
rect 14403 -22341 14413 -22281
rect 14791 -22211 14801 -22161
rect 15257 -22151 15317 -21849
rect 14861 -22211 14871 -22161
rect 14791 -22281 14871 -22211
rect 14791 -22341 14801 -22281
rect 14861 -22341 14871 -22281
rect 15247 -22211 15257 -22161
rect 15317 -22211 15327 -22161
rect 15247 -22281 15327 -22211
rect 15247 -22341 15257 -22281
rect 15317 -22341 15327 -22281
rect 171 -22638 231 -22341
rect 627 -22638 687 -22341
rect 1083 -22638 1143 -22341
rect 1541 -22638 1601 -22341
rect 1997 -22638 2057 -22341
rect 2453 -22638 2513 -22341
rect 2911 -22638 2971 -22341
rect 3367 -22638 3427 -22341
rect 3823 -22638 3883 -22341
rect 4281 -22638 4341 -22341
rect 4737 -22638 4797 -22341
rect 5193 -22638 5253 -22341
rect 5651 -22638 5711 -22341
rect 6107 -22638 6167 -22341
rect 6563 -22638 6623 -22341
rect 7021 -22638 7081 -22341
rect 7477 -22638 7537 -22341
rect 7933 -22638 7993 -22341
rect 8407 -22638 8467 -22341
rect 8863 -22638 8923 -22341
rect 9321 -22638 9381 -22341
rect 9777 -22638 9837 -22341
rect 10233 -22638 10293 -22341
rect 10691 -22638 10751 -22341
rect 11147 -22638 11207 -22341
rect 11603 -22638 11663 -22341
rect 12061 -22638 12121 -22341
rect 12517 -22638 12577 -22341
rect 12973 -22638 13033 -22341
rect 13431 -22638 13491 -22341
rect 13887 -22638 13947 -22341
rect 14343 -22638 14403 -22341
rect 14801 -22638 14861 -22341
rect 15257 -22638 15317 -22341
rect 161 -22698 171 -22638
rect 231 -22698 241 -22638
rect 161 -22768 241 -22698
rect 161 -22818 171 -22768
rect 231 -22818 241 -22768
rect 617 -22698 627 -22638
rect 687 -22698 697 -22638
rect 617 -22768 697 -22698
rect 617 -22818 627 -22768
rect 171 -23140 231 -22828
rect 687 -22818 697 -22768
rect 1073 -22698 1083 -22638
rect 1143 -22698 1153 -22638
rect 1073 -22768 1153 -22698
rect 1073 -22818 1083 -22768
rect 627 -23140 687 -22828
rect 1143 -22818 1153 -22768
rect 1531 -22698 1541 -22638
rect 1601 -22698 1611 -22638
rect 1531 -22768 1611 -22698
rect 1531 -22818 1541 -22768
rect 1083 -23140 1143 -22828
rect 1601 -22818 1611 -22768
rect 1987 -22698 1997 -22638
rect 2057 -22698 2067 -22638
rect 1987 -22768 2067 -22698
rect 1987 -22818 1997 -22768
rect 1541 -23140 1601 -22828
rect 2057 -22818 2067 -22768
rect 2443 -22698 2453 -22638
rect 2513 -22698 2523 -22638
rect 2443 -22768 2523 -22698
rect 2443 -22818 2453 -22768
rect 1997 -23140 2057 -22828
rect 2513 -22818 2523 -22768
rect 2901 -22698 2911 -22638
rect 2971 -22698 2981 -22638
rect 2901 -22768 2981 -22698
rect 2901 -22818 2911 -22768
rect 2453 -23140 2513 -22828
rect 2971 -22818 2981 -22768
rect 3357 -22698 3367 -22638
rect 3427 -22698 3437 -22638
rect 3357 -22768 3437 -22698
rect 3357 -22818 3367 -22768
rect 2911 -23140 2971 -22828
rect 3427 -22818 3437 -22768
rect 3813 -22698 3823 -22638
rect 3883 -22698 3893 -22638
rect 3813 -22768 3893 -22698
rect 3813 -22818 3823 -22768
rect 3367 -23140 3427 -22828
rect 3883 -22818 3893 -22768
rect 4271 -22698 4281 -22638
rect 4341 -22698 4351 -22638
rect 4271 -22768 4351 -22698
rect 4271 -22818 4281 -22768
rect 3823 -23140 3883 -22828
rect 4341 -22818 4351 -22768
rect 4727 -22698 4737 -22638
rect 4797 -22698 4807 -22638
rect 4727 -22768 4807 -22698
rect 4727 -22818 4737 -22768
rect 4281 -23140 4341 -22828
rect 4797 -22818 4807 -22768
rect 5183 -22698 5193 -22638
rect 5253 -22698 5263 -22638
rect 5183 -22768 5263 -22698
rect 5183 -22818 5193 -22768
rect 4737 -23140 4797 -22828
rect 5253 -22818 5263 -22768
rect 5641 -22698 5651 -22638
rect 5711 -22698 5721 -22638
rect 5641 -22768 5721 -22698
rect 5641 -22818 5651 -22768
rect 5193 -23140 5253 -22828
rect 5711 -22818 5721 -22768
rect 6097 -22698 6107 -22638
rect 6167 -22698 6177 -22638
rect 6097 -22768 6177 -22698
rect 6097 -22818 6107 -22768
rect 5651 -23140 5711 -22828
rect 6167 -22818 6177 -22768
rect 6553 -22698 6563 -22638
rect 6623 -22698 6633 -22638
rect 6553 -22768 6633 -22698
rect 6553 -22818 6563 -22768
rect 6107 -23140 6167 -22828
rect 6623 -22818 6633 -22768
rect 7011 -22698 7021 -22638
rect 7081 -22698 7091 -22638
rect 7011 -22768 7091 -22698
rect 7011 -22818 7021 -22768
rect 6563 -23140 6623 -22828
rect 7081 -22818 7091 -22768
rect 7467 -22698 7477 -22638
rect 7537 -22698 7547 -22638
rect 7467 -22768 7547 -22698
rect 7467 -22818 7477 -22768
rect 7021 -23140 7081 -22828
rect 7537 -22818 7547 -22768
rect 7923 -22698 7933 -22638
rect 7993 -22698 8003 -22638
rect 7923 -22768 8003 -22698
rect 7923 -22818 7933 -22768
rect 7477 -23140 7537 -22828
rect 7993 -22818 8003 -22768
rect 8397 -22698 8407 -22638
rect 8467 -22698 8477 -22638
rect 8397 -22768 8477 -22698
rect 8397 -22818 8407 -22768
rect 7933 -23140 7993 -22828
rect 8467 -22818 8477 -22768
rect 8853 -22698 8863 -22638
rect 8923 -22698 8933 -22638
rect 8853 -22768 8933 -22698
rect 8853 -22818 8863 -22768
rect 8407 -23140 8467 -22828
rect 8923 -22818 8933 -22768
rect 9311 -22698 9321 -22638
rect 9381 -22698 9391 -22638
rect 9311 -22768 9391 -22698
rect 9311 -22818 9321 -22768
rect 8863 -23140 8923 -22828
rect 9381 -22818 9391 -22768
rect 9767 -22698 9777 -22638
rect 9837 -22698 9847 -22638
rect 9767 -22768 9847 -22698
rect 9767 -22818 9777 -22768
rect 9321 -23140 9381 -22828
rect 9837 -22818 9847 -22768
rect 10223 -22698 10233 -22638
rect 10293 -22698 10303 -22638
rect 10223 -22768 10303 -22698
rect 10223 -22818 10233 -22768
rect 9777 -23140 9837 -22828
rect 10293 -22818 10303 -22768
rect 10681 -22698 10691 -22638
rect 10751 -22698 10761 -22638
rect 10681 -22768 10761 -22698
rect 10681 -22818 10691 -22768
rect 10233 -23140 10293 -22828
rect 10751 -22818 10761 -22768
rect 11137 -22698 11147 -22638
rect 11207 -22698 11217 -22638
rect 11137 -22768 11217 -22698
rect 11137 -22818 11147 -22768
rect 10691 -23140 10751 -22828
rect 11207 -22818 11217 -22768
rect 11593 -22698 11603 -22638
rect 11663 -22698 11673 -22638
rect 11593 -22768 11673 -22698
rect 11593 -22818 11603 -22768
rect 11147 -23140 11207 -22828
rect 11663 -22818 11673 -22768
rect 12051 -22698 12061 -22638
rect 12121 -22698 12131 -22638
rect 12051 -22768 12131 -22698
rect 12051 -22818 12061 -22768
rect 11603 -23140 11663 -22828
rect 12121 -22818 12131 -22768
rect 12507 -22698 12517 -22638
rect 12577 -22698 12587 -22638
rect 12507 -22768 12587 -22698
rect 12507 -22818 12517 -22768
rect 12061 -23140 12121 -22828
rect 12577 -22818 12587 -22768
rect 12963 -22698 12973 -22638
rect 13033 -22698 13043 -22638
rect 12963 -22768 13043 -22698
rect 12963 -22818 12973 -22768
rect 12517 -23140 12577 -22828
rect 13033 -22818 13043 -22768
rect 13421 -22698 13431 -22638
rect 13491 -22698 13501 -22638
rect 13421 -22768 13501 -22698
rect 13421 -22818 13431 -22768
rect 12973 -23140 13033 -22828
rect 13491 -22818 13501 -22768
rect 13877 -22698 13887 -22638
rect 13947 -22698 13957 -22638
rect 13877 -22768 13957 -22698
rect 13877 -22818 13887 -22768
rect 13431 -23140 13491 -22828
rect 13947 -22818 13957 -22768
rect 14333 -22698 14343 -22638
rect 14403 -22698 14413 -22638
rect 14333 -22768 14413 -22698
rect 14333 -22818 14343 -22768
rect 13887 -23140 13947 -22828
rect 14403 -22818 14413 -22768
rect 14791 -22698 14801 -22638
rect 14861 -22698 14871 -22638
rect 14791 -22768 14871 -22698
rect 14791 -22818 14801 -22768
rect 14343 -23140 14403 -22828
rect 14861 -22818 14871 -22768
rect 15247 -22698 15257 -22638
rect 15317 -22698 15327 -22638
rect 15247 -22768 15327 -22698
rect 15247 -22818 15257 -22768
rect 14801 -23140 14861 -22828
rect 15317 -22818 15327 -22768
rect 15257 -23140 15317 -22828
rect 161 -23200 171 -23140
rect 231 -23200 241 -23140
rect 161 -23270 241 -23200
rect 161 -23320 171 -23270
rect 231 -23320 241 -23270
rect 617 -23200 627 -23140
rect 687 -23200 697 -23140
rect 617 -23270 697 -23200
rect 617 -23320 627 -23270
rect 171 -23634 231 -23330
rect 687 -23320 697 -23270
rect 1073 -23200 1083 -23140
rect 1143 -23200 1153 -23140
rect 1073 -23270 1153 -23200
rect 1073 -23320 1083 -23270
rect 627 -23634 687 -23330
rect 1143 -23320 1153 -23270
rect 1531 -23200 1541 -23140
rect 1601 -23200 1611 -23140
rect 1531 -23270 1611 -23200
rect 1531 -23320 1541 -23270
rect 1083 -23634 1143 -23330
rect 1601 -23320 1611 -23270
rect 1987 -23200 1997 -23140
rect 2057 -23200 2067 -23140
rect 1987 -23270 2067 -23200
rect 1987 -23320 1997 -23270
rect 1541 -23634 1601 -23330
rect 2057 -23320 2067 -23270
rect 2443 -23200 2453 -23140
rect 2513 -23200 2523 -23140
rect 2443 -23270 2523 -23200
rect 2443 -23320 2453 -23270
rect 1997 -23634 2057 -23330
rect 2513 -23320 2523 -23270
rect 2901 -23200 2911 -23140
rect 2971 -23200 2981 -23140
rect 2901 -23270 2981 -23200
rect 2901 -23320 2911 -23270
rect 2453 -23634 2513 -23330
rect 2971 -23320 2981 -23270
rect 3357 -23200 3367 -23140
rect 3427 -23200 3437 -23140
rect 3357 -23270 3437 -23200
rect 3357 -23320 3367 -23270
rect 2911 -23634 2971 -23330
rect 3427 -23320 3437 -23270
rect 3813 -23200 3823 -23140
rect 3883 -23200 3893 -23140
rect 3813 -23270 3893 -23200
rect 3813 -23320 3823 -23270
rect 3367 -23634 3427 -23330
rect 3883 -23320 3893 -23270
rect 4271 -23200 4281 -23140
rect 4341 -23200 4351 -23140
rect 4271 -23270 4351 -23200
rect 4271 -23320 4281 -23270
rect 3823 -23634 3883 -23330
rect 4341 -23320 4351 -23270
rect 4727 -23200 4737 -23140
rect 4797 -23200 4807 -23140
rect 4727 -23270 4807 -23200
rect 4727 -23320 4737 -23270
rect 4281 -23634 4341 -23330
rect 4797 -23320 4807 -23270
rect 5183 -23200 5193 -23140
rect 5253 -23200 5263 -23140
rect 5183 -23270 5263 -23200
rect 5183 -23320 5193 -23270
rect 4737 -23634 4797 -23330
rect 5253 -23320 5263 -23270
rect 5641 -23200 5651 -23140
rect 5711 -23200 5721 -23140
rect 5641 -23270 5721 -23200
rect 5641 -23320 5651 -23270
rect 5193 -23634 5253 -23330
rect 5711 -23320 5721 -23270
rect 6097 -23200 6107 -23140
rect 6167 -23200 6177 -23140
rect 6097 -23270 6177 -23200
rect 6097 -23320 6107 -23270
rect 5651 -23634 5711 -23330
rect 6167 -23320 6177 -23270
rect 6553 -23200 6563 -23140
rect 6623 -23200 6633 -23140
rect 6553 -23270 6633 -23200
rect 6553 -23320 6563 -23270
rect 6107 -23634 6167 -23330
rect 6623 -23320 6633 -23270
rect 7011 -23200 7021 -23140
rect 7081 -23200 7091 -23140
rect 7011 -23270 7091 -23200
rect 7011 -23320 7021 -23270
rect 6563 -23634 6623 -23330
rect 7081 -23320 7091 -23270
rect 7467 -23200 7477 -23140
rect 7537 -23200 7547 -23140
rect 7467 -23270 7547 -23200
rect 7467 -23320 7477 -23270
rect 7021 -23634 7081 -23330
rect 7537 -23320 7547 -23270
rect 7923 -23200 7933 -23140
rect 7993 -23200 8003 -23140
rect 7923 -23270 8003 -23200
rect 7923 -23320 7933 -23270
rect 7477 -23634 7537 -23330
rect 7993 -23320 8003 -23270
rect 8397 -23200 8407 -23140
rect 8467 -23200 8477 -23140
rect 8397 -23270 8477 -23200
rect 8397 -23320 8407 -23270
rect 7933 -23634 7993 -23330
rect 8467 -23320 8477 -23270
rect 8853 -23200 8863 -23140
rect 8923 -23200 8933 -23140
rect 8853 -23270 8933 -23200
rect 8853 -23320 8863 -23270
rect 8407 -23634 8467 -23330
rect 8923 -23320 8933 -23270
rect 9311 -23200 9321 -23140
rect 9381 -23200 9391 -23140
rect 9311 -23270 9391 -23200
rect 9311 -23320 9321 -23270
rect 8863 -23634 8923 -23330
rect 9381 -23320 9391 -23270
rect 9767 -23200 9777 -23140
rect 9837 -23200 9847 -23140
rect 9767 -23270 9847 -23200
rect 9767 -23320 9777 -23270
rect 9321 -23634 9381 -23330
rect 9837 -23320 9847 -23270
rect 10223 -23200 10233 -23140
rect 10293 -23200 10303 -23140
rect 10223 -23270 10303 -23200
rect 10223 -23320 10233 -23270
rect 9777 -23634 9837 -23330
rect 10293 -23320 10303 -23270
rect 10681 -23200 10691 -23140
rect 10751 -23200 10761 -23140
rect 10681 -23270 10761 -23200
rect 10681 -23320 10691 -23270
rect 10233 -23634 10293 -23330
rect 10751 -23320 10761 -23270
rect 11137 -23200 11147 -23140
rect 11207 -23200 11217 -23140
rect 11137 -23270 11217 -23200
rect 11137 -23320 11147 -23270
rect 10691 -23634 10751 -23330
rect 11207 -23320 11217 -23270
rect 11593 -23200 11603 -23140
rect 11663 -23200 11673 -23140
rect 11593 -23270 11673 -23200
rect 11593 -23320 11603 -23270
rect 11147 -23634 11207 -23330
rect 11663 -23320 11673 -23270
rect 12051 -23200 12061 -23140
rect 12121 -23200 12131 -23140
rect 12051 -23270 12131 -23200
rect 12051 -23320 12061 -23270
rect 11603 -23634 11663 -23330
rect 12121 -23320 12131 -23270
rect 12507 -23200 12517 -23140
rect 12577 -23200 12587 -23140
rect 12507 -23270 12587 -23200
rect 12507 -23320 12517 -23270
rect 12061 -23634 12121 -23330
rect 12577 -23320 12587 -23270
rect 12963 -23200 12973 -23140
rect 13033 -23200 13043 -23140
rect 12963 -23270 13043 -23200
rect 12963 -23320 12973 -23270
rect 12517 -23634 12577 -23330
rect 13033 -23320 13043 -23270
rect 13421 -23200 13431 -23140
rect 13491 -23200 13501 -23140
rect 13421 -23270 13501 -23200
rect 13421 -23320 13431 -23270
rect 12973 -23634 13033 -23330
rect 13491 -23320 13501 -23270
rect 13877 -23200 13887 -23140
rect 13947 -23200 13957 -23140
rect 13877 -23270 13957 -23200
rect 13877 -23320 13887 -23270
rect 13431 -23634 13491 -23330
rect 13947 -23320 13957 -23270
rect 14333 -23200 14343 -23140
rect 14403 -23200 14413 -23140
rect 14333 -23270 14413 -23200
rect 14333 -23320 14343 -23270
rect 13887 -23634 13947 -23330
rect 14403 -23320 14413 -23270
rect 14791 -23200 14801 -23140
rect 14861 -23200 14871 -23140
rect 14791 -23270 14871 -23200
rect 14791 -23320 14801 -23270
rect 14343 -23634 14403 -23330
rect 14861 -23320 14871 -23270
rect 15247 -23200 15257 -23140
rect 15317 -23200 15327 -23140
rect 15247 -23270 15327 -23200
rect 15247 -23320 15257 -23270
rect 14801 -23634 14861 -23330
rect 15317 -23320 15327 -23270
rect 15257 -23634 15317 -23330
rect 161 -23694 171 -23634
rect 231 -23694 241 -23634
rect 161 -23764 241 -23694
rect 161 -23814 171 -23764
rect 231 -23814 241 -23764
rect 617 -23694 627 -23634
rect 687 -23694 697 -23634
rect 617 -23764 697 -23694
rect 617 -23814 627 -23764
rect 171 -24126 231 -23824
rect 687 -23814 697 -23764
rect 1073 -23694 1083 -23634
rect 1143 -23694 1153 -23634
rect 1073 -23764 1153 -23694
rect 1073 -23814 1083 -23764
rect 627 -24126 687 -23824
rect 1143 -23814 1153 -23764
rect 1531 -23694 1541 -23634
rect 1601 -23694 1611 -23634
rect 1531 -23764 1611 -23694
rect 1531 -23814 1541 -23764
rect 1083 -24126 1143 -23824
rect 1601 -23814 1611 -23764
rect 1987 -23694 1997 -23634
rect 2057 -23694 2067 -23634
rect 1987 -23764 2067 -23694
rect 1987 -23814 1997 -23764
rect 1541 -24126 1601 -23824
rect 2057 -23814 2067 -23764
rect 2443 -23694 2453 -23634
rect 2513 -23694 2523 -23634
rect 2443 -23764 2523 -23694
rect 2443 -23814 2453 -23764
rect 1997 -24126 2057 -23824
rect 2513 -23814 2523 -23764
rect 2901 -23694 2911 -23634
rect 2971 -23694 2981 -23634
rect 2901 -23764 2981 -23694
rect 2901 -23814 2911 -23764
rect 2453 -24126 2513 -23824
rect 2971 -23814 2981 -23764
rect 3357 -23694 3367 -23634
rect 3427 -23694 3437 -23634
rect 3357 -23764 3437 -23694
rect 3357 -23814 3367 -23764
rect 2911 -24126 2971 -23824
rect 3427 -23814 3437 -23764
rect 3813 -23694 3823 -23634
rect 3883 -23694 3893 -23634
rect 3813 -23764 3893 -23694
rect 3813 -23814 3823 -23764
rect 3367 -24126 3427 -23824
rect 3883 -23814 3893 -23764
rect 4271 -23694 4281 -23634
rect 4341 -23694 4351 -23634
rect 4271 -23764 4351 -23694
rect 4271 -23814 4281 -23764
rect 3823 -24126 3883 -23824
rect 4341 -23814 4351 -23764
rect 4727 -23694 4737 -23634
rect 4797 -23694 4807 -23634
rect 4727 -23764 4807 -23694
rect 4727 -23814 4737 -23764
rect 4281 -24126 4341 -23824
rect 4797 -23814 4807 -23764
rect 5183 -23694 5193 -23634
rect 5253 -23694 5263 -23634
rect 5183 -23764 5263 -23694
rect 5183 -23814 5193 -23764
rect 4737 -24126 4797 -23824
rect 5253 -23814 5263 -23764
rect 5641 -23694 5651 -23634
rect 5711 -23694 5721 -23634
rect 5641 -23764 5721 -23694
rect 5641 -23814 5651 -23764
rect 5193 -24126 5253 -23824
rect 5711 -23814 5721 -23764
rect 6097 -23694 6107 -23634
rect 6167 -23694 6177 -23634
rect 6097 -23764 6177 -23694
rect 6097 -23814 6107 -23764
rect 5651 -24126 5711 -23824
rect 6167 -23814 6177 -23764
rect 6553 -23694 6563 -23634
rect 6623 -23694 6633 -23634
rect 6553 -23764 6633 -23694
rect 6553 -23814 6563 -23764
rect 6107 -24126 6167 -23824
rect 6623 -23814 6633 -23764
rect 7011 -23694 7021 -23634
rect 7081 -23694 7091 -23634
rect 7011 -23764 7091 -23694
rect 7011 -23814 7021 -23764
rect 6563 -24126 6623 -23824
rect 7081 -23814 7091 -23764
rect 7467 -23694 7477 -23634
rect 7537 -23694 7547 -23634
rect 7467 -23764 7547 -23694
rect 7467 -23814 7477 -23764
rect 7021 -24126 7081 -23824
rect 7537 -23814 7547 -23764
rect 7923 -23694 7933 -23634
rect 7993 -23694 8003 -23634
rect 7923 -23764 8003 -23694
rect 7923 -23814 7933 -23764
rect 7477 -24126 7537 -23824
rect 7993 -23814 8003 -23764
rect 8397 -23694 8407 -23634
rect 8467 -23694 8477 -23634
rect 8397 -23764 8477 -23694
rect 8397 -23814 8407 -23764
rect 7933 -24126 7993 -23824
rect 8467 -23814 8477 -23764
rect 8853 -23694 8863 -23634
rect 8923 -23694 8933 -23634
rect 8853 -23764 8933 -23694
rect 8853 -23814 8863 -23764
rect 8407 -24126 8467 -23824
rect 8923 -23814 8933 -23764
rect 9311 -23694 9321 -23634
rect 9381 -23694 9391 -23634
rect 9311 -23764 9391 -23694
rect 9311 -23814 9321 -23764
rect 8863 -24126 8923 -23824
rect 9381 -23814 9391 -23764
rect 9767 -23694 9777 -23634
rect 9837 -23694 9847 -23634
rect 9767 -23764 9847 -23694
rect 9767 -23814 9777 -23764
rect 9321 -24126 9381 -23824
rect 9837 -23814 9847 -23764
rect 10223 -23694 10233 -23634
rect 10293 -23694 10303 -23634
rect 10223 -23764 10303 -23694
rect 10223 -23814 10233 -23764
rect 9777 -24126 9837 -23824
rect 10293 -23814 10303 -23764
rect 10681 -23694 10691 -23634
rect 10751 -23694 10761 -23634
rect 10681 -23764 10761 -23694
rect 10681 -23814 10691 -23764
rect 10233 -24126 10293 -23824
rect 10751 -23814 10761 -23764
rect 11137 -23694 11147 -23634
rect 11207 -23694 11217 -23634
rect 11137 -23764 11217 -23694
rect 11137 -23814 11147 -23764
rect 10691 -24126 10751 -23824
rect 11207 -23814 11217 -23764
rect 11593 -23694 11603 -23634
rect 11663 -23694 11673 -23634
rect 11593 -23764 11673 -23694
rect 11593 -23814 11603 -23764
rect 11147 -24126 11207 -23824
rect 11663 -23814 11673 -23764
rect 12051 -23694 12061 -23634
rect 12121 -23694 12131 -23634
rect 12051 -23764 12131 -23694
rect 12051 -23814 12061 -23764
rect 11603 -24126 11663 -23824
rect 12121 -23814 12131 -23764
rect 12507 -23694 12517 -23634
rect 12577 -23694 12587 -23634
rect 12507 -23764 12587 -23694
rect 12507 -23814 12517 -23764
rect 12061 -24126 12121 -23824
rect 12577 -23814 12587 -23764
rect 12963 -23694 12973 -23634
rect 13033 -23694 13043 -23634
rect 12963 -23764 13043 -23694
rect 12963 -23814 12973 -23764
rect 12517 -24126 12577 -23824
rect 13033 -23814 13043 -23764
rect 13421 -23694 13431 -23634
rect 13491 -23694 13501 -23634
rect 13421 -23764 13501 -23694
rect 13421 -23814 13431 -23764
rect 12973 -24126 13033 -23824
rect 13491 -23814 13501 -23764
rect 13877 -23694 13887 -23634
rect 13947 -23694 13957 -23634
rect 13877 -23764 13957 -23694
rect 13877 -23814 13887 -23764
rect 13431 -24126 13491 -23824
rect 13947 -23814 13957 -23764
rect 14333 -23694 14343 -23634
rect 14403 -23694 14413 -23634
rect 14333 -23764 14413 -23694
rect 14333 -23814 14343 -23764
rect 13887 -24126 13947 -23824
rect 14403 -23814 14413 -23764
rect 14791 -23694 14801 -23634
rect 14861 -23694 14871 -23634
rect 14791 -23764 14871 -23694
rect 14791 -23814 14801 -23764
rect 14343 -24126 14403 -23824
rect 14861 -23814 14871 -23764
rect 15247 -23694 15257 -23634
rect 15317 -23694 15327 -23634
rect 15247 -23764 15327 -23694
rect 15247 -23814 15257 -23764
rect 14801 -24126 14861 -23824
rect 15317 -23814 15327 -23764
rect 15257 -24126 15317 -23824
rect 161 -24186 171 -24126
rect 231 -24186 241 -24126
rect 161 -24256 241 -24186
rect 161 -24306 171 -24256
rect 231 -24306 241 -24256
rect 617 -24186 627 -24126
rect 687 -24186 697 -24126
rect 617 -24256 697 -24186
rect 617 -24306 627 -24256
rect 171 -24628 231 -24316
rect 687 -24306 697 -24256
rect 1073 -24186 1083 -24126
rect 1143 -24186 1153 -24126
rect 1073 -24256 1153 -24186
rect 1073 -24306 1083 -24256
rect 627 -24628 687 -24316
rect 1143 -24306 1153 -24256
rect 1531 -24186 1541 -24126
rect 1601 -24186 1611 -24126
rect 1531 -24256 1611 -24186
rect 1531 -24306 1541 -24256
rect 1083 -24628 1143 -24316
rect 1601 -24306 1611 -24256
rect 1987 -24186 1997 -24126
rect 2057 -24186 2067 -24126
rect 1987 -24256 2067 -24186
rect 1987 -24306 1997 -24256
rect 1541 -24628 1601 -24316
rect 2057 -24306 2067 -24256
rect 2443 -24186 2453 -24126
rect 2513 -24186 2523 -24126
rect 2443 -24256 2523 -24186
rect 2443 -24306 2453 -24256
rect 1997 -24628 2057 -24316
rect 2513 -24306 2523 -24256
rect 2901 -24186 2911 -24126
rect 2971 -24186 2981 -24126
rect 2901 -24256 2981 -24186
rect 2901 -24306 2911 -24256
rect 2453 -24628 2513 -24316
rect 2971 -24306 2981 -24256
rect 3357 -24186 3367 -24126
rect 3427 -24186 3437 -24126
rect 3357 -24256 3437 -24186
rect 3357 -24306 3367 -24256
rect 2911 -24628 2971 -24316
rect 3427 -24306 3437 -24256
rect 3813 -24186 3823 -24126
rect 3883 -24186 3893 -24126
rect 3813 -24256 3893 -24186
rect 3813 -24306 3823 -24256
rect 3367 -24628 3427 -24316
rect 3883 -24306 3893 -24256
rect 4271 -24186 4281 -24126
rect 4341 -24186 4351 -24126
rect 4271 -24256 4351 -24186
rect 4271 -24306 4281 -24256
rect 3823 -24628 3883 -24316
rect 4341 -24306 4351 -24256
rect 4727 -24186 4737 -24126
rect 4797 -24186 4807 -24126
rect 4727 -24256 4807 -24186
rect 4727 -24306 4737 -24256
rect 4281 -24628 4341 -24316
rect 4797 -24306 4807 -24256
rect 5183 -24186 5193 -24126
rect 5253 -24186 5263 -24126
rect 5183 -24256 5263 -24186
rect 5183 -24306 5193 -24256
rect 4737 -24628 4797 -24316
rect 5253 -24306 5263 -24256
rect 5641 -24186 5651 -24126
rect 5711 -24186 5721 -24126
rect 5641 -24256 5721 -24186
rect 5641 -24306 5651 -24256
rect 5193 -24628 5253 -24316
rect 5711 -24306 5721 -24256
rect 6097 -24186 6107 -24126
rect 6167 -24186 6177 -24126
rect 6097 -24256 6177 -24186
rect 6097 -24306 6107 -24256
rect 5651 -24628 5711 -24316
rect 6167 -24306 6177 -24256
rect 6553 -24186 6563 -24126
rect 6623 -24186 6633 -24126
rect 6553 -24256 6633 -24186
rect 6553 -24306 6563 -24256
rect 6107 -24628 6167 -24316
rect 6623 -24306 6633 -24256
rect 7011 -24186 7021 -24126
rect 7081 -24186 7091 -24126
rect 7011 -24256 7091 -24186
rect 7011 -24306 7021 -24256
rect 6563 -24628 6623 -24316
rect 7081 -24306 7091 -24256
rect 7467 -24186 7477 -24126
rect 7537 -24186 7547 -24126
rect 7467 -24256 7547 -24186
rect 7467 -24306 7477 -24256
rect 7021 -24628 7081 -24316
rect 7537 -24306 7547 -24256
rect 7923 -24186 7933 -24126
rect 7993 -24186 8003 -24126
rect 7923 -24256 8003 -24186
rect 7923 -24306 7933 -24256
rect 7477 -24628 7537 -24316
rect 7993 -24306 8003 -24256
rect 8397 -24186 8407 -24126
rect 8467 -24186 8477 -24126
rect 8397 -24256 8477 -24186
rect 8397 -24306 8407 -24256
rect 7933 -24628 7993 -24316
rect 8467 -24306 8477 -24256
rect 8853 -24186 8863 -24126
rect 8923 -24186 8933 -24126
rect 8853 -24256 8933 -24186
rect 8853 -24306 8863 -24256
rect 8407 -24628 8467 -24316
rect 8923 -24306 8933 -24256
rect 9311 -24186 9321 -24126
rect 9381 -24186 9391 -24126
rect 9311 -24256 9391 -24186
rect 9311 -24306 9321 -24256
rect 8863 -24628 8923 -24316
rect 9381 -24306 9391 -24256
rect 9767 -24186 9777 -24126
rect 9837 -24186 9847 -24126
rect 9767 -24256 9847 -24186
rect 9767 -24306 9777 -24256
rect 9321 -24628 9381 -24316
rect 9837 -24306 9847 -24256
rect 10223 -24186 10233 -24126
rect 10293 -24186 10303 -24126
rect 10223 -24256 10303 -24186
rect 10223 -24306 10233 -24256
rect 9777 -24628 9837 -24316
rect 10293 -24306 10303 -24256
rect 10681 -24186 10691 -24126
rect 10751 -24186 10761 -24126
rect 10681 -24256 10761 -24186
rect 10681 -24306 10691 -24256
rect 10233 -24628 10293 -24316
rect 10751 -24306 10761 -24256
rect 11137 -24186 11147 -24126
rect 11207 -24186 11217 -24126
rect 11137 -24256 11217 -24186
rect 11137 -24306 11147 -24256
rect 10691 -24628 10751 -24316
rect 11207 -24306 11217 -24256
rect 11593 -24186 11603 -24126
rect 11663 -24186 11673 -24126
rect 11593 -24256 11673 -24186
rect 11593 -24306 11603 -24256
rect 11147 -24628 11207 -24316
rect 11663 -24306 11673 -24256
rect 12051 -24186 12061 -24126
rect 12121 -24186 12131 -24126
rect 12051 -24256 12131 -24186
rect 12051 -24306 12061 -24256
rect 11603 -24628 11663 -24316
rect 12121 -24306 12131 -24256
rect 12507 -24186 12517 -24126
rect 12577 -24186 12587 -24126
rect 12507 -24256 12587 -24186
rect 12507 -24306 12517 -24256
rect 12061 -24628 12121 -24316
rect 12577 -24306 12587 -24256
rect 12963 -24186 12973 -24126
rect 13033 -24186 13043 -24126
rect 12963 -24256 13043 -24186
rect 12963 -24306 12973 -24256
rect 12517 -24628 12577 -24316
rect 13033 -24306 13043 -24256
rect 13421 -24186 13431 -24126
rect 13491 -24186 13501 -24126
rect 13421 -24256 13501 -24186
rect 13421 -24306 13431 -24256
rect 12973 -24628 13033 -24316
rect 13491 -24306 13501 -24256
rect 13877 -24186 13887 -24126
rect 13947 -24186 13957 -24126
rect 13877 -24256 13957 -24186
rect 13877 -24306 13887 -24256
rect 13431 -24628 13491 -24316
rect 13947 -24306 13957 -24256
rect 14333 -24186 14343 -24126
rect 14403 -24186 14413 -24126
rect 14333 -24256 14413 -24186
rect 14333 -24306 14343 -24256
rect 13887 -24628 13947 -24316
rect 14403 -24306 14413 -24256
rect 14791 -24186 14801 -24126
rect 14861 -24186 14871 -24126
rect 14791 -24256 14871 -24186
rect 14791 -24306 14801 -24256
rect 14343 -24628 14403 -24316
rect 14861 -24306 14871 -24256
rect 15247 -24186 15257 -24126
rect 15317 -24186 15327 -24126
rect 15247 -24256 15327 -24186
rect 15247 -24306 15257 -24256
rect 14801 -24628 14861 -24316
rect 15317 -24306 15327 -24256
rect 15257 -24628 15317 -24316
rect 161 -24688 171 -24628
rect 231 -24688 241 -24628
rect 161 -24758 241 -24688
rect 161 -24808 171 -24758
rect 231 -24808 241 -24758
rect 617 -24688 627 -24628
rect 687 -24688 697 -24628
rect 617 -24758 697 -24688
rect 617 -24808 627 -24758
rect 171 -25144 231 -24818
rect 687 -24808 697 -24758
rect 1073 -24688 1083 -24628
rect 1143 -24688 1153 -24628
rect 1073 -24758 1153 -24688
rect 1073 -24808 1083 -24758
rect 627 -25144 687 -24818
rect 1143 -24808 1153 -24758
rect 1531 -24688 1541 -24628
rect 1601 -24688 1611 -24628
rect 1531 -24758 1611 -24688
rect 1531 -24808 1541 -24758
rect 1083 -25144 1143 -24818
rect 1601 -24808 1611 -24758
rect 1987 -24688 1997 -24628
rect 2057 -24688 2067 -24628
rect 1987 -24758 2067 -24688
rect 1987 -24808 1997 -24758
rect 1541 -25144 1601 -24818
rect 2057 -24808 2067 -24758
rect 2443 -24688 2453 -24628
rect 2513 -24688 2523 -24628
rect 2443 -24758 2523 -24688
rect 2443 -24808 2453 -24758
rect 1997 -25144 2057 -24818
rect 2513 -24808 2523 -24758
rect 2901 -24688 2911 -24628
rect 2971 -24688 2981 -24628
rect 2901 -24758 2981 -24688
rect 2901 -24808 2911 -24758
rect 2453 -25144 2513 -24818
rect 2971 -24808 2981 -24758
rect 3357 -24688 3367 -24628
rect 3427 -24688 3437 -24628
rect 3357 -24758 3437 -24688
rect 3357 -24808 3367 -24758
rect 2911 -25144 2971 -24818
rect 3427 -24808 3437 -24758
rect 3813 -24688 3823 -24628
rect 3883 -24688 3893 -24628
rect 3813 -24758 3893 -24688
rect 3813 -24808 3823 -24758
rect 3367 -25144 3427 -24818
rect 3883 -24808 3893 -24758
rect 4271 -24688 4281 -24628
rect 4341 -24688 4351 -24628
rect 4271 -24758 4351 -24688
rect 4271 -24808 4281 -24758
rect 3823 -25144 3883 -24818
rect 4341 -24808 4351 -24758
rect 4727 -24688 4737 -24628
rect 4797 -24688 4807 -24628
rect 4727 -24758 4807 -24688
rect 4727 -24808 4737 -24758
rect 4281 -25144 4341 -24818
rect 4797 -24808 4807 -24758
rect 5183 -24688 5193 -24628
rect 5253 -24688 5263 -24628
rect 5183 -24758 5263 -24688
rect 5183 -24808 5193 -24758
rect 4737 -25144 4797 -24818
rect 5253 -24808 5263 -24758
rect 5641 -24688 5651 -24628
rect 5711 -24688 5721 -24628
rect 5641 -24758 5721 -24688
rect 5641 -24808 5651 -24758
rect 5193 -25144 5253 -24818
rect 5711 -24808 5721 -24758
rect 6097 -24688 6107 -24628
rect 6167 -24688 6177 -24628
rect 6097 -24758 6177 -24688
rect 6097 -24808 6107 -24758
rect 5651 -25144 5711 -24818
rect 6167 -24808 6177 -24758
rect 6553 -24688 6563 -24628
rect 6623 -24688 6633 -24628
rect 6553 -24758 6633 -24688
rect 6553 -24808 6563 -24758
rect 6107 -25144 6167 -24818
rect 6623 -24808 6633 -24758
rect 7011 -24688 7021 -24628
rect 7081 -24688 7091 -24628
rect 7011 -24758 7091 -24688
rect 7011 -24808 7021 -24758
rect 6563 -25144 6623 -24818
rect 7081 -24808 7091 -24758
rect 7467 -24688 7477 -24628
rect 7537 -24688 7547 -24628
rect 7467 -24758 7547 -24688
rect 7467 -24808 7477 -24758
rect 7021 -25144 7081 -24818
rect 7537 -24808 7547 -24758
rect 7923 -24688 7933 -24628
rect 7993 -24688 8003 -24628
rect 7923 -24758 8003 -24688
rect 7923 -24808 7933 -24758
rect 7477 -25144 7537 -24818
rect 7993 -24808 8003 -24758
rect 8397 -24688 8407 -24628
rect 8467 -24688 8477 -24628
rect 8397 -24758 8477 -24688
rect 8397 -24808 8407 -24758
rect 7933 -25144 7993 -24818
rect 8467 -24808 8477 -24758
rect 8853 -24688 8863 -24628
rect 8923 -24688 8933 -24628
rect 8853 -24758 8933 -24688
rect 8853 -24808 8863 -24758
rect 8407 -25144 8467 -24818
rect 8923 -24808 8933 -24758
rect 9311 -24688 9321 -24628
rect 9381 -24688 9391 -24628
rect 9311 -24758 9391 -24688
rect 9311 -24808 9321 -24758
rect 8863 -25144 8923 -24818
rect 9381 -24808 9391 -24758
rect 9767 -24688 9777 -24628
rect 9837 -24688 9847 -24628
rect 9767 -24758 9847 -24688
rect 9767 -24808 9777 -24758
rect 9321 -25144 9381 -24818
rect 9837 -24808 9847 -24758
rect 10223 -24688 10233 -24628
rect 10293 -24688 10303 -24628
rect 10223 -24758 10303 -24688
rect 10223 -24808 10233 -24758
rect 9777 -25144 9837 -24818
rect 10293 -24808 10303 -24758
rect 10681 -24688 10691 -24628
rect 10751 -24688 10761 -24628
rect 10681 -24758 10761 -24688
rect 10681 -24808 10691 -24758
rect 10233 -25144 10293 -24818
rect 10751 -24808 10761 -24758
rect 11137 -24688 11147 -24628
rect 11207 -24688 11217 -24628
rect 11137 -24758 11217 -24688
rect 11137 -24808 11147 -24758
rect 10691 -25144 10751 -24818
rect 11207 -24808 11217 -24758
rect 11593 -24688 11603 -24628
rect 11663 -24688 11673 -24628
rect 11593 -24758 11673 -24688
rect 11593 -24808 11603 -24758
rect 11147 -25144 11207 -24818
rect 11663 -24808 11673 -24758
rect 12051 -24688 12061 -24628
rect 12121 -24688 12131 -24628
rect 12051 -24758 12131 -24688
rect 12051 -24808 12061 -24758
rect 11603 -25144 11663 -24818
rect 12121 -24808 12131 -24758
rect 12507 -24688 12517 -24628
rect 12577 -24688 12587 -24628
rect 12507 -24758 12587 -24688
rect 12507 -24808 12517 -24758
rect 12061 -25144 12121 -24818
rect 12577 -24808 12587 -24758
rect 12963 -24688 12973 -24628
rect 13033 -24688 13043 -24628
rect 12963 -24758 13043 -24688
rect 12963 -24808 12973 -24758
rect 12517 -25144 12577 -24818
rect 13033 -24808 13043 -24758
rect 13421 -24688 13431 -24628
rect 13491 -24688 13501 -24628
rect 13421 -24758 13501 -24688
rect 13421 -24808 13431 -24758
rect 12973 -25144 13033 -24818
rect 13491 -24808 13501 -24758
rect 13877 -24688 13887 -24628
rect 13947 -24688 13957 -24628
rect 13877 -24758 13957 -24688
rect 13877 -24808 13887 -24758
rect 13431 -25144 13491 -24818
rect 13947 -24808 13957 -24758
rect 14333 -24688 14343 -24628
rect 14403 -24688 14413 -24628
rect 14333 -24758 14413 -24688
rect 14333 -24808 14343 -24758
rect 13887 -25144 13947 -24818
rect 14403 -24808 14413 -24758
rect 14791 -24688 14801 -24628
rect 14861 -24688 14871 -24628
rect 14791 -24758 14871 -24688
rect 14791 -24808 14801 -24758
rect 14343 -25144 14403 -24818
rect 14861 -24808 14871 -24758
rect 15247 -24688 15257 -24628
rect 15317 -24688 15327 -24628
rect 15247 -24758 15327 -24688
rect 15247 -24808 15257 -24758
rect 14801 -25144 14861 -24818
rect 15317 -24808 15327 -24758
rect 15257 -25144 15317 -24818
rect 161 -25204 171 -25144
rect 231 -25204 241 -25144
rect 161 -25274 241 -25204
rect 161 -25324 171 -25274
rect 231 -25324 241 -25274
rect 617 -25204 627 -25144
rect 687 -25204 697 -25144
rect 617 -25274 697 -25204
rect 617 -25324 627 -25274
rect 171 -25636 231 -25334
rect 687 -25324 697 -25274
rect 1073 -25204 1083 -25144
rect 1143 -25204 1153 -25144
rect 1073 -25274 1153 -25204
rect 1073 -25324 1083 -25274
rect 627 -25636 687 -25334
rect 1143 -25324 1153 -25274
rect 1531 -25204 1541 -25144
rect 1601 -25204 1611 -25144
rect 1531 -25274 1611 -25204
rect 1531 -25324 1541 -25274
rect 1083 -25636 1143 -25334
rect 1601 -25324 1611 -25274
rect 1987 -25204 1997 -25144
rect 2057 -25204 2067 -25144
rect 1987 -25274 2067 -25204
rect 1987 -25324 1997 -25274
rect 1541 -25636 1601 -25334
rect 2057 -25324 2067 -25274
rect 2443 -25204 2453 -25144
rect 2513 -25204 2523 -25144
rect 2443 -25274 2523 -25204
rect 2443 -25324 2453 -25274
rect 1997 -25636 2057 -25334
rect 2513 -25324 2523 -25274
rect 2901 -25204 2911 -25144
rect 2971 -25204 2981 -25144
rect 2901 -25274 2981 -25204
rect 2901 -25324 2911 -25274
rect 2453 -25636 2513 -25334
rect 2971 -25324 2981 -25274
rect 3357 -25204 3367 -25144
rect 3427 -25204 3437 -25144
rect 3357 -25274 3437 -25204
rect 3357 -25324 3367 -25274
rect 2911 -25636 2971 -25334
rect 3427 -25324 3437 -25274
rect 3813 -25204 3823 -25144
rect 3883 -25204 3893 -25144
rect 3813 -25274 3893 -25204
rect 3813 -25324 3823 -25274
rect 3367 -25636 3427 -25334
rect 3883 -25324 3893 -25274
rect 4271 -25204 4281 -25144
rect 4341 -25204 4351 -25144
rect 4271 -25274 4351 -25204
rect 4271 -25324 4281 -25274
rect 3823 -25636 3883 -25334
rect 4341 -25324 4351 -25274
rect 4727 -25204 4737 -25144
rect 4797 -25204 4807 -25144
rect 4727 -25274 4807 -25204
rect 4727 -25324 4737 -25274
rect 4281 -25636 4341 -25334
rect 4797 -25324 4807 -25274
rect 5183 -25204 5193 -25144
rect 5253 -25204 5263 -25144
rect 5183 -25274 5263 -25204
rect 5183 -25324 5193 -25274
rect 4737 -25636 4797 -25334
rect 5253 -25324 5263 -25274
rect 5641 -25204 5651 -25144
rect 5711 -25204 5721 -25144
rect 5641 -25274 5721 -25204
rect 5641 -25324 5651 -25274
rect 5193 -25636 5253 -25334
rect 5711 -25324 5721 -25274
rect 6097 -25204 6107 -25144
rect 6167 -25204 6177 -25144
rect 6097 -25274 6177 -25204
rect 6097 -25324 6107 -25274
rect 5651 -25636 5711 -25334
rect 6167 -25324 6177 -25274
rect 6553 -25204 6563 -25144
rect 6623 -25204 6633 -25144
rect 6553 -25274 6633 -25204
rect 6553 -25324 6563 -25274
rect 6107 -25636 6167 -25334
rect 6623 -25324 6633 -25274
rect 7011 -25204 7021 -25144
rect 7081 -25204 7091 -25144
rect 7011 -25274 7091 -25204
rect 7011 -25324 7021 -25274
rect 6563 -25636 6623 -25334
rect 7081 -25324 7091 -25274
rect 7467 -25204 7477 -25144
rect 7537 -25204 7547 -25144
rect 7467 -25274 7547 -25204
rect 7467 -25324 7477 -25274
rect 7021 -25636 7081 -25334
rect 7537 -25324 7547 -25274
rect 7923 -25204 7933 -25144
rect 7993 -25204 8003 -25144
rect 7923 -25274 8003 -25204
rect 7923 -25324 7933 -25274
rect 7477 -25636 7537 -25334
rect 7993 -25324 8003 -25274
rect 8397 -25204 8407 -25144
rect 8467 -25204 8477 -25144
rect 8397 -25274 8477 -25204
rect 8397 -25324 8407 -25274
rect 7933 -25636 7993 -25334
rect 8467 -25324 8477 -25274
rect 8853 -25204 8863 -25144
rect 8923 -25204 8933 -25144
rect 8853 -25274 8933 -25204
rect 8853 -25324 8863 -25274
rect 8407 -25636 8467 -25334
rect 8923 -25324 8933 -25274
rect 9311 -25204 9321 -25144
rect 9381 -25204 9391 -25144
rect 9311 -25274 9391 -25204
rect 9311 -25324 9321 -25274
rect 8863 -25636 8923 -25334
rect 9381 -25324 9391 -25274
rect 9767 -25204 9777 -25144
rect 9837 -25204 9847 -25144
rect 9767 -25274 9847 -25204
rect 9767 -25324 9777 -25274
rect 9321 -25636 9381 -25334
rect 9837 -25324 9847 -25274
rect 10223 -25204 10233 -25144
rect 10293 -25204 10303 -25144
rect 10223 -25274 10303 -25204
rect 10223 -25324 10233 -25274
rect 9777 -25636 9837 -25334
rect 10293 -25324 10303 -25274
rect 10681 -25204 10691 -25144
rect 10751 -25204 10761 -25144
rect 10681 -25274 10761 -25204
rect 10681 -25324 10691 -25274
rect 10233 -25636 10293 -25334
rect 10751 -25324 10761 -25274
rect 11137 -25204 11147 -25144
rect 11207 -25204 11217 -25144
rect 11137 -25274 11217 -25204
rect 11137 -25324 11147 -25274
rect 10691 -25636 10751 -25334
rect 11207 -25324 11217 -25274
rect 11593 -25204 11603 -25144
rect 11663 -25204 11673 -25144
rect 11593 -25274 11673 -25204
rect 11593 -25324 11603 -25274
rect 11147 -25636 11207 -25334
rect 11663 -25324 11673 -25274
rect 12051 -25204 12061 -25144
rect 12121 -25204 12131 -25144
rect 12051 -25274 12131 -25204
rect 12051 -25324 12061 -25274
rect 11603 -25636 11663 -25334
rect 12121 -25324 12131 -25274
rect 12507 -25204 12517 -25144
rect 12577 -25204 12587 -25144
rect 12507 -25274 12587 -25204
rect 12507 -25324 12517 -25274
rect 12061 -25636 12121 -25334
rect 12577 -25324 12587 -25274
rect 12963 -25204 12973 -25144
rect 13033 -25204 13043 -25144
rect 12963 -25274 13043 -25204
rect 12963 -25324 12973 -25274
rect 12517 -25636 12577 -25334
rect 13033 -25324 13043 -25274
rect 13421 -25204 13431 -25144
rect 13491 -25204 13501 -25144
rect 13421 -25274 13501 -25204
rect 13421 -25324 13431 -25274
rect 12973 -25636 13033 -25334
rect 13491 -25324 13501 -25274
rect 13877 -25204 13887 -25144
rect 13947 -25204 13957 -25144
rect 13877 -25274 13957 -25204
rect 13877 -25324 13887 -25274
rect 13431 -25636 13491 -25334
rect 13947 -25324 13957 -25274
rect 14333 -25204 14343 -25144
rect 14403 -25204 14413 -25144
rect 14333 -25274 14413 -25204
rect 14333 -25324 14343 -25274
rect 13887 -25636 13947 -25334
rect 14403 -25324 14413 -25274
rect 14791 -25204 14801 -25144
rect 14861 -25204 14871 -25144
rect 14791 -25274 14871 -25204
rect 14791 -25324 14801 -25274
rect 14343 -25636 14403 -25334
rect 14861 -25324 14871 -25274
rect 15247 -25204 15257 -25144
rect 15317 -25204 15327 -25144
rect 15247 -25274 15327 -25204
rect 15247 -25324 15257 -25274
rect 14801 -25636 14861 -25334
rect 15317 -25324 15327 -25274
rect 15257 -25636 15317 -25334
rect 161 -25696 171 -25636
rect 231 -25696 241 -25636
rect 161 -25766 241 -25696
rect 161 -25816 171 -25766
rect 231 -25816 241 -25766
rect 617 -25696 627 -25636
rect 687 -25696 697 -25636
rect 617 -25766 697 -25696
rect 617 -25816 627 -25766
rect 171 -25993 231 -25826
rect 687 -25816 697 -25766
rect 1073 -25696 1083 -25636
rect 1143 -25696 1153 -25636
rect 1073 -25766 1153 -25696
rect 1073 -25816 1083 -25766
rect 627 -25993 687 -25826
rect 1143 -25816 1153 -25766
rect 1531 -25696 1541 -25636
rect 1601 -25696 1611 -25636
rect 1531 -25766 1611 -25696
rect 1531 -25816 1541 -25766
rect 1083 -25993 1143 -25826
rect 1601 -25816 1611 -25766
rect 1987 -25696 1997 -25636
rect 2057 -25696 2067 -25636
rect 1987 -25766 2067 -25696
rect 1987 -25816 1997 -25766
rect 1541 -25993 1601 -25826
rect 2057 -25816 2067 -25766
rect 2443 -25696 2453 -25636
rect 2513 -25696 2523 -25636
rect 2443 -25766 2523 -25696
rect 2443 -25816 2453 -25766
rect 1997 -25993 2057 -25826
rect 2513 -25816 2523 -25766
rect 2901 -25696 2911 -25636
rect 2971 -25696 2981 -25636
rect 2901 -25766 2981 -25696
rect 2901 -25816 2911 -25766
rect 2453 -25993 2513 -25826
rect 2971 -25816 2981 -25766
rect 3357 -25696 3367 -25636
rect 3427 -25696 3437 -25636
rect 3357 -25766 3437 -25696
rect 3357 -25816 3367 -25766
rect 2911 -25993 2971 -25826
rect 3427 -25816 3437 -25766
rect 3813 -25696 3823 -25636
rect 3883 -25696 3893 -25636
rect 3813 -25766 3893 -25696
rect 3813 -25816 3823 -25766
rect 3367 -25993 3427 -25826
rect 3883 -25816 3893 -25766
rect 4271 -25696 4281 -25636
rect 4341 -25696 4351 -25636
rect 4271 -25766 4351 -25696
rect 4271 -25816 4281 -25766
rect 3823 -25993 3883 -25826
rect 4341 -25816 4351 -25766
rect 4727 -25696 4737 -25636
rect 4797 -25696 4807 -25636
rect 4727 -25766 4807 -25696
rect 4727 -25816 4737 -25766
rect 4281 -25993 4341 -25826
rect 4797 -25816 4807 -25766
rect 5183 -25696 5193 -25636
rect 5253 -25696 5263 -25636
rect 5183 -25766 5263 -25696
rect 5183 -25816 5193 -25766
rect 4737 -25993 4797 -25826
rect 5253 -25816 5263 -25766
rect 5641 -25696 5651 -25636
rect 5711 -25696 5721 -25636
rect 5641 -25766 5721 -25696
rect 5641 -25816 5651 -25766
rect 5193 -25993 5253 -25826
rect 5711 -25816 5721 -25766
rect 6097 -25696 6107 -25636
rect 6167 -25696 6177 -25636
rect 6097 -25766 6177 -25696
rect 6097 -25816 6107 -25766
rect 5651 -25993 5711 -25826
rect 6167 -25816 6177 -25766
rect 6553 -25696 6563 -25636
rect 6623 -25696 6633 -25636
rect 6553 -25766 6633 -25696
rect 6553 -25816 6563 -25766
rect 6107 -25993 6167 -25826
rect 6623 -25816 6633 -25766
rect 7011 -25696 7021 -25636
rect 7081 -25696 7091 -25636
rect 7011 -25766 7091 -25696
rect 7011 -25816 7021 -25766
rect 6563 -25993 6623 -25826
rect 7081 -25816 7091 -25766
rect 7467 -25696 7477 -25636
rect 7537 -25696 7547 -25636
rect 7467 -25766 7547 -25696
rect 7467 -25816 7477 -25766
rect 7021 -25993 7081 -25826
rect 7537 -25816 7547 -25766
rect 7923 -25696 7933 -25636
rect 7993 -25696 8003 -25636
rect 7923 -25766 8003 -25696
rect 7923 -25816 7933 -25766
rect 7477 -25993 7537 -25826
rect 7993 -25816 8003 -25766
rect 8397 -25696 8407 -25636
rect 8467 -25696 8477 -25636
rect 8397 -25766 8477 -25696
rect 8397 -25816 8407 -25766
rect 7933 -25993 7993 -25826
rect 8467 -25816 8477 -25766
rect 8853 -25696 8863 -25636
rect 8923 -25696 8933 -25636
rect 8853 -25766 8933 -25696
rect 8853 -25816 8863 -25766
rect 8407 -25993 8467 -25826
rect 8923 -25816 8933 -25766
rect 9311 -25696 9321 -25636
rect 9381 -25696 9391 -25636
rect 9311 -25766 9391 -25696
rect 9311 -25816 9321 -25766
rect 8863 -25993 8923 -25826
rect 9381 -25816 9391 -25766
rect 9767 -25696 9777 -25636
rect 9837 -25696 9847 -25636
rect 9767 -25766 9847 -25696
rect 9767 -25816 9777 -25766
rect 9321 -25993 9381 -25826
rect 9837 -25816 9847 -25766
rect 10223 -25696 10233 -25636
rect 10293 -25696 10303 -25636
rect 10223 -25766 10303 -25696
rect 10223 -25816 10233 -25766
rect 9777 -25993 9837 -25826
rect 10293 -25816 10303 -25766
rect 10681 -25696 10691 -25636
rect 10751 -25696 10761 -25636
rect 10681 -25766 10761 -25696
rect 10681 -25816 10691 -25766
rect 10233 -25993 10293 -25826
rect 10751 -25816 10761 -25766
rect 11137 -25696 11147 -25636
rect 11207 -25696 11217 -25636
rect 11137 -25766 11217 -25696
rect 11137 -25816 11147 -25766
rect 10691 -25993 10751 -25826
rect 11207 -25816 11217 -25766
rect 11593 -25696 11603 -25636
rect 11663 -25696 11673 -25636
rect 11593 -25766 11673 -25696
rect 11593 -25816 11603 -25766
rect 11147 -25993 11207 -25826
rect 11663 -25816 11673 -25766
rect 12051 -25696 12061 -25636
rect 12121 -25696 12131 -25636
rect 12051 -25766 12131 -25696
rect 12051 -25816 12061 -25766
rect 11603 -25993 11663 -25826
rect 12121 -25816 12131 -25766
rect 12507 -25696 12517 -25636
rect 12577 -25696 12587 -25636
rect 12507 -25766 12587 -25696
rect 12507 -25816 12517 -25766
rect 12061 -25993 12121 -25826
rect 12577 -25816 12587 -25766
rect 12963 -25696 12973 -25636
rect 13033 -25696 13043 -25636
rect 12963 -25766 13043 -25696
rect 12963 -25816 12973 -25766
rect 12517 -25993 12577 -25826
rect 13033 -25816 13043 -25766
rect 13421 -25696 13431 -25636
rect 13491 -25696 13501 -25636
rect 13421 -25766 13501 -25696
rect 13421 -25816 13431 -25766
rect 12973 -25993 13033 -25826
rect 13491 -25816 13501 -25766
rect 13877 -25696 13887 -25636
rect 13947 -25696 13957 -25636
rect 13877 -25766 13957 -25696
rect 13877 -25816 13887 -25766
rect 13431 -25993 13491 -25826
rect 13947 -25816 13957 -25766
rect 14333 -25696 14343 -25636
rect 14403 -25696 14413 -25636
rect 14333 -25766 14413 -25696
rect 14333 -25816 14343 -25766
rect 13887 -25993 13947 -25826
rect 14403 -25816 14413 -25766
rect 14791 -25696 14801 -25636
rect 14861 -25696 14871 -25636
rect 14791 -25766 14871 -25696
rect 14791 -25816 14801 -25766
rect 14343 -25993 14403 -25826
rect 14861 -25816 14871 -25766
rect 15247 -25696 15257 -25636
rect 15317 -25696 15327 -25636
rect 15247 -25766 15327 -25696
rect 15247 -25816 15257 -25766
rect 14801 -25993 14861 -25826
rect 15317 -25816 15327 -25766
rect 15257 -25993 15317 -25826
rect 170 -25997 231 -25993
rect 626 -25997 687 -25993
rect 1082 -25997 1143 -25993
rect 1540 -25997 1601 -25993
rect 1996 -25997 2057 -25993
rect 2452 -25997 2513 -25993
rect 2910 -25997 2971 -25993
rect 3366 -25997 3427 -25993
rect 3822 -25997 3883 -25993
rect 4280 -25997 4341 -25993
rect 4736 -25997 4797 -25993
rect 5192 -25997 5253 -25993
rect 5650 -25997 5711 -25993
rect 6106 -25997 6167 -25993
rect 6562 -25997 6623 -25993
rect 7020 -25997 7081 -25993
rect 7476 -25997 7537 -25993
rect 7932 -25997 7993 -25993
rect 8406 -25997 8467 -25993
rect 8862 -25997 8923 -25993
rect 9320 -25997 9381 -25993
rect 9776 -25997 9837 -25993
rect 10232 -25997 10293 -25993
rect 10690 -25997 10751 -25993
rect 11146 -25997 11207 -25993
rect 11602 -25997 11663 -25993
rect 12060 -25997 12121 -25993
rect 12516 -25997 12577 -25993
rect 12972 -25997 13033 -25993
rect 13430 -25997 13491 -25993
rect 13886 -25997 13947 -25993
rect 14342 -25997 14403 -25993
rect 14800 -25997 14861 -25993
rect 15256 -25997 15317 -25993
rect 170 -26133 230 -25997
rect 626 -26133 686 -25997
rect 1082 -26133 1142 -25997
rect 1540 -26133 1600 -25997
rect 1996 -26133 2056 -25997
rect 2452 -26133 2512 -25997
rect 2910 -26133 2970 -25997
rect 3366 -26133 3426 -25997
rect 3822 -26133 3882 -25997
rect 4280 -26133 4340 -25997
rect 4736 -26133 4796 -25997
rect 5192 -26133 5252 -25997
rect 5650 -26133 5710 -25997
rect 6106 -26133 6166 -25997
rect 6562 -26133 6622 -25997
rect 7020 -26133 7080 -25997
rect 7476 -26133 7536 -25997
rect 7932 -26133 7992 -25997
rect 8406 -26133 8466 -25997
rect 8862 -26133 8922 -25997
rect 9320 -26133 9380 -25997
rect 9776 -26133 9836 -25997
rect 10232 -26133 10292 -25997
rect 10690 -26133 10750 -25997
rect 11146 -26133 11206 -25997
rect 11602 -26133 11662 -25997
rect 12060 -26133 12120 -25997
rect 12516 -26133 12576 -25997
rect 12972 -26133 13032 -25997
rect 13430 -26133 13490 -25997
rect 13886 -26133 13946 -25997
rect 14342 -26133 14402 -25997
rect 14800 -26133 14860 -25997
rect 15256 -26133 15316 -25997
rect 160 -26193 170 -26133
rect 230 -26193 240 -26133
rect 160 -26263 240 -26193
rect 160 -26313 170 -26263
rect 230 -26313 240 -26263
rect 616 -26193 626 -26133
rect 686 -26193 696 -26133
rect 616 -26263 696 -26193
rect 616 -26313 626 -26263
rect 170 -26625 230 -26323
rect 686 -26313 696 -26263
rect 1072 -26193 1082 -26133
rect 1142 -26193 1152 -26133
rect 1072 -26263 1152 -26193
rect 1072 -26313 1082 -26263
rect 626 -26625 686 -26323
rect 1142 -26313 1152 -26263
rect 1530 -26193 1540 -26133
rect 1600 -26193 1610 -26133
rect 1530 -26263 1610 -26193
rect 1530 -26313 1540 -26263
rect 1082 -26625 1142 -26323
rect 1600 -26313 1610 -26263
rect 1986 -26193 1996 -26133
rect 2056 -26193 2066 -26133
rect 1986 -26263 2066 -26193
rect 1986 -26313 1996 -26263
rect 1540 -26625 1600 -26323
rect 2056 -26313 2066 -26263
rect 2442 -26193 2452 -26133
rect 2512 -26193 2522 -26133
rect 2442 -26263 2522 -26193
rect 2442 -26313 2452 -26263
rect 1996 -26625 2056 -26323
rect 2512 -26313 2522 -26263
rect 2900 -26193 2910 -26133
rect 2970 -26193 2980 -26133
rect 2900 -26263 2980 -26193
rect 2900 -26313 2910 -26263
rect 2452 -26625 2512 -26323
rect 2970 -26313 2980 -26263
rect 3356 -26193 3366 -26133
rect 3426 -26193 3436 -26133
rect 3356 -26263 3436 -26193
rect 3356 -26313 3366 -26263
rect 2910 -26625 2970 -26323
rect 3426 -26313 3436 -26263
rect 3812 -26193 3822 -26133
rect 3882 -26193 3892 -26133
rect 3812 -26263 3892 -26193
rect 3812 -26313 3822 -26263
rect 3366 -26625 3426 -26323
rect 3882 -26313 3892 -26263
rect 4270 -26193 4280 -26133
rect 4340 -26193 4350 -26133
rect 4270 -26263 4350 -26193
rect 4270 -26313 4280 -26263
rect 3822 -26625 3882 -26323
rect 4340 -26313 4350 -26263
rect 4726 -26193 4736 -26133
rect 4796 -26193 4806 -26133
rect 4726 -26263 4806 -26193
rect 4726 -26313 4736 -26263
rect 4280 -26625 4340 -26323
rect 4796 -26313 4806 -26263
rect 5182 -26193 5192 -26133
rect 5252 -26193 5262 -26133
rect 5182 -26263 5262 -26193
rect 5182 -26313 5192 -26263
rect 4736 -26625 4796 -26323
rect 5252 -26313 5262 -26263
rect 5640 -26193 5650 -26133
rect 5710 -26193 5720 -26133
rect 5640 -26263 5720 -26193
rect 5640 -26313 5650 -26263
rect 5192 -26625 5252 -26323
rect 5710 -26313 5720 -26263
rect 6096 -26193 6106 -26133
rect 6166 -26193 6176 -26133
rect 6096 -26263 6176 -26193
rect 6096 -26313 6106 -26263
rect 5650 -26625 5710 -26323
rect 6166 -26313 6176 -26263
rect 6552 -26193 6562 -26133
rect 6622 -26193 6632 -26133
rect 6552 -26263 6632 -26193
rect 6552 -26313 6562 -26263
rect 6106 -26625 6166 -26323
rect 6622 -26313 6632 -26263
rect 7010 -26193 7020 -26133
rect 7080 -26193 7090 -26133
rect 7010 -26263 7090 -26193
rect 7010 -26313 7020 -26263
rect 6562 -26625 6622 -26323
rect 7080 -26313 7090 -26263
rect 7466 -26193 7476 -26133
rect 7536 -26193 7546 -26133
rect 7466 -26263 7546 -26193
rect 7466 -26313 7476 -26263
rect 7020 -26625 7080 -26323
rect 7536 -26313 7546 -26263
rect 7922 -26193 7932 -26133
rect 7992 -26193 8002 -26133
rect 7922 -26263 8002 -26193
rect 7922 -26313 7932 -26263
rect 7476 -26625 7536 -26323
rect 7992 -26313 8002 -26263
rect 8396 -26193 8406 -26133
rect 8466 -26193 8476 -26133
rect 8396 -26263 8476 -26193
rect 8396 -26313 8406 -26263
rect 7932 -26625 7992 -26323
rect 8466 -26313 8476 -26263
rect 8852 -26193 8862 -26133
rect 8922 -26193 8932 -26133
rect 8852 -26263 8932 -26193
rect 8852 -26313 8862 -26263
rect 8406 -26625 8466 -26323
rect 8922 -26313 8932 -26263
rect 9310 -26193 9320 -26133
rect 9380 -26193 9390 -26133
rect 9310 -26263 9390 -26193
rect 9310 -26313 9320 -26263
rect 8862 -26625 8922 -26323
rect 9380 -26313 9390 -26263
rect 9766 -26193 9776 -26133
rect 9836 -26193 9846 -26133
rect 9766 -26263 9846 -26193
rect 9766 -26313 9776 -26263
rect 9320 -26625 9380 -26323
rect 9836 -26313 9846 -26263
rect 10222 -26193 10232 -26133
rect 10292 -26193 10302 -26133
rect 10222 -26263 10302 -26193
rect 10222 -26313 10232 -26263
rect 9776 -26625 9836 -26323
rect 10292 -26313 10302 -26263
rect 10680 -26193 10690 -26133
rect 10750 -26193 10760 -26133
rect 10680 -26263 10760 -26193
rect 10680 -26313 10690 -26263
rect 10232 -26625 10292 -26323
rect 10750 -26313 10760 -26263
rect 11136 -26193 11146 -26133
rect 11206 -26193 11216 -26133
rect 11136 -26263 11216 -26193
rect 11136 -26313 11146 -26263
rect 10690 -26625 10750 -26323
rect 11206 -26313 11216 -26263
rect 11592 -26193 11602 -26133
rect 11662 -26193 11672 -26133
rect 11592 -26263 11672 -26193
rect 11592 -26313 11602 -26263
rect 11146 -26625 11206 -26323
rect 11662 -26313 11672 -26263
rect 12050 -26193 12060 -26133
rect 12120 -26193 12130 -26133
rect 12050 -26263 12130 -26193
rect 12050 -26313 12060 -26263
rect 11602 -26625 11662 -26323
rect 12120 -26313 12130 -26263
rect 12506 -26193 12516 -26133
rect 12576 -26193 12586 -26133
rect 12506 -26263 12586 -26193
rect 12506 -26313 12516 -26263
rect 12060 -26625 12120 -26323
rect 12576 -26313 12586 -26263
rect 12962 -26193 12972 -26133
rect 13032 -26193 13042 -26133
rect 12962 -26263 13042 -26193
rect 12962 -26313 12972 -26263
rect 12516 -26625 12576 -26323
rect 13032 -26313 13042 -26263
rect 13420 -26193 13430 -26133
rect 13490 -26193 13500 -26133
rect 13420 -26263 13500 -26193
rect 13420 -26313 13430 -26263
rect 12972 -26625 13032 -26323
rect 13490 -26313 13500 -26263
rect 13876 -26193 13886 -26133
rect 13946 -26193 13956 -26133
rect 13876 -26263 13956 -26193
rect 13876 -26313 13886 -26263
rect 13430 -26625 13490 -26323
rect 13946 -26313 13956 -26263
rect 14332 -26193 14342 -26133
rect 14402 -26193 14412 -26133
rect 14332 -26263 14412 -26193
rect 14332 -26313 14342 -26263
rect 13886 -26625 13946 -26323
rect 14402 -26313 14412 -26263
rect 14790 -26193 14800 -26133
rect 14860 -26193 14870 -26133
rect 14790 -26263 14870 -26193
rect 14790 -26313 14800 -26263
rect 14342 -26625 14402 -26323
rect 14860 -26313 14870 -26263
rect 15246 -26193 15256 -26133
rect 15316 -26193 15326 -26133
rect 15246 -26263 15326 -26193
rect 15246 -26313 15256 -26263
rect 14800 -26625 14860 -26323
rect 15316 -26313 15326 -26263
rect 15256 -26625 15316 -26323
rect 160 -26685 170 -26625
rect 230 -26685 240 -26625
rect 160 -26755 240 -26685
rect 160 -26805 170 -26755
rect 230 -26805 240 -26755
rect 616 -26685 626 -26625
rect 686 -26685 696 -26625
rect 616 -26755 696 -26685
rect 616 -26805 626 -26755
rect 170 -27127 230 -26815
rect 686 -26805 696 -26755
rect 1072 -26685 1082 -26625
rect 1142 -26685 1152 -26625
rect 1072 -26755 1152 -26685
rect 1072 -26805 1082 -26755
rect 626 -27127 686 -26815
rect 1142 -26805 1152 -26755
rect 1530 -26685 1540 -26625
rect 1600 -26685 1610 -26625
rect 1530 -26755 1610 -26685
rect 1530 -26805 1540 -26755
rect 1082 -27127 1142 -26815
rect 1600 -26805 1610 -26755
rect 1986 -26685 1996 -26625
rect 2056 -26685 2066 -26625
rect 1986 -26755 2066 -26685
rect 1986 -26805 1996 -26755
rect 1540 -27127 1600 -26815
rect 2056 -26805 2066 -26755
rect 2442 -26685 2452 -26625
rect 2512 -26685 2522 -26625
rect 2442 -26755 2522 -26685
rect 2442 -26805 2452 -26755
rect 1996 -27127 2056 -26815
rect 2512 -26805 2522 -26755
rect 2900 -26685 2910 -26625
rect 2970 -26685 2980 -26625
rect 2900 -26755 2980 -26685
rect 2900 -26805 2910 -26755
rect 2452 -27127 2512 -26815
rect 2970 -26805 2980 -26755
rect 3356 -26685 3366 -26625
rect 3426 -26685 3436 -26625
rect 3356 -26755 3436 -26685
rect 3356 -26805 3366 -26755
rect 2910 -27127 2970 -26815
rect 3426 -26805 3436 -26755
rect 3812 -26685 3822 -26625
rect 3882 -26685 3892 -26625
rect 3812 -26755 3892 -26685
rect 3812 -26805 3822 -26755
rect 3366 -27127 3426 -26815
rect 3882 -26805 3892 -26755
rect 4270 -26685 4280 -26625
rect 4340 -26685 4350 -26625
rect 4270 -26755 4350 -26685
rect 4270 -26805 4280 -26755
rect 3822 -27127 3882 -26815
rect 4340 -26805 4350 -26755
rect 4726 -26685 4736 -26625
rect 4796 -26685 4806 -26625
rect 4726 -26755 4806 -26685
rect 4726 -26805 4736 -26755
rect 4280 -27127 4340 -26815
rect 4796 -26805 4806 -26755
rect 5182 -26685 5192 -26625
rect 5252 -26685 5262 -26625
rect 5182 -26755 5262 -26685
rect 5182 -26805 5192 -26755
rect 4736 -27127 4796 -26815
rect 5252 -26805 5262 -26755
rect 5640 -26685 5650 -26625
rect 5710 -26685 5720 -26625
rect 5640 -26755 5720 -26685
rect 5640 -26805 5650 -26755
rect 5192 -27127 5252 -26815
rect 5710 -26805 5720 -26755
rect 6096 -26685 6106 -26625
rect 6166 -26685 6176 -26625
rect 6096 -26755 6176 -26685
rect 6096 -26805 6106 -26755
rect 5650 -27127 5710 -26815
rect 6166 -26805 6176 -26755
rect 6552 -26685 6562 -26625
rect 6622 -26685 6632 -26625
rect 6552 -26755 6632 -26685
rect 6552 -26805 6562 -26755
rect 6106 -27127 6166 -26815
rect 6622 -26805 6632 -26755
rect 7010 -26685 7020 -26625
rect 7080 -26685 7090 -26625
rect 7010 -26755 7090 -26685
rect 7010 -26805 7020 -26755
rect 6562 -27127 6622 -26815
rect 7080 -26805 7090 -26755
rect 7466 -26685 7476 -26625
rect 7536 -26685 7546 -26625
rect 7466 -26755 7546 -26685
rect 7466 -26805 7476 -26755
rect 7020 -27127 7080 -26815
rect 7536 -26805 7546 -26755
rect 7922 -26685 7932 -26625
rect 7992 -26685 8002 -26625
rect 7922 -26755 8002 -26685
rect 7922 -26805 7932 -26755
rect 7476 -27127 7536 -26815
rect 7992 -26805 8002 -26755
rect 8396 -26685 8406 -26625
rect 8466 -26685 8476 -26625
rect 8396 -26755 8476 -26685
rect 8396 -26805 8406 -26755
rect 7932 -27127 7992 -26815
rect 8466 -26805 8476 -26755
rect 8852 -26685 8862 -26625
rect 8922 -26685 8932 -26625
rect 8852 -26755 8932 -26685
rect 8852 -26805 8862 -26755
rect 8406 -27127 8466 -26815
rect 8922 -26805 8932 -26755
rect 9310 -26685 9320 -26625
rect 9380 -26685 9390 -26625
rect 9310 -26755 9390 -26685
rect 9310 -26805 9320 -26755
rect 8862 -27127 8922 -26815
rect 9380 -26805 9390 -26755
rect 9766 -26685 9776 -26625
rect 9836 -26685 9846 -26625
rect 9766 -26755 9846 -26685
rect 9766 -26805 9776 -26755
rect 9320 -27127 9380 -26815
rect 9836 -26805 9846 -26755
rect 10222 -26685 10232 -26625
rect 10292 -26685 10302 -26625
rect 10222 -26755 10302 -26685
rect 10222 -26805 10232 -26755
rect 9776 -27127 9836 -26815
rect 10292 -26805 10302 -26755
rect 10680 -26685 10690 -26625
rect 10750 -26685 10760 -26625
rect 10680 -26755 10760 -26685
rect 10680 -26805 10690 -26755
rect 10232 -27127 10292 -26815
rect 10750 -26805 10760 -26755
rect 11136 -26685 11146 -26625
rect 11206 -26685 11216 -26625
rect 11136 -26755 11216 -26685
rect 11136 -26805 11146 -26755
rect 10690 -27127 10750 -26815
rect 11206 -26805 11216 -26755
rect 11592 -26685 11602 -26625
rect 11662 -26685 11672 -26625
rect 11592 -26755 11672 -26685
rect 11592 -26805 11602 -26755
rect 11146 -27127 11206 -26815
rect 11662 -26805 11672 -26755
rect 12050 -26685 12060 -26625
rect 12120 -26685 12130 -26625
rect 12050 -26755 12130 -26685
rect 12050 -26805 12060 -26755
rect 11602 -27127 11662 -26815
rect 12120 -26805 12130 -26755
rect 12506 -26685 12516 -26625
rect 12576 -26685 12586 -26625
rect 12506 -26755 12586 -26685
rect 12506 -26805 12516 -26755
rect 12060 -27127 12120 -26815
rect 12576 -26805 12586 -26755
rect 12962 -26685 12972 -26625
rect 13032 -26685 13042 -26625
rect 12962 -26755 13042 -26685
rect 12962 -26805 12972 -26755
rect 12516 -27127 12576 -26815
rect 13032 -26805 13042 -26755
rect 13420 -26685 13430 -26625
rect 13490 -26685 13500 -26625
rect 13420 -26755 13500 -26685
rect 13420 -26805 13430 -26755
rect 12972 -27127 13032 -26815
rect 13490 -26805 13500 -26755
rect 13876 -26685 13886 -26625
rect 13946 -26685 13956 -26625
rect 13876 -26755 13956 -26685
rect 13876 -26805 13886 -26755
rect 13430 -27127 13490 -26815
rect 13946 -26805 13956 -26755
rect 14332 -26685 14342 -26625
rect 14402 -26685 14412 -26625
rect 14332 -26755 14412 -26685
rect 14332 -26805 14342 -26755
rect 13886 -27127 13946 -26815
rect 14402 -26805 14412 -26755
rect 14790 -26685 14800 -26625
rect 14860 -26685 14870 -26625
rect 14790 -26755 14870 -26685
rect 14790 -26805 14800 -26755
rect 14342 -27127 14402 -26815
rect 14860 -26805 14870 -26755
rect 15246 -26685 15256 -26625
rect 15316 -26685 15326 -26625
rect 15246 -26755 15326 -26685
rect 15246 -26805 15256 -26755
rect 14800 -27127 14860 -26815
rect 15316 -26805 15326 -26755
rect 15256 -27127 15316 -26815
rect 160 -27187 170 -27127
rect 230 -27187 240 -27127
rect 160 -27257 240 -27187
rect 160 -27307 170 -27257
rect 230 -27307 240 -27257
rect 616 -27187 626 -27127
rect 686 -27187 696 -27127
rect 616 -27257 696 -27187
rect 616 -27307 626 -27257
rect 170 -27643 230 -27317
rect 686 -27307 696 -27257
rect 1072 -27187 1082 -27127
rect 1142 -27187 1152 -27127
rect 1072 -27257 1152 -27187
rect 1072 -27307 1082 -27257
rect 626 -27643 686 -27317
rect 1142 -27307 1152 -27257
rect 1530 -27187 1540 -27127
rect 1600 -27187 1610 -27127
rect 1530 -27257 1610 -27187
rect 1530 -27307 1540 -27257
rect 1082 -27643 1142 -27317
rect 1600 -27307 1610 -27257
rect 1986 -27187 1996 -27127
rect 2056 -27187 2066 -27127
rect 1986 -27257 2066 -27187
rect 1986 -27307 1996 -27257
rect 1540 -27643 1600 -27317
rect 2056 -27307 2066 -27257
rect 2442 -27187 2452 -27127
rect 2512 -27187 2522 -27127
rect 2442 -27257 2522 -27187
rect 2442 -27307 2452 -27257
rect 1996 -27643 2056 -27317
rect 2512 -27307 2522 -27257
rect 2900 -27187 2910 -27127
rect 2970 -27187 2980 -27127
rect 2900 -27257 2980 -27187
rect 2900 -27307 2910 -27257
rect 2452 -27643 2512 -27317
rect 2970 -27307 2980 -27257
rect 3356 -27187 3366 -27127
rect 3426 -27187 3436 -27127
rect 3356 -27257 3436 -27187
rect 3356 -27307 3366 -27257
rect 2910 -27643 2970 -27317
rect 3426 -27307 3436 -27257
rect 3812 -27187 3822 -27127
rect 3882 -27187 3892 -27127
rect 3812 -27257 3892 -27187
rect 3812 -27307 3822 -27257
rect 3366 -27643 3426 -27317
rect 3882 -27307 3892 -27257
rect 4270 -27187 4280 -27127
rect 4340 -27187 4350 -27127
rect 4270 -27257 4350 -27187
rect 4270 -27307 4280 -27257
rect 3822 -27643 3882 -27317
rect 4340 -27307 4350 -27257
rect 4726 -27187 4736 -27127
rect 4796 -27187 4806 -27127
rect 4726 -27257 4806 -27187
rect 4726 -27307 4736 -27257
rect 4280 -27643 4340 -27317
rect 4796 -27307 4806 -27257
rect 5182 -27187 5192 -27127
rect 5252 -27187 5262 -27127
rect 5182 -27257 5262 -27187
rect 5182 -27307 5192 -27257
rect 4736 -27643 4796 -27317
rect 5252 -27307 5262 -27257
rect 5640 -27187 5650 -27127
rect 5710 -27187 5720 -27127
rect 5640 -27257 5720 -27187
rect 5640 -27307 5650 -27257
rect 5192 -27643 5252 -27317
rect 5710 -27307 5720 -27257
rect 6096 -27187 6106 -27127
rect 6166 -27187 6176 -27127
rect 6096 -27257 6176 -27187
rect 6096 -27307 6106 -27257
rect 5650 -27643 5710 -27317
rect 6166 -27307 6176 -27257
rect 6552 -27187 6562 -27127
rect 6622 -27187 6632 -27127
rect 6552 -27257 6632 -27187
rect 6552 -27307 6562 -27257
rect 6106 -27643 6166 -27317
rect 6622 -27307 6632 -27257
rect 7010 -27187 7020 -27127
rect 7080 -27187 7090 -27127
rect 7010 -27257 7090 -27187
rect 7010 -27307 7020 -27257
rect 6562 -27643 6622 -27317
rect 7080 -27307 7090 -27257
rect 7466 -27187 7476 -27127
rect 7536 -27187 7546 -27127
rect 7466 -27257 7546 -27187
rect 7466 -27307 7476 -27257
rect 7020 -27643 7080 -27317
rect 7536 -27307 7546 -27257
rect 7922 -27187 7932 -27127
rect 7992 -27187 8002 -27127
rect 7922 -27257 8002 -27187
rect 7922 -27307 7932 -27257
rect 7476 -27643 7536 -27317
rect 7992 -27307 8002 -27257
rect 8396 -27187 8406 -27127
rect 8466 -27187 8476 -27127
rect 8396 -27257 8476 -27187
rect 8396 -27307 8406 -27257
rect 7932 -27643 7992 -27317
rect 8466 -27307 8476 -27257
rect 8852 -27187 8862 -27127
rect 8922 -27187 8932 -27127
rect 8852 -27257 8932 -27187
rect 8852 -27307 8862 -27257
rect 8406 -27643 8466 -27317
rect 8922 -27307 8932 -27257
rect 9310 -27187 9320 -27127
rect 9380 -27187 9390 -27127
rect 9310 -27257 9390 -27187
rect 9310 -27307 9320 -27257
rect 8862 -27643 8922 -27317
rect 9380 -27307 9390 -27257
rect 9766 -27187 9776 -27127
rect 9836 -27187 9846 -27127
rect 9766 -27257 9846 -27187
rect 9766 -27307 9776 -27257
rect 9320 -27643 9380 -27317
rect 9836 -27307 9846 -27257
rect 10222 -27187 10232 -27127
rect 10292 -27187 10302 -27127
rect 10222 -27257 10302 -27187
rect 10222 -27307 10232 -27257
rect 9776 -27643 9836 -27317
rect 10292 -27307 10302 -27257
rect 10680 -27187 10690 -27127
rect 10750 -27187 10760 -27127
rect 10680 -27257 10760 -27187
rect 10680 -27307 10690 -27257
rect 10232 -27643 10292 -27317
rect 10750 -27307 10760 -27257
rect 11136 -27187 11146 -27127
rect 11206 -27187 11216 -27127
rect 11136 -27257 11216 -27187
rect 11136 -27307 11146 -27257
rect 10690 -27643 10750 -27317
rect 11206 -27307 11216 -27257
rect 11592 -27187 11602 -27127
rect 11662 -27187 11672 -27127
rect 11592 -27257 11672 -27187
rect 11592 -27307 11602 -27257
rect 11146 -27643 11206 -27317
rect 11662 -27307 11672 -27257
rect 12050 -27187 12060 -27127
rect 12120 -27187 12130 -27127
rect 12050 -27257 12130 -27187
rect 12050 -27307 12060 -27257
rect 11602 -27643 11662 -27317
rect 12120 -27307 12130 -27257
rect 12506 -27187 12516 -27127
rect 12576 -27187 12586 -27127
rect 12506 -27257 12586 -27187
rect 12506 -27307 12516 -27257
rect 12060 -27643 12120 -27317
rect 12576 -27307 12586 -27257
rect 12962 -27187 12972 -27127
rect 13032 -27187 13042 -27127
rect 12962 -27257 13042 -27187
rect 12962 -27307 12972 -27257
rect 12516 -27643 12576 -27317
rect 13032 -27307 13042 -27257
rect 13420 -27187 13430 -27127
rect 13490 -27187 13500 -27127
rect 13420 -27257 13500 -27187
rect 13420 -27307 13430 -27257
rect 12972 -27643 13032 -27317
rect 13490 -27307 13500 -27257
rect 13876 -27187 13886 -27127
rect 13946 -27187 13956 -27127
rect 13876 -27257 13956 -27187
rect 13876 -27307 13886 -27257
rect 13430 -27643 13490 -27317
rect 13946 -27307 13956 -27257
rect 14332 -27187 14342 -27127
rect 14402 -27187 14412 -27127
rect 14332 -27257 14412 -27187
rect 14332 -27307 14342 -27257
rect 13886 -27643 13946 -27317
rect 14402 -27307 14412 -27257
rect 14790 -27187 14800 -27127
rect 14860 -27187 14870 -27127
rect 14790 -27257 14870 -27187
rect 14790 -27307 14800 -27257
rect 14342 -27643 14402 -27317
rect 14860 -27307 14870 -27257
rect 15246 -27187 15256 -27127
rect 15316 -27187 15326 -27127
rect 15246 -27257 15326 -27187
rect 15246 -27307 15256 -27257
rect 14800 -27643 14860 -27317
rect 15316 -27307 15326 -27257
rect 15256 -27643 15316 -27317
rect 160 -27703 170 -27643
rect 230 -27703 240 -27643
rect 160 -27773 240 -27703
rect 160 -27823 170 -27773
rect 230 -27823 240 -27773
rect 616 -27703 626 -27643
rect 686 -27703 696 -27643
rect 616 -27773 696 -27703
rect 616 -27823 626 -27773
rect 170 -28135 230 -27833
rect 686 -27823 696 -27773
rect 1072 -27703 1082 -27643
rect 1142 -27703 1152 -27643
rect 1072 -27773 1152 -27703
rect 1072 -27823 1082 -27773
rect 626 -28135 686 -27833
rect 1142 -27823 1152 -27773
rect 1530 -27703 1540 -27643
rect 1600 -27703 1610 -27643
rect 1530 -27773 1610 -27703
rect 1530 -27823 1540 -27773
rect 1082 -28135 1142 -27833
rect 1600 -27823 1610 -27773
rect 1986 -27703 1996 -27643
rect 2056 -27703 2066 -27643
rect 1986 -27773 2066 -27703
rect 1986 -27823 1996 -27773
rect 1540 -28135 1600 -27833
rect 2056 -27823 2066 -27773
rect 2442 -27703 2452 -27643
rect 2512 -27703 2522 -27643
rect 2442 -27773 2522 -27703
rect 2442 -27823 2452 -27773
rect 1996 -28135 2056 -27833
rect 2512 -27823 2522 -27773
rect 2900 -27703 2910 -27643
rect 2970 -27703 2980 -27643
rect 2900 -27773 2980 -27703
rect 2900 -27823 2910 -27773
rect 2452 -28135 2512 -27833
rect 2970 -27823 2980 -27773
rect 3356 -27703 3366 -27643
rect 3426 -27703 3436 -27643
rect 3356 -27773 3436 -27703
rect 3356 -27823 3366 -27773
rect 2910 -28135 2970 -27833
rect 3426 -27823 3436 -27773
rect 3812 -27703 3822 -27643
rect 3882 -27703 3892 -27643
rect 3812 -27773 3892 -27703
rect 3812 -27823 3822 -27773
rect 3366 -28135 3426 -27833
rect 3882 -27823 3892 -27773
rect 4270 -27703 4280 -27643
rect 4340 -27703 4350 -27643
rect 4270 -27773 4350 -27703
rect 4270 -27823 4280 -27773
rect 3822 -28135 3882 -27833
rect 4340 -27823 4350 -27773
rect 4726 -27703 4736 -27643
rect 4796 -27703 4806 -27643
rect 4726 -27773 4806 -27703
rect 4726 -27823 4736 -27773
rect 4280 -28135 4340 -27833
rect 4796 -27823 4806 -27773
rect 5182 -27703 5192 -27643
rect 5252 -27703 5262 -27643
rect 5182 -27773 5262 -27703
rect 5182 -27823 5192 -27773
rect 4736 -28135 4796 -27833
rect 5252 -27823 5262 -27773
rect 5640 -27703 5650 -27643
rect 5710 -27703 5720 -27643
rect 5640 -27773 5720 -27703
rect 5640 -27823 5650 -27773
rect 5192 -28135 5252 -27833
rect 5710 -27823 5720 -27773
rect 6096 -27703 6106 -27643
rect 6166 -27703 6176 -27643
rect 6096 -27773 6176 -27703
rect 6096 -27823 6106 -27773
rect 5650 -28135 5710 -27833
rect 6166 -27823 6176 -27773
rect 6552 -27703 6562 -27643
rect 6622 -27703 6632 -27643
rect 6552 -27773 6632 -27703
rect 6552 -27823 6562 -27773
rect 6106 -28135 6166 -27833
rect 6622 -27823 6632 -27773
rect 7010 -27703 7020 -27643
rect 7080 -27703 7090 -27643
rect 7010 -27773 7090 -27703
rect 7010 -27823 7020 -27773
rect 6562 -28135 6622 -27833
rect 7080 -27823 7090 -27773
rect 7466 -27703 7476 -27643
rect 7536 -27703 7546 -27643
rect 7466 -27773 7546 -27703
rect 7466 -27823 7476 -27773
rect 7020 -28135 7080 -27833
rect 7536 -27823 7546 -27773
rect 7922 -27703 7932 -27643
rect 7992 -27703 8002 -27643
rect 7922 -27773 8002 -27703
rect 7922 -27823 7932 -27773
rect 7476 -28135 7536 -27833
rect 7992 -27823 8002 -27773
rect 8396 -27703 8406 -27643
rect 8466 -27703 8476 -27643
rect 8396 -27773 8476 -27703
rect 8396 -27823 8406 -27773
rect 7932 -28135 7992 -27833
rect 8466 -27823 8476 -27773
rect 8852 -27703 8862 -27643
rect 8922 -27703 8932 -27643
rect 8852 -27773 8932 -27703
rect 8852 -27823 8862 -27773
rect 8406 -28135 8466 -27833
rect 8922 -27823 8932 -27773
rect 9310 -27703 9320 -27643
rect 9380 -27703 9390 -27643
rect 9310 -27773 9390 -27703
rect 9310 -27823 9320 -27773
rect 8862 -28135 8922 -27833
rect 9380 -27823 9390 -27773
rect 9766 -27703 9776 -27643
rect 9836 -27703 9846 -27643
rect 9766 -27773 9846 -27703
rect 9766 -27823 9776 -27773
rect 9320 -28135 9380 -27833
rect 9836 -27823 9846 -27773
rect 10222 -27703 10232 -27643
rect 10292 -27703 10302 -27643
rect 10222 -27773 10302 -27703
rect 10222 -27823 10232 -27773
rect 9776 -28135 9836 -27833
rect 10292 -27823 10302 -27773
rect 10680 -27703 10690 -27643
rect 10750 -27703 10760 -27643
rect 10680 -27773 10760 -27703
rect 10680 -27823 10690 -27773
rect 10232 -28135 10292 -27833
rect 10750 -27823 10760 -27773
rect 11136 -27703 11146 -27643
rect 11206 -27703 11216 -27643
rect 11136 -27773 11216 -27703
rect 11136 -27823 11146 -27773
rect 10690 -28135 10750 -27833
rect 11206 -27823 11216 -27773
rect 11592 -27703 11602 -27643
rect 11662 -27703 11672 -27643
rect 11592 -27773 11672 -27703
rect 11592 -27823 11602 -27773
rect 11146 -28135 11206 -27833
rect 11662 -27823 11672 -27773
rect 12050 -27703 12060 -27643
rect 12120 -27703 12130 -27643
rect 12050 -27773 12130 -27703
rect 12050 -27823 12060 -27773
rect 11602 -28135 11662 -27833
rect 12120 -27823 12130 -27773
rect 12506 -27703 12516 -27643
rect 12576 -27703 12586 -27643
rect 12506 -27773 12586 -27703
rect 12506 -27823 12516 -27773
rect 12060 -28135 12120 -27833
rect 12576 -27823 12586 -27773
rect 12962 -27703 12972 -27643
rect 13032 -27703 13042 -27643
rect 12962 -27773 13042 -27703
rect 12962 -27823 12972 -27773
rect 12516 -28135 12576 -27833
rect 13032 -27823 13042 -27773
rect 13420 -27703 13430 -27643
rect 13490 -27703 13500 -27643
rect 13420 -27773 13500 -27703
rect 13420 -27823 13430 -27773
rect 12972 -28135 13032 -27833
rect 13490 -27823 13500 -27773
rect 13876 -27703 13886 -27643
rect 13946 -27703 13956 -27643
rect 13876 -27773 13956 -27703
rect 13876 -27823 13886 -27773
rect 13430 -28135 13490 -27833
rect 13946 -27823 13956 -27773
rect 14332 -27703 14342 -27643
rect 14402 -27703 14412 -27643
rect 14332 -27773 14412 -27703
rect 14332 -27823 14342 -27773
rect 13886 -28135 13946 -27833
rect 14402 -27823 14412 -27773
rect 14790 -27703 14800 -27643
rect 14860 -27703 14870 -27643
rect 14790 -27773 14870 -27703
rect 14790 -27823 14800 -27773
rect 14342 -28135 14402 -27833
rect 14860 -27823 14870 -27773
rect 15246 -27703 15256 -27643
rect 15316 -27703 15326 -27643
rect 15246 -27773 15326 -27703
rect 15246 -27823 15256 -27773
rect 14800 -28135 14860 -27833
rect 15316 -27823 15326 -27773
rect 15256 -28135 15316 -27833
rect 160 -28195 170 -28135
rect 230 -28195 240 -28135
rect 160 -28265 240 -28195
rect 160 -28315 170 -28265
rect 230 -28315 240 -28265
rect 616 -28195 626 -28135
rect 686 -28195 696 -28135
rect 616 -28265 696 -28195
rect 616 -28315 626 -28265
rect 170 -28637 230 -28325
rect 686 -28315 696 -28265
rect 1072 -28195 1082 -28135
rect 1142 -28195 1152 -28135
rect 1072 -28265 1152 -28195
rect 1072 -28315 1082 -28265
rect 626 -28637 686 -28325
rect 1142 -28315 1152 -28265
rect 1530 -28195 1540 -28135
rect 1600 -28195 1610 -28135
rect 1530 -28265 1610 -28195
rect 1530 -28315 1540 -28265
rect 1082 -28637 1142 -28325
rect 1600 -28315 1610 -28265
rect 1986 -28195 1996 -28135
rect 2056 -28195 2066 -28135
rect 1986 -28265 2066 -28195
rect 1986 -28315 1996 -28265
rect 1540 -28637 1600 -28325
rect 2056 -28315 2066 -28265
rect 2442 -28195 2452 -28135
rect 2512 -28195 2522 -28135
rect 2442 -28265 2522 -28195
rect 2442 -28315 2452 -28265
rect 1996 -28637 2056 -28325
rect 2512 -28315 2522 -28265
rect 2900 -28195 2910 -28135
rect 2970 -28195 2980 -28135
rect 2900 -28265 2980 -28195
rect 2900 -28315 2910 -28265
rect 2452 -28637 2512 -28325
rect 2970 -28315 2980 -28265
rect 3356 -28195 3366 -28135
rect 3426 -28195 3436 -28135
rect 3356 -28265 3436 -28195
rect 3356 -28315 3366 -28265
rect 2910 -28637 2970 -28325
rect 3426 -28315 3436 -28265
rect 3812 -28195 3822 -28135
rect 3882 -28195 3892 -28135
rect 3812 -28265 3892 -28195
rect 3812 -28315 3822 -28265
rect 3366 -28637 3426 -28325
rect 3882 -28315 3892 -28265
rect 4270 -28195 4280 -28135
rect 4340 -28195 4350 -28135
rect 4270 -28265 4350 -28195
rect 4270 -28315 4280 -28265
rect 3822 -28637 3882 -28325
rect 4340 -28315 4350 -28265
rect 4726 -28195 4736 -28135
rect 4796 -28195 4806 -28135
rect 4726 -28265 4806 -28195
rect 4726 -28315 4736 -28265
rect 4280 -28637 4340 -28325
rect 4796 -28315 4806 -28265
rect 5182 -28195 5192 -28135
rect 5252 -28195 5262 -28135
rect 5182 -28265 5262 -28195
rect 5182 -28315 5192 -28265
rect 4736 -28637 4796 -28325
rect 5252 -28315 5262 -28265
rect 5640 -28195 5650 -28135
rect 5710 -28195 5720 -28135
rect 5640 -28265 5720 -28195
rect 5640 -28315 5650 -28265
rect 5192 -28637 5252 -28325
rect 5710 -28315 5720 -28265
rect 6096 -28195 6106 -28135
rect 6166 -28195 6176 -28135
rect 6096 -28265 6176 -28195
rect 6096 -28315 6106 -28265
rect 5650 -28637 5710 -28325
rect 6166 -28315 6176 -28265
rect 6552 -28195 6562 -28135
rect 6622 -28195 6632 -28135
rect 6552 -28265 6632 -28195
rect 6552 -28315 6562 -28265
rect 6106 -28637 6166 -28325
rect 6622 -28315 6632 -28265
rect 7010 -28195 7020 -28135
rect 7080 -28195 7090 -28135
rect 7010 -28265 7090 -28195
rect 7010 -28315 7020 -28265
rect 6562 -28637 6622 -28325
rect 7080 -28315 7090 -28265
rect 7466 -28195 7476 -28135
rect 7536 -28195 7546 -28135
rect 7466 -28265 7546 -28195
rect 7466 -28315 7476 -28265
rect 7020 -28637 7080 -28325
rect 7536 -28315 7546 -28265
rect 7922 -28195 7932 -28135
rect 7992 -28195 8002 -28135
rect 7922 -28265 8002 -28195
rect 7922 -28315 7932 -28265
rect 7476 -28637 7536 -28325
rect 7992 -28315 8002 -28265
rect 8396 -28195 8406 -28135
rect 8466 -28195 8476 -28135
rect 8396 -28265 8476 -28195
rect 8396 -28315 8406 -28265
rect 7932 -28637 7992 -28325
rect 8466 -28315 8476 -28265
rect 8852 -28195 8862 -28135
rect 8922 -28195 8932 -28135
rect 8852 -28265 8932 -28195
rect 8852 -28315 8862 -28265
rect 8406 -28637 8466 -28325
rect 8922 -28315 8932 -28265
rect 9310 -28195 9320 -28135
rect 9380 -28195 9390 -28135
rect 9310 -28265 9390 -28195
rect 9310 -28315 9320 -28265
rect 8862 -28637 8922 -28325
rect 9380 -28315 9390 -28265
rect 9766 -28195 9776 -28135
rect 9836 -28195 9846 -28135
rect 9766 -28265 9846 -28195
rect 9766 -28315 9776 -28265
rect 9320 -28637 9380 -28325
rect 9836 -28315 9846 -28265
rect 10222 -28195 10232 -28135
rect 10292 -28195 10302 -28135
rect 10222 -28265 10302 -28195
rect 10222 -28315 10232 -28265
rect 9776 -28637 9836 -28325
rect 10292 -28315 10302 -28265
rect 10680 -28195 10690 -28135
rect 10750 -28195 10760 -28135
rect 10680 -28265 10760 -28195
rect 10680 -28315 10690 -28265
rect 10232 -28637 10292 -28325
rect 10750 -28315 10760 -28265
rect 11136 -28195 11146 -28135
rect 11206 -28195 11216 -28135
rect 11136 -28265 11216 -28195
rect 11136 -28315 11146 -28265
rect 10690 -28637 10750 -28325
rect 11206 -28315 11216 -28265
rect 11592 -28195 11602 -28135
rect 11662 -28195 11672 -28135
rect 11592 -28265 11672 -28195
rect 11592 -28315 11602 -28265
rect 11146 -28637 11206 -28325
rect 11662 -28315 11672 -28265
rect 12050 -28195 12060 -28135
rect 12120 -28195 12130 -28135
rect 12050 -28265 12130 -28195
rect 12050 -28315 12060 -28265
rect 11602 -28637 11662 -28325
rect 12120 -28315 12130 -28265
rect 12506 -28195 12516 -28135
rect 12576 -28195 12586 -28135
rect 12506 -28265 12586 -28195
rect 12506 -28315 12516 -28265
rect 12060 -28637 12120 -28325
rect 12576 -28315 12586 -28265
rect 12962 -28195 12972 -28135
rect 13032 -28195 13042 -28135
rect 12962 -28265 13042 -28195
rect 12962 -28315 12972 -28265
rect 12516 -28637 12576 -28325
rect 13032 -28315 13042 -28265
rect 13420 -28195 13430 -28135
rect 13490 -28195 13500 -28135
rect 13420 -28265 13500 -28195
rect 13420 -28315 13430 -28265
rect 12972 -28637 13032 -28325
rect 13490 -28315 13500 -28265
rect 13876 -28195 13886 -28135
rect 13946 -28195 13956 -28135
rect 13876 -28265 13956 -28195
rect 13876 -28315 13886 -28265
rect 13430 -28637 13490 -28325
rect 13946 -28315 13956 -28265
rect 14332 -28195 14342 -28135
rect 14402 -28195 14412 -28135
rect 14332 -28265 14412 -28195
rect 14332 -28315 14342 -28265
rect 13886 -28637 13946 -28325
rect 14402 -28315 14412 -28265
rect 14790 -28195 14800 -28135
rect 14860 -28195 14870 -28135
rect 14790 -28265 14870 -28195
rect 14790 -28315 14800 -28265
rect 14342 -28637 14402 -28325
rect 14860 -28315 14870 -28265
rect 15246 -28195 15256 -28135
rect 15316 -28195 15326 -28135
rect 15246 -28265 15326 -28195
rect 15246 -28315 15256 -28265
rect 14800 -28637 14860 -28325
rect 15316 -28315 15326 -28265
rect 15256 -28637 15316 -28325
rect 160 -28697 170 -28637
rect 230 -28697 240 -28637
rect 160 -28767 240 -28697
rect 160 -28817 170 -28767
rect 230 -28817 240 -28767
rect 616 -28697 626 -28637
rect 686 -28697 696 -28637
rect 616 -28767 696 -28697
rect 616 -28817 626 -28767
rect 170 -29131 230 -28827
rect 686 -28817 696 -28767
rect 1072 -28697 1082 -28637
rect 1142 -28697 1152 -28637
rect 1072 -28767 1152 -28697
rect 1072 -28817 1082 -28767
rect 626 -29131 686 -28827
rect 1142 -28817 1152 -28767
rect 1530 -28697 1540 -28637
rect 1600 -28697 1610 -28637
rect 1530 -28767 1610 -28697
rect 1530 -28817 1540 -28767
rect 1082 -29131 1142 -28827
rect 1600 -28817 1610 -28767
rect 1986 -28697 1996 -28637
rect 2056 -28697 2066 -28637
rect 1986 -28767 2066 -28697
rect 1986 -28817 1996 -28767
rect 1540 -29131 1600 -28827
rect 2056 -28817 2066 -28767
rect 2442 -28697 2452 -28637
rect 2512 -28697 2522 -28637
rect 2442 -28767 2522 -28697
rect 2442 -28817 2452 -28767
rect 1996 -29131 2056 -28827
rect 2512 -28817 2522 -28767
rect 2900 -28697 2910 -28637
rect 2970 -28697 2980 -28637
rect 2900 -28767 2980 -28697
rect 2900 -28817 2910 -28767
rect 2452 -29131 2512 -28827
rect 2970 -28817 2980 -28767
rect 3356 -28697 3366 -28637
rect 3426 -28697 3436 -28637
rect 3356 -28767 3436 -28697
rect 3356 -28817 3366 -28767
rect 2910 -29131 2970 -28827
rect 3426 -28817 3436 -28767
rect 3812 -28697 3822 -28637
rect 3882 -28697 3892 -28637
rect 3812 -28767 3892 -28697
rect 3812 -28817 3822 -28767
rect 3366 -29131 3426 -28827
rect 3882 -28817 3892 -28767
rect 4270 -28697 4280 -28637
rect 4340 -28697 4350 -28637
rect 4270 -28767 4350 -28697
rect 4270 -28817 4280 -28767
rect 3822 -29131 3882 -28827
rect 4340 -28817 4350 -28767
rect 4726 -28697 4736 -28637
rect 4796 -28697 4806 -28637
rect 4726 -28767 4806 -28697
rect 4726 -28817 4736 -28767
rect 4280 -29131 4340 -28827
rect 4796 -28817 4806 -28767
rect 5182 -28697 5192 -28637
rect 5252 -28697 5262 -28637
rect 5182 -28767 5262 -28697
rect 5182 -28817 5192 -28767
rect 4736 -29131 4796 -28827
rect 5252 -28817 5262 -28767
rect 5640 -28697 5650 -28637
rect 5710 -28697 5720 -28637
rect 5640 -28767 5720 -28697
rect 5640 -28817 5650 -28767
rect 5192 -29131 5252 -28827
rect 5710 -28817 5720 -28767
rect 6096 -28697 6106 -28637
rect 6166 -28697 6176 -28637
rect 6096 -28767 6176 -28697
rect 6096 -28817 6106 -28767
rect 5650 -29131 5710 -28827
rect 6166 -28817 6176 -28767
rect 6552 -28697 6562 -28637
rect 6622 -28697 6632 -28637
rect 6552 -28767 6632 -28697
rect 6552 -28817 6562 -28767
rect 6106 -29131 6166 -28827
rect 6622 -28817 6632 -28767
rect 7010 -28697 7020 -28637
rect 7080 -28697 7090 -28637
rect 7010 -28767 7090 -28697
rect 7010 -28817 7020 -28767
rect 6562 -29131 6622 -28827
rect 7080 -28817 7090 -28767
rect 7466 -28697 7476 -28637
rect 7536 -28697 7546 -28637
rect 7466 -28767 7546 -28697
rect 7466 -28817 7476 -28767
rect 7020 -29131 7080 -28827
rect 7536 -28817 7546 -28767
rect 7922 -28697 7932 -28637
rect 7992 -28697 8002 -28637
rect 7922 -28767 8002 -28697
rect 7922 -28817 7932 -28767
rect 7476 -29131 7536 -28827
rect 7992 -28817 8002 -28767
rect 8396 -28697 8406 -28637
rect 8466 -28697 8476 -28637
rect 8396 -28767 8476 -28697
rect 8396 -28817 8406 -28767
rect 7932 -29131 7992 -28827
rect 8466 -28817 8476 -28767
rect 8852 -28697 8862 -28637
rect 8922 -28697 8932 -28637
rect 8852 -28767 8932 -28697
rect 8852 -28817 8862 -28767
rect 8406 -29131 8466 -28827
rect 8922 -28817 8932 -28767
rect 9310 -28697 9320 -28637
rect 9380 -28697 9390 -28637
rect 9310 -28767 9390 -28697
rect 9310 -28817 9320 -28767
rect 8862 -29131 8922 -28827
rect 9380 -28817 9390 -28767
rect 9766 -28697 9776 -28637
rect 9836 -28697 9846 -28637
rect 9766 -28767 9846 -28697
rect 9766 -28817 9776 -28767
rect 9320 -29131 9380 -28827
rect 9836 -28817 9846 -28767
rect 10222 -28697 10232 -28637
rect 10292 -28697 10302 -28637
rect 10222 -28767 10302 -28697
rect 10222 -28817 10232 -28767
rect 9776 -29131 9836 -28827
rect 10292 -28817 10302 -28767
rect 10680 -28697 10690 -28637
rect 10750 -28697 10760 -28637
rect 10680 -28767 10760 -28697
rect 10680 -28817 10690 -28767
rect 10232 -29131 10292 -28827
rect 10750 -28817 10760 -28767
rect 11136 -28697 11146 -28637
rect 11206 -28697 11216 -28637
rect 11136 -28767 11216 -28697
rect 11136 -28817 11146 -28767
rect 10690 -29131 10750 -28827
rect 11206 -28817 11216 -28767
rect 11592 -28697 11602 -28637
rect 11662 -28697 11672 -28637
rect 11592 -28767 11672 -28697
rect 11592 -28817 11602 -28767
rect 11146 -29131 11206 -28827
rect 11662 -28817 11672 -28767
rect 12050 -28697 12060 -28637
rect 12120 -28697 12130 -28637
rect 12050 -28767 12130 -28697
rect 12050 -28817 12060 -28767
rect 11602 -29131 11662 -28827
rect 12120 -28817 12130 -28767
rect 12506 -28697 12516 -28637
rect 12576 -28697 12586 -28637
rect 12506 -28767 12586 -28697
rect 12506 -28817 12516 -28767
rect 12060 -29131 12120 -28827
rect 12576 -28817 12586 -28767
rect 12962 -28697 12972 -28637
rect 13032 -28697 13042 -28637
rect 12962 -28767 13042 -28697
rect 12962 -28817 12972 -28767
rect 12516 -29131 12576 -28827
rect 13032 -28817 13042 -28767
rect 13420 -28697 13430 -28637
rect 13490 -28697 13500 -28637
rect 13420 -28767 13500 -28697
rect 13420 -28817 13430 -28767
rect 12972 -29131 13032 -28827
rect 13490 -28817 13500 -28767
rect 13876 -28697 13886 -28637
rect 13946 -28697 13956 -28637
rect 13876 -28767 13956 -28697
rect 13876 -28817 13886 -28767
rect 13430 -29131 13490 -28827
rect 13946 -28817 13956 -28767
rect 14332 -28697 14342 -28637
rect 14402 -28697 14412 -28637
rect 14332 -28767 14412 -28697
rect 14332 -28817 14342 -28767
rect 13886 -29131 13946 -28827
rect 14402 -28817 14412 -28767
rect 14790 -28697 14800 -28637
rect 14860 -28697 14870 -28637
rect 14790 -28767 14870 -28697
rect 14790 -28817 14800 -28767
rect 14342 -29131 14402 -28827
rect 14860 -28817 14870 -28767
rect 15246 -28697 15256 -28637
rect 15316 -28697 15326 -28637
rect 15246 -28767 15326 -28697
rect 15246 -28817 15256 -28767
rect 14800 -29131 14860 -28827
rect 15316 -28817 15326 -28767
rect 15256 -29131 15316 -28827
rect 160 -29191 170 -29131
rect 230 -29191 240 -29131
rect 160 -29261 240 -29191
rect 160 -29311 170 -29261
rect 230 -29311 240 -29261
rect 616 -29191 626 -29131
rect 686 -29191 696 -29131
rect 616 -29261 696 -29191
rect 616 -29311 626 -29261
rect 170 -29623 230 -29321
rect 686 -29311 696 -29261
rect 1072 -29191 1082 -29131
rect 1142 -29191 1152 -29131
rect 1072 -29261 1152 -29191
rect 1072 -29311 1082 -29261
rect 626 -29623 686 -29321
rect 1142 -29311 1152 -29261
rect 1530 -29191 1540 -29131
rect 1600 -29191 1610 -29131
rect 1530 -29261 1610 -29191
rect 1530 -29311 1540 -29261
rect 1082 -29623 1142 -29321
rect 1600 -29311 1610 -29261
rect 1986 -29191 1996 -29131
rect 2056 -29191 2066 -29131
rect 1986 -29261 2066 -29191
rect 1986 -29311 1996 -29261
rect 1540 -29623 1600 -29321
rect 2056 -29311 2066 -29261
rect 2442 -29191 2452 -29131
rect 2512 -29191 2522 -29131
rect 2442 -29261 2522 -29191
rect 2442 -29311 2452 -29261
rect 1996 -29623 2056 -29321
rect 2512 -29311 2522 -29261
rect 2900 -29191 2910 -29131
rect 2970 -29191 2980 -29131
rect 2900 -29261 2980 -29191
rect 2900 -29311 2910 -29261
rect 2452 -29623 2512 -29321
rect 2970 -29311 2980 -29261
rect 3356 -29191 3366 -29131
rect 3426 -29191 3436 -29131
rect 3356 -29261 3436 -29191
rect 3356 -29311 3366 -29261
rect 2910 -29623 2970 -29321
rect 3426 -29311 3436 -29261
rect 3812 -29191 3822 -29131
rect 3882 -29191 3892 -29131
rect 3812 -29261 3892 -29191
rect 3812 -29311 3822 -29261
rect 3366 -29623 3426 -29321
rect 3882 -29311 3892 -29261
rect 4270 -29191 4280 -29131
rect 4340 -29191 4350 -29131
rect 4270 -29261 4350 -29191
rect 4270 -29311 4280 -29261
rect 3822 -29623 3882 -29321
rect 4340 -29311 4350 -29261
rect 4726 -29191 4736 -29131
rect 4796 -29191 4806 -29131
rect 4726 -29261 4806 -29191
rect 4726 -29311 4736 -29261
rect 4280 -29623 4340 -29321
rect 4796 -29311 4806 -29261
rect 5182 -29191 5192 -29131
rect 5252 -29191 5262 -29131
rect 5182 -29261 5262 -29191
rect 5182 -29311 5192 -29261
rect 4736 -29623 4796 -29321
rect 5252 -29311 5262 -29261
rect 5640 -29191 5650 -29131
rect 5710 -29191 5720 -29131
rect 5640 -29261 5720 -29191
rect 5640 -29311 5650 -29261
rect 5192 -29623 5252 -29321
rect 5710 -29311 5720 -29261
rect 6096 -29191 6106 -29131
rect 6166 -29191 6176 -29131
rect 6096 -29261 6176 -29191
rect 6096 -29311 6106 -29261
rect 5650 -29623 5710 -29321
rect 6166 -29311 6176 -29261
rect 6552 -29191 6562 -29131
rect 6622 -29191 6632 -29131
rect 6552 -29261 6632 -29191
rect 6552 -29311 6562 -29261
rect 6106 -29623 6166 -29321
rect 6622 -29311 6632 -29261
rect 7010 -29191 7020 -29131
rect 7080 -29191 7090 -29131
rect 7010 -29261 7090 -29191
rect 7010 -29311 7020 -29261
rect 6562 -29623 6622 -29321
rect 7080 -29311 7090 -29261
rect 7466 -29191 7476 -29131
rect 7536 -29191 7546 -29131
rect 7466 -29261 7546 -29191
rect 7466 -29311 7476 -29261
rect 7020 -29623 7080 -29321
rect 7536 -29311 7546 -29261
rect 7922 -29191 7932 -29131
rect 7992 -29191 8002 -29131
rect 7922 -29261 8002 -29191
rect 7922 -29311 7932 -29261
rect 7476 -29623 7536 -29321
rect 7992 -29311 8002 -29261
rect 8396 -29191 8406 -29131
rect 8466 -29191 8476 -29131
rect 8396 -29261 8476 -29191
rect 8396 -29311 8406 -29261
rect 7932 -29623 7992 -29321
rect 8466 -29311 8476 -29261
rect 8852 -29191 8862 -29131
rect 8922 -29191 8932 -29131
rect 8852 -29261 8932 -29191
rect 8852 -29311 8862 -29261
rect 8406 -29623 8466 -29321
rect 8922 -29311 8932 -29261
rect 9310 -29191 9320 -29131
rect 9380 -29191 9390 -29131
rect 9310 -29261 9390 -29191
rect 9310 -29311 9320 -29261
rect 8862 -29623 8922 -29321
rect 9380 -29311 9390 -29261
rect 9766 -29191 9776 -29131
rect 9836 -29191 9846 -29131
rect 9766 -29261 9846 -29191
rect 9766 -29311 9776 -29261
rect 9320 -29623 9380 -29321
rect 9836 -29311 9846 -29261
rect 10222 -29191 10232 -29131
rect 10292 -29191 10302 -29131
rect 10222 -29261 10302 -29191
rect 10222 -29311 10232 -29261
rect 9776 -29623 9836 -29321
rect 10292 -29311 10302 -29261
rect 10680 -29191 10690 -29131
rect 10750 -29191 10760 -29131
rect 10680 -29261 10760 -29191
rect 10680 -29311 10690 -29261
rect 10232 -29623 10292 -29321
rect 10750 -29311 10760 -29261
rect 11136 -29191 11146 -29131
rect 11206 -29191 11216 -29131
rect 11136 -29261 11216 -29191
rect 11136 -29311 11146 -29261
rect 10690 -29623 10750 -29321
rect 11206 -29311 11216 -29261
rect 11592 -29191 11602 -29131
rect 11662 -29191 11672 -29131
rect 11592 -29261 11672 -29191
rect 11592 -29311 11602 -29261
rect 11146 -29623 11206 -29321
rect 11662 -29311 11672 -29261
rect 12050 -29191 12060 -29131
rect 12120 -29191 12130 -29131
rect 12050 -29261 12130 -29191
rect 12050 -29311 12060 -29261
rect 11602 -29623 11662 -29321
rect 12120 -29311 12130 -29261
rect 12506 -29191 12516 -29131
rect 12576 -29191 12586 -29131
rect 12506 -29261 12586 -29191
rect 12506 -29311 12516 -29261
rect 12060 -29623 12120 -29321
rect 12576 -29311 12586 -29261
rect 12962 -29191 12972 -29131
rect 13032 -29191 13042 -29131
rect 12962 -29261 13042 -29191
rect 12962 -29311 12972 -29261
rect 12516 -29623 12576 -29321
rect 13032 -29311 13042 -29261
rect 13420 -29191 13430 -29131
rect 13490 -29191 13500 -29131
rect 13420 -29261 13500 -29191
rect 13420 -29311 13430 -29261
rect 12972 -29623 13032 -29321
rect 13490 -29311 13500 -29261
rect 13876 -29191 13886 -29131
rect 13946 -29191 13956 -29131
rect 13876 -29261 13956 -29191
rect 13876 -29311 13886 -29261
rect 13430 -29623 13490 -29321
rect 13946 -29311 13956 -29261
rect 14332 -29191 14342 -29131
rect 14402 -29191 14412 -29131
rect 14332 -29261 14412 -29191
rect 14332 -29311 14342 -29261
rect 13886 -29623 13946 -29321
rect 14402 -29311 14412 -29261
rect 14790 -29191 14800 -29131
rect 14860 -29191 14870 -29131
rect 14790 -29261 14870 -29191
rect 14790 -29311 14800 -29261
rect 14342 -29623 14402 -29321
rect 14860 -29311 14870 -29261
rect 15246 -29191 15256 -29131
rect 15316 -29191 15326 -29131
rect 15246 -29261 15326 -29191
rect 15246 -29311 15256 -29261
rect 14800 -29623 14860 -29321
rect 15316 -29311 15326 -29261
rect 15256 -29623 15316 -29321
rect 160 -29683 170 -29623
rect 230 -29683 240 -29623
rect 160 -29753 240 -29683
rect 160 -29803 170 -29753
rect 230 -29803 240 -29753
rect 616 -29683 626 -29623
rect 686 -29683 696 -29623
rect 616 -29753 696 -29683
rect 616 -29803 626 -29753
rect 170 -30125 230 -29813
rect 686 -29803 696 -29753
rect 1072 -29683 1082 -29623
rect 1142 -29683 1152 -29623
rect 1072 -29753 1152 -29683
rect 1072 -29803 1082 -29753
rect 626 -30125 686 -29813
rect 1142 -29803 1152 -29753
rect 1530 -29683 1540 -29623
rect 1600 -29683 1610 -29623
rect 1530 -29753 1610 -29683
rect 1530 -29803 1540 -29753
rect 1082 -30125 1142 -29813
rect 1600 -29803 1610 -29753
rect 1986 -29683 1996 -29623
rect 2056 -29683 2066 -29623
rect 1986 -29753 2066 -29683
rect 1986 -29803 1996 -29753
rect 1540 -30125 1600 -29813
rect 2056 -29803 2066 -29753
rect 2442 -29683 2452 -29623
rect 2512 -29683 2522 -29623
rect 2442 -29753 2522 -29683
rect 2442 -29803 2452 -29753
rect 1996 -30125 2056 -29813
rect 2512 -29803 2522 -29753
rect 2900 -29683 2910 -29623
rect 2970 -29683 2980 -29623
rect 2900 -29753 2980 -29683
rect 2900 -29803 2910 -29753
rect 2452 -30125 2512 -29813
rect 2970 -29803 2980 -29753
rect 3356 -29683 3366 -29623
rect 3426 -29683 3436 -29623
rect 3356 -29753 3436 -29683
rect 3356 -29803 3366 -29753
rect 2910 -30125 2970 -29813
rect 3426 -29803 3436 -29753
rect 3812 -29683 3822 -29623
rect 3882 -29683 3892 -29623
rect 3812 -29753 3892 -29683
rect 3812 -29803 3822 -29753
rect 3366 -30125 3426 -29813
rect 3882 -29803 3892 -29753
rect 4270 -29683 4280 -29623
rect 4340 -29683 4350 -29623
rect 4270 -29753 4350 -29683
rect 4270 -29803 4280 -29753
rect 3822 -30125 3882 -29813
rect 4340 -29803 4350 -29753
rect 4726 -29683 4736 -29623
rect 4796 -29683 4806 -29623
rect 4726 -29753 4806 -29683
rect 4726 -29803 4736 -29753
rect 4280 -30125 4340 -29813
rect 4796 -29803 4806 -29753
rect 5182 -29683 5192 -29623
rect 5252 -29683 5262 -29623
rect 5182 -29753 5262 -29683
rect 5182 -29803 5192 -29753
rect 4736 -30125 4796 -29813
rect 5252 -29803 5262 -29753
rect 5640 -29683 5650 -29623
rect 5710 -29683 5720 -29623
rect 5640 -29753 5720 -29683
rect 5640 -29803 5650 -29753
rect 5192 -30125 5252 -29813
rect 5710 -29803 5720 -29753
rect 6096 -29683 6106 -29623
rect 6166 -29683 6176 -29623
rect 6096 -29753 6176 -29683
rect 6096 -29803 6106 -29753
rect 5650 -30125 5710 -29813
rect 6166 -29803 6176 -29753
rect 6552 -29683 6562 -29623
rect 6622 -29683 6632 -29623
rect 6552 -29753 6632 -29683
rect 6552 -29803 6562 -29753
rect 6106 -30125 6166 -29813
rect 6622 -29803 6632 -29753
rect 7010 -29683 7020 -29623
rect 7080 -29683 7090 -29623
rect 7010 -29753 7090 -29683
rect 7010 -29803 7020 -29753
rect 6562 -30125 6622 -29813
rect 7080 -29803 7090 -29753
rect 7466 -29683 7476 -29623
rect 7536 -29683 7546 -29623
rect 7466 -29753 7546 -29683
rect 7466 -29803 7476 -29753
rect 7020 -30125 7080 -29813
rect 7536 -29803 7546 -29753
rect 7922 -29683 7932 -29623
rect 7992 -29683 8002 -29623
rect 7922 -29753 8002 -29683
rect 7922 -29803 7932 -29753
rect 7476 -30125 7536 -29813
rect 7992 -29803 8002 -29753
rect 8396 -29683 8406 -29623
rect 8466 -29683 8476 -29623
rect 8396 -29753 8476 -29683
rect 8396 -29803 8406 -29753
rect 7932 -30125 7992 -29813
rect 8466 -29803 8476 -29753
rect 8852 -29683 8862 -29623
rect 8922 -29683 8932 -29623
rect 8852 -29753 8932 -29683
rect 8852 -29803 8862 -29753
rect 8406 -30125 8466 -29813
rect 8922 -29803 8932 -29753
rect 9310 -29683 9320 -29623
rect 9380 -29683 9390 -29623
rect 9310 -29753 9390 -29683
rect 9310 -29803 9320 -29753
rect 8862 -30125 8922 -29813
rect 9380 -29803 9390 -29753
rect 9766 -29683 9776 -29623
rect 9836 -29683 9846 -29623
rect 9766 -29753 9846 -29683
rect 9766 -29803 9776 -29753
rect 9320 -30125 9380 -29813
rect 9836 -29803 9846 -29753
rect 10222 -29683 10232 -29623
rect 10292 -29683 10302 -29623
rect 10222 -29753 10302 -29683
rect 10222 -29803 10232 -29753
rect 9776 -30125 9836 -29813
rect 10292 -29803 10302 -29753
rect 10680 -29683 10690 -29623
rect 10750 -29683 10760 -29623
rect 10680 -29753 10760 -29683
rect 10680 -29803 10690 -29753
rect 10232 -30125 10292 -29813
rect 10750 -29803 10760 -29753
rect 11136 -29683 11146 -29623
rect 11206 -29683 11216 -29623
rect 11136 -29753 11216 -29683
rect 11136 -29803 11146 -29753
rect 10690 -30125 10750 -29813
rect 11206 -29803 11216 -29753
rect 11592 -29683 11602 -29623
rect 11662 -29683 11672 -29623
rect 11592 -29753 11672 -29683
rect 11592 -29803 11602 -29753
rect 11146 -30125 11206 -29813
rect 11662 -29803 11672 -29753
rect 12050 -29683 12060 -29623
rect 12120 -29683 12130 -29623
rect 12050 -29753 12130 -29683
rect 12050 -29803 12060 -29753
rect 11602 -30125 11662 -29813
rect 12120 -29803 12130 -29753
rect 12506 -29683 12516 -29623
rect 12576 -29683 12586 -29623
rect 12506 -29753 12586 -29683
rect 12506 -29803 12516 -29753
rect 12060 -30125 12120 -29813
rect 12576 -29803 12586 -29753
rect 12962 -29683 12972 -29623
rect 13032 -29683 13042 -29623
rect 12962 -29753 13042 -29683
rect 12962 -29803 12972 -29753
rect 12516 -30125 12576 -29813
rect 13032 -29803 13042 -29753
rect 13420 -29683 13430 -29623
rect 13490 -29683 13500 -29623
rect 13420 -29753 13500 -29683
rect 13420 -29803 13430 -29753
rect 12972 -30125 13032 -29813
rect 13490 -29803 13500 -29753
rect 13876 -29683 13886 -29623
rect 13946 -29683 13956 -29623
rect 13876 -29753 13956 -29683
rect 13876 -29803 13886 -29753
rect 13430 -30125 13490 -29813
rect 13946 -29803 13956 -29753
rect 14332 -29683 14342 -29623
rect 14402 -29683 14412 -29623
rect 14332 -29753 14412 -29683
rect 14332 -29803 14342 -29753
rect 13886 -30125 13946 -29813
rect 14402 -29803 14412 -29753
rect 14790 -29683 14800 -29623
rect 14860 -29683 14870 -29623
rect 14790 -29753 14870 -29683
rect 14790 -29803 14800 -29753
rect 14342 -30125 14402 -29813
rect 14860 -29803 14870 -29753
rect 15246 -29683 15256 -29623
rect 15316 -29683 15326 -29623
rect 15246 -29753 15326 -29683
rect 15246 -29803 15256 -29753
rect 14800 -30125 14860 -29813
rect 15316 -29803 15326 -29753
rect 15256 -30125 15316 -29813
rect 160 -30185 170 -30125
rect 230 -30185 240 -30125
rect 160 -30255 240 -30185
rect 160 -30305 170 -30255
rect 230 -30305 240 -30255
rect 616 -30185 626 -30125
rect 686 -30185 696 -30125
rect 616 -30255 696 -30185
rect 616 -30305 626 -30255
rect 170 -30641 230 -30315
rect 686 -30305 696 -30255
rect 1072 -30185 1082 -30125
rect 1142 -30185 1152 -30125
rect 1072 -30255 1152 -30185
rect 1072 -30305 1082 -30255
rect 626 -30641 686 -30315
rect 1142 -30305 1152 -30255
rect 1530 -30185 1540 -30125
rect 1600 -30185 1610 -30125
rect 1530 -30255 1610 -30185
rect 1530 -30305 1540 -30255
rect 1082 -30641 1142 -30315
rect 1600 -30305 1610 -30255
rect 1986 -30185 1996 -30125
rect 2056 -30185 2066 -30125
rect 1986 -30255 2066 -30185
rect 1986 -30305 1996 -30255
rect 1540 -30641 1600 -30315
rect 2056 -30305 2066 -30255
rect 2442 -30185 2452 -30125
rect 2512 -30185 2522 -30125
rect 2442 -30255 2522 -30185
rect 2442 -30305 2452 -30255
rect 1996 -30641 2056 -30315
rect 2512 -30305 2522 -30255
rect 2900 -30185 2910 -30125
rect 2970 -30185 2980 -30125
rect 2900 -30255 2980 -30185
rect 2900 -30305 2910 -30255
rect 2452 -30641 2512 -30315
rect 2970 -30305 2980 -30255
rect 3356 -30185 3366 -30125
rect 3426 -30185 3436 -30125
rect 3356 -30255 3436 -30185
rect 3356 -30305 3366 -30255
rect 2910 -30641 2970 -30315
rect 3426 -30305 3436 -30255
rect 3812 -30185 3822 -30125
rect 3882 -30185 3892 -30125
rect 3812 -30255 3892 -30185
rect 3812 -30305 3822 -30255
rect 3366 -30641 3426 -30315
rect 3882 -30305 3892 -30255
rect 4270 -30185 4280 -30125
rect 4340 -30185 4350 -30125
rect 4270 -30255 4350 -30185
rect 4270 -30305 4280 -30255
rect 3822 -30641 3882 -30315
rect 4340 -30305 4350 -30255
rect 4726 -30185 4736 -30125
rect 4796 -30185 4806 -30125
rect 4726 -30255 4806 -30185
rect 4726 -30305 4736 -30255
rect 4280 -30641 4340 -30315
rect 4796 -30305 4806 -30255
rect 5182 -30185 5192 -30125
rect 5252 -30185 5262 -30125
rect 5182 -30255 5262 -30185
rect 5182 -30305 5192 -30255
rect 4736 -30641 4796 -30315
rect 5252 -30305 5262 -30255
rect 5640 -30185 5650 -30125
rect 5710 -30185 5720 -30125
rect 5640 -30255 5720 -30185
rect 5640 -30305 5650 -30255
rect 5192 -30641 5252 -30315
rect 5710 -30305 5720 -30255
rect 6096 -30185 6106 -30125
rect 6166 -30185 6176 -30125
rect 6096 -30255 6176 -30185
rect 6096 -30305 6106 -30255
rect 5650 -30641 5710 -30315
rect 6166 -30305 6176 -30255
rect 6552 -30185 6562 -30125
rect 6622 -30185 6632 -30125
rect 6552 -30255 6632 -30185
rect 6552 -30305 6562 -30255
rect 6106 -30641 6166 -30315
rect 6622 -30305 6632 -30255
rect 7010 -30185 7020 -30125
rect 7080 -30185 7090 -30125
rect 7010 -30255 7090 -30185
rect 7010 -30305 7020 -30255
rect 6562 -30641 6622 -30315
rect 7080 -30305 7090 -30255
rect 7466 -30185 7476 -30125
rect 7536 -30185 7546 -30125
rect 7466 -30255 7546 -30185
rect 7466 -30305 7476 -30255
rect 7020 -30641 7080 -30315
rect 7536 -30305 7546 -30255
rect 7922 -30185 7932 -30125
rect 7992 -30185 8002 -30125
rect 7922 -30255 8002 -30185
rect 7922 -30305 7932 -30255
rect 7476 -30641 7536 -30315
rect 7992 -30305 8002 -30255
rect 8396 -30185 8406 -30125
rect 8466 -30185 8476 -30125
rect 8396 -30255 8476 -30185
rect 8396 -30305 8406 -30255
rect 7932 -30641 7992 -30315
rect 8466 -30305 8476 -30255
rect 8852 -30185 8862 -30125
rect 8922 -30185 8932 -30125
rect 8852 -30255 8932 -30185
rect 8852 -30305 8862 -30255
rect 8406 -30641 8466 -30315
rect 8922 -30305 8932 -30255
rect 9310 -30185 9320 -30125
rect 9380 -30185 9390 -30125
rect 9310 -30255 9390 -30185
rect 9310 -30305 9320 -30255
rect 8862 -30641 8922 -30315
rect 9380 -30305 9390 -30255
rect 9766 -30185 9776 -30125
rect 9836 -30185 9846 -30125
rect 9766 -30255 9846 -30185
rect 9766 -30305 9776 -30255
rect 9320 -30641 9380 -30315
rect 9836 -30305 9846 -30255
rect 10222 -30185 10232 -30125
rect 10292 -30185 10302 -30125
rect 10222 -30255 10302 -30185
rect 10222 -30305 10232 -30255
rect 9776 -30641 9836 -30315
rect 10292 -30305 10302 -30255
rect 10680 -30185 10690 -30125
rect 10750 -30185 10760 -30125
rect 10680 -30255 10760 -30185
rect 10680 -30305 10690 -30255
rect 10232 -30641 10292 -30315
rect 10750 -30305 10760 -30255
rect 11136 -30185 11146 -30125
rect 11206 -30185 11216 -30125
rect 11136 -30255 11216 -30185
rect 11136 -30305 11146 -30255
rect 10690 -30641 10750 -30315
rect 11206 -30305 11216 -30255
rect 11592 -30185 11602 -30125
rect 11662 -30185 11672 -30125
rect 11592 -30255 11672 -30185
rect 11592 -30305 11602 -30255
rect 11146 -30641 11206 -30315
rect 11662 -30305 11672 -30255
rect 12050 -30185 12060 -30125
rect 12120 -30185 12130 -30125
rect 12050 -30255 12130 -30185
rect 12050 -30305 12060 -30255
rect 11602 -30641 11662 -30315
rect 12120 -30305 12130 -30255
rect 12506 -30185 12516 -30125
rect 12576 -30185 12586 -30125
rect 12506 -30255 12586 -30185
rect 12506 -30305 12516 -30255
rect 12060 -30641 12120 -30315
rect 12576 -30305 12586 -30255
rect 12962 -30185 12972 -30125
rect 13032 -30185 13042 -30125
rect 12962 -30255 13042 -30185
rect 12962 -30305 12972 -30255
rect 12516 -30641 12576 -30315
rect 13032 -30305 13042 -30255
rect 13420 -30185 13430 -30125
rect 13490 -30185 13500 -30125
rect 13420 -30255 13500 -30185
rect 13420 -30305 13430 -30255
rect 12972 -30641 13032 -30315
rect 13490 -30305 13500 -30255
rect 13876 -30185 13886 -30125
rect 13946 -30185 13956 -30125
rect 13876 -30255 13956 -30185
rect 13876 -30305 13886 -30255
rect 13430 -30641 13490 -30315
rect 13946 -30305 13956 -30255
rect 14332 -30185 14342 -30125
rect 14402 -30185 14412 -30125
rect 14332 -30255 14412 -30185
rect 14332 -30305 14342 -30255
rect 13886 -30641 13946 -30315
rect 14402 -30305 14412 -30255
rect 14790 -30185 14800 -30125
rect 14860 -30185 14870 -30125
rect 14790 -30255 14870 -30185
rect 14790 -30305 14800 -30255
rect 14342 -30641 14402 -30315
rect 14860 -30305 14870 -30255
rect 15246 -30185 15256 -30125
rect 15316 -30185 15326 -30125
rect 15246 -30255 15326 -30185
rect 15246 -30305 15256 -30255
rect 14800 -30641 14860 -30315
rect 15316 -30305 15326 -30255
rect 15256 -30641 15316 -30315
rect 160 -30701 170 -30641
rect 230 -30701 240 -30641
rect 160 -30771 240 -30701
rect 160 -30821 170 -30771
rect 230 -30821 240 -30771
rect 616 -30701 626 -30641
rect 686 -30701 696 -30641
rect 616 -30771 696 -30701
rect 616 -30821 626 -30771
rect 170 -31133 230 -30831
rect 686 -30821 696 -30771
rect 1072 -30701 1082 -30641
rect 1142 -30701 1152 -30641
rect 1072 -30771 1152 -30701
rect 1072 -30821 1082 -30771
rect 626 -31133 686 -30831
rect 1142 -30821 1152 -30771
rect 1530 -30701 1540 -30641
rect 1600 -30701 1610 -30641
rect 1530 -30771 1610 -30701
rect 1530 -30821 1540 -30771
rect 1082 -31133 1142 -30831
rect 1600 -30821 1610 -30771
rect 1986 -30701 1996 -30641
rect 2056 -30701 2066 -30641
rect 1986 -30771 2066 -30701
rect 1986 -30821 1996 -30771
rect 1540 -31133 1600 -30831
rect 2056 -30821 2066 -30771
rect 2442 -30701 2452 -30641
rect 2512 -30701 2522 -30641
rect 2442 -30771 2522 -30701
rect 2442 -30821 2452 -30771
rect 1996 -31133 2056 -30831
rect 2512 -30821 2522 -30771
rect 2900 -30701 2910 -30641
rect 2970 -30701 2980 -30641
rect 2900 -30771 2980 -30701
rect 2900 -30821 2910 -30771
rect 2452 -31133 2512 -30831
rect 2970 -30821 2980 -30771
rect 3356 -30701 3366 -30641
rect 3426 -30701 3436 -30641
rect 3356 -30771 3436 -30701
rect 3356 -30821 3366 -30771
rect 2910 -31133 2970 -30831
rect 3426 -30821 3436 -30771
rect 3812 -30701 3822 -30641
rect 3882 -30701 3892 -30641
rect 3812 -30771 3892 -30701
rect 3812 -30821 3822 -30771
rect 3366 -31133 3426 -30831
rect 3882 -30821 3892 -30771
rect 4270 -30701 4280 -30641
rect 4340 -30701 4350 -30641
rect 4270 -30771 4350 -30701
rect 4270 -30821 4280 -30771
rect 3822 -31133 3882 -30831
rect 4340 -30821 4350 -30771
rect 4726 -30701 4736 -30641
rect 4796 -30701 4806 -30641
rect 4726 -30771 4806 -30701
rect 4726 -30821 4736 -30771
rect 4280 -31133 4340 -30831
rect 4796 -30821 4806 -30771
rect 5182 -30701 5192 -30641
rect 5252 -30701 5262 -30641
rect 5182 -30771 5262 -30701
rect 5182 -30821 5192 -30771
rect 4736 -31133 4796 -30831
rect 5252 -30821 5262 -30771
rect 5640 -30701 5650 -30641
rect 5710 -30701 5720 -30641
rect 5640 -30771 5720 -30701
rect 5640 -30821 5650 -30771
rect 5192 -31133 5252 -30831
rect 5710 -30821 5720 -30771
rect 6096 -30701 6106 -30641
rect 6166 -30701 6176 -30641
rect 6096 -30771 6176 -30701
rect 6096 -30821 6106 -30771
rect 5650 -31133 5710 -30831
rect 6166 -30821 6176 -30771
rect 6552 -30701 6562 -30641
rect 6622 -30701 6632 -30641
rect 6552 -30771 6632 -30701
rect 6552 -30821 6562 -30771
rect 6106 -31133 6166 -30831
rect 6622 -30821 6632 -30771
rect 7010 -30701 7020 -30641
rect 7080 -30701 7090 -30641
rect 7010 -30771 7090 -30701
rect 7010 -30821 7020 -30771
rect 6562 -31133 6622 -30831
rect 7080 -30821 7090 -30771
rect 7466 -30701 7476 -30641
rect 7536 -30701 7546 -30641
rect 7466 -30771 7546 -30701
rect 7466 -30821 7476 -30771
rect 7020 -31133 7080 -30831
rect 7536 -30821 7546 -30771
rect 7922 -30701 7932 -30641
rect 7992 -30701 8002 -30641
rect 7922 -30771 8002 -30701
rect 7922 -30821 7932 -30771
rect 7476 -31133 7536 -30831
rect 7992 -30821 8002 -30771
rect 8396 -30701 8406 -30641
rect 8466 -30701 8476 -30641
rect 8396 -30771 8476 -30701
rect 8396 -30821 8406 -30771
rect 7932 -31133 7992 -30831
rect 8466 -30821 8476 -30771
rect 8852 -30701 8862 -30641
rect 8922 -30701 8932 -30641
rect 8852 -30771 8932 -30701
rect 8852 -30821 8862 -30771
rect 8406 -31133 8466 -30831
rect 8922 -30821 8932 -30771
rect 9310 -30701 9320 -30641
rect 9380 -30701 9390 -30641
rect 9310 -30771 9390 -30701
rect 9310 -30821 9320 -30771
rect 8862 -31133 8922 -30831
rect 9380 -30821 9390 -30771
rect 9766 -30701 9776 -30641
rect 9836 -30701 9846 -30641
rect 9766 -30771 9846 -30701
rect 9766 -30821 9776 -30771
rect 9320 -31133 9380 -30831
rect 9836 -30821 9846 -30771
rect 10222 -30701 10232 -30641
rect 10292 -30701 10302 -30641
rect 10222 -30771 10302 -30701
rect 10222 -30821 10232 -30771
rect 9776 -31133 9836 -30831
rect 10292 -30821 10302 -30771
rect 10680 -30701 10690 -30641
rect 10750 -30701 10760 -30641
rect 10680 -30771 10760 -30701
rect 10680 -30821 10690 -30771
rect 10232 -31133 10292 -30831
rect 10750 -30821 10760 -30771
rect 11136 -30701 11146 -30641
rect 11206 -30701 11216 -30641
rect 11136 -30771 11216 -30701
rect 11136 -30821 11146 -30771
rect 10690 -31133 10750 -30831
rect 11206 -30821 11216 -30771
rect 11592 -30701 11602 -30641
rect 11662 -30701 11672 -30641
rect 11592 -30771 11672 -30701
rect 11592 -30821 11602 -30771
rect 11146 -31133 11206 -30831
rect 11662 -30821 11672 -30771
rect 12050 -30701 12060 -30641
rect 12120 -30701 12130 -30641
rect 12050 -30771 12130 -30701
rect 12050 -30821 12060 -30771
rect 11602 -31133 11662 -30831
rect 12120 -30821 12130 -30771
rect 12506 -30701 12516 -30641
rect 12576 -30701 12586 -30641
rect 12506 -30771 12586 -30701
rect 12506 -30821 12516 -30771
rect 12060 -31133 12120 -30831
rect 12576 -30821 12586 -30771
rect 12962 -30701 12972 -30641
rect 13032 -30701 13042 -30641
rect 12962 -30771 13042 -30701
rect 12962 -30821 12972 -30771
rect 12516 -31133 12576 -30831
rect 13032 -30821 13042 -30771
rect 13420 -30701 13430 -30641
rect 13490 -30701 13500 -30641
rect 13420 -30771 13500 -30701
rect 13420 -30821 13430 -30771
rect 12972 -31133 13032 -30831
rect 13490 -30821 13500 -30771
rect 13876 -30701 13886 -30641
rect 13946 -30701 13956 -30641
rect 13876 -30771 13956 -30701
rect 13876 -30821 13886 -30771
rect 13430 -31133 13490 -30831
rect 13946 -30821 13956 -30771
rect 14332 -30701 14342 -30641
rect 14402 -30701 14412 -30641
rect 14332 -30771 14412 -30701
rect 14332 -30821 14342 -30771
rect 13886 -31133 13946 -30831
rect 14402 -30821 14412 -30771
rect 14790 -30701 14800 -30641
rect 14860 -30701 14870 -30641
rect 14790 -30771 14870 -30701
rect 14790 -30821 14800 -30771
rect 14342 -31133 14402 -30831
rect 14860 -30821 14870 -30771
rect 15246 -30701 15256 -30641
rect 15316 -30701 15326 -30641
rect 15246 -30771 15326 -30701
rect 15246 -30821 15256 -30771
rect 14800 -31133 14860 -30831
rect 15316 -30821 15326 -30771
rect 15256 -31133 15316 -30831
rect 160 -31193 170 -31133
rect 230 -31193 240 -31133
rect 160 -31263 240 -31193
rect 160 -31313 170 -31263
rect 230 -31313 240 -31263
rect 616 -31193 626 -31133
rect 686 -31193 696 -31133
rect 616 -31263 696 -31193
rect 616 -31313 626 -31263
rect 170 -31635 230 -31323
rect 686 -31313 696 -31263
rect 1072 -31193 1082 -31133
rect 1142 -31193 1152 -31133
rect 1072 -31263 1152 -31193
rect 1072 -31313 1082 -31263
rect 626 -31635 686 -31323
rect 1142 -31313 1152 -31263
rect 1530 -31193 1540 -31133
rect 1600 -31193 1610 -31133
rect 1530 -31263 1610 -31193
rect 1530 -31313 1540 -31263
rect 1082 -31635 1142 -31323
rect 1600 -31313 1610 -31263
rect 1986 -31193 1996 -31133
rect 2056 -31193 2066 -31133
rect 1986 -31263 2066 -31193
rect 1986 -31313 1996 -31263
rect 1540 -31635 1600 -31323
rect 2056 -31313 2066 -31263
rect 2442 -31193 2452 -31133
rect 2512 -31193 2522 -31133
rect 2442 -31263 2522 -31193
rect 2442 -31313 2452 -31263
rect 1996 -31635 2056 -31323
rect 2512 -31313 2522 -31263
rect 2900 -31193 2910 -31133
rect 2970 -31193 2980 -31133
rect 2900 -31263 2980 -31193
rect 2900 -31313 2910 -31263
rect 2452 -31635 2512 -31323
rect 2970 -31313 2980 -31263
rect 3356 -31193 3366 -31133
rect 3426 -31193 3436 -31133
rect 3356 -31263 3436 -31193
rect 3356 -31313 3366 -31263
rect 2910 -31635 2970 -31323
rect 3426 -31313 3436 -31263
rect 3812 -31193 3822 -31133
rect 3882 -31193 3892 -31133
rect 3812 -31263 3892 -31193
rect 3812 -31313 3822 -31263
rect 3366 -31635 3426 -31323
rect 3882 -31313 3892 -31263
rect 4270 -31193 4280 -31133
rect 4340 -31193 4350 -31133
rect 4270 -31263 4350 -31193
rect 4270 -31313 4280 -31263
rect 3822 -31635 3882 -31323
rect 4340 -31313 4350 -31263
rect 4726 -31193 4736 -31133
rect 4796 -31193 4806 -31133
rect 4726 -31263 4806 -31193
rect 4726 -31313 4736 -31263
rect 4280 -31635 4340 -31323
rect 4796 -31313 4806 -31263
rect 5182 -31193 5192 -31133
rect 5252 -31193 5262 -31133
rect 5182 -31263 5262 -31193
rect 5182 -31313 5192 -31263
rect 4736 -31635 4796 -31323
rect 5252 -31313 5262 -31263
rect 5640 -31193 5650 -31133
rect 5710 -31193 5720 -31133
rect 5640 -31263 5720 -31193
rect 5640 -31313 5650 -31263
rect 5192 -31635 5252 -31323
rect 5710 -31313 5720 -31263
rect 6096 -31193 6106 -31133
rect 6166 -31193 6176 -31133
rect 6096 -31263 6176 -31193
rect 6096 -31313 6106 -31263
rect 5650 -31635 5710 -31323
rect 6166 -31313 6176 -31263
rect 6552 -31193 6562 -31133
rect 6622 -31193 6632 -31133
rect 6552 -31263 6632 -31193
rect 6552 -31313 6562 -31263
rect 6106 -31635 6166 -31323
rect 6622 -31313 6632 -31263
rect 7010 -31193 7020 -31133
rect 7080 -31193 7090 -31133
rect 7010 -31263 7090 -31193
rect 7010 -31313 7020 -31263
rect 6562 -31635 6622 -31323
rect 7080 -31313 7090 -31263
rect 7466 -31193 7476 -31133
rect 7536 -31193 7546 -31133
rect 7466 -31263 7546 -31193
rect 7466 -31313 7476 -31263
rect 7020 -31635 7080 -31323
rect 7536 -31313 7546 -31263
rect 7922 -31193 7932 -31133
rect 7992 -31193 8002 -31133
rect 7922 -31263 8002 -31193
rect 7922 -31313 7932 -31263
rect 7476 -31635 7536 -31323
rect 7992 -31313 8002 -31263
rect 8396 -31193 8406 -31133
rect 8466 -31193 8476 -31133
rect 8396 -31263 8476 -31193
rect 8396 -31313 8406 -31263
rect 7932 -31635 7992 -31323
rect 8466 -31313 8476 -31263
rect 8852 -31193 8862 -31133
rect 8922 -31193 8932 -31133
rect 8852 -31263 8932 -31193
rect 8852 -31313 8862 -31263
rect 8406 -31635 8466 -31323
rect 8922 -31313 8932 -31263
rect 9310 -31193 9320 -31133
rect 9380 -31193 9390 -31133
rect 9310 -31263 9390 -31193
rect 9310 -31313 9320 -31263
rect 8862 -31635 8922 -31323
rect 9380 -31313 9390 -31263
rect 9766 -31193 9776 -31133
rect 9836 -31193 9846 -31133
rect 9766 -31263 9846 -31193
rect 9766 -31313 9776 -31263
rect 9320 -31635 9380 -31323
rect 9836 -31313 9846 -31263
rect 10222 -31193 10232 -31133
rect 10292 -31193 10302 -31133
rect 10222 -31263 10302 -31193
rect 10222 -31313 10232 -31263
rect 9776 -31635 9836 -31323
rect 10292 -31313 10302 -31263
rect 10680 -31193 10690 -31133
rect 10750 -31193 10760 -31133
rect 10680 -31263 10760 -31193
rect 10680 -31313 10690 -31263
rect 10232 -31635 10292 -31323
rect 10750 -31313 10760 -31263
rect 11136 -31193 11146 -31133
rect 11206 -31193 11216 -31133
rect 11136 -31263 11216 -31193
rect 11136 -31313 11146 -31263
rect 10690 -31635 10750 -31323
rect 11206 -31313 11216 -31263
rect 11592 -31193 11602 -31133
rect 11662 -31193 11672 -31133
rect 11592 -31263 11672 -31193
rect 11592 -31313 11602 -31263
rect 11146 -31635 11206 -31323
rect 11662 -31313 11672 -31263
rect 12050 -31193 12060 -31133
rect 12120 -31193 12130 -31133
rect 12050 -31263 12130 -31193
rect 12050 -31313 12060 -31263
rect 11602 -31635 11662 -31323
rect 12120 -31313 12130 -31263
rect 12506 -31193 12516 -31133
rect 12576 -31193 12586 -31133
rect 12506 -31263 12586 -31193
rect 12506 -31313 12516 -31263
rect 12060 -31635 12120 -31323
rect 12576 -31313 12586 -31263
rect 12962 -31193 12972 -31133
rect 13032 -31193 13042 -31133
rect 12962 -31263 13042 -31193
rect 12962 -31313 12972 -31263
rect 12516 -31635 12576 -31323
rect 13032 -31313 13042 -31263
rect 13420 -31193 13430 -31133
rect 13490 -31193 13500 -31133
rect 13420 -31263 13500 -31193
rect 13420 -31313 13430 -31263
rect 12972 -31635 13032 -31323
rect 13490 -31313 13500 -31263
rect 13876 -31193 13886 -31133
rect 13946 -31193 13956 -31133
rect 13876 -31263 13956 -31193
rect 13876 -31313 13886 -31263
rect 13430 -31635 13490 -31323
rect 13946 -31313 13956 -31263
rect 14332 -31193 14342 -31133
rect 14402 -31193 14412 -31133
rect 14332 -31263 14412 -31193
rect 14332 -31313 14342 -31263
rect 13886 -31635 13946 -31323
rect 14402 -31313 14412 -31263
rect 14790 -31193 14800 -31133
rect 14860 -31193 14870 -31133
rect 14790 -31263 14870 -31193
rect 14790 -31313 14800 -31263
rect 14342 -31635 14402 -31323
rect 14860 -31313 14870 -31263
rect 15246 -31193 15256 -31133
rect 15316 -31193 15326 -31133
rect 15246 -31263 15326 -31193
rect 15246 -31313 15256 -31263
rect 14800 -31635 14860 -31323
rect 15316 -31313 15326 -31263
rect 15256 -31635 15316 -31323
rect 160 -31695 170 -31635
rect 230 -31695 240 -31635
rect 160 -31765 240 -31695
rect 160 -31815 170 -31765
rect 230 -31815 240 -31765
rect 616 -31695 626 -31635
rect 686 -31695 696 -31635
rect 616 -31765 696 -31695
rect 616 -31815 626 -31765
rect 170 -32127 230 -31825
rect 686 -31815 696 -31765
rect 1072 -31695 1082 -31635
rect 1142 -31695 1152 -31635
rect 1072 -31765 1152 -31695
rect 1072 -31815 1082 -31765
rect 626 -32127 686 -31825
rect 1142 -31815 1152 -31765
rect 1530 -31695 1540 -31635
rect 1600 -31695 1610 -31635
rect 1530 -31765 1610 -31695
rect 1530 -31815 1540 -31765
rect 1082 -32127 1142 -31825
rect 1600 -31815 1610 -31765
rect 1986 -31695 1996 -31635
rect 2056 -31695 2066 -31635
rect 1986 -31765 2066 -31695
rect 1986 -31815 1996 -31765
rect 1540 -32127 1600 -31825
rect 2056 -31815 2066 -31765
rect 2442 -31695 2452 -31635
rect 2512 -31695 2522 -31635
rect 2442 -31765 2522 -31695
rect 2442 -31815 2452 -31765
rect 1996 -32127 2056 -31825
rect 2512 -31815 2522 -31765
rect 2900 -31695 2910 -31635
rect 2970 -31695 2980 -31635
rect 2900 -31765 2980 -31695
rect 2900 -31815 2910 -31765
rect 2452 -32127 2512 -31825
rect 2970 -31815 2980 -31765
rect 3356 -31695 3366 -31635
rect 3426 -31695 3436 -31635
rect 3356 -31765 3436 -31695
rect 3356 -31815 3366 -31765
rect 2910 -32127 2970 -31825
rect 3426 -31815 3436 -31765
rect 3812 -31695 3822 -31635
rect 3882 -31695 3892 -31635
rect 3812 -31765 3892 -31695
rect 3812 -31815 3822 -31765
rect 3366 -32127 3426 -31825
rect 3882 -31815 3892 -31765
rect 4270 -31695 4280 -31635
rect 4340 -31695 4350 -31635
rect 4270 -31765 4350 -31695
rect 4270 -31815 4280 -31765
rect 3822 -32127 3882 -31825
rect 4340 -31815 4350 -31765
rect 4726 -31695 4736 -31635
rect 4796 -31695 4806 -31635
rect 4726 -31765 4806 -31695
rect 4726 -31815 4736 -31765
rect 4280 -32127 4340 -31825
rect 4796 -31815 4806 -31765
rect 5182 -31695 5192 -31635
rect 5252 -31695 5262 -31635
rect 5182 -31765 5262 -31695
rect 5182 -31815 5192 -31765
rect 4736 -32127 4796 -31825
rect 5252 -31815 5262 -31765
rect 5640 -31695 5650 -31635
rect 5710 -31695 5720 -31635
rect 5640 -31765 5720 -31695
rect 5640 -31815 5650 -31765
rect 5192 -32127 5252 -31825
rect 5710 -31815 5720 -31765
rect 6096 -31695 6106 -31635
rect 6166 -31695 6176 -31635
rect 6096 -31765 6176 -31695
rect 6096 -31815 6106 -31765
rect 5650 -32127 5710 -31825
rect 6166 -31815 6176 -31765
rect 6552 -31695 6562 -31635
rect 6622 -31695 6632 -31635
rect 6552 -31765 6632 -31695
rect 6552 -31815 6562 -31765
rect 6106 -32127 6166 -31825
rect 6622 -31815 6632 -31765
rect 7010 -31695 7020 -31635
rect 7080 -31695 7090 -31635
rect 7010 -31765 7090 -31695
rect 7010 -31815 7020 -31765
rect 6562 -32127 6622 -31825
rect 7080 -31815 7090 -31765
rect 7466 -31695 7476 -31635
rect 7536 -31695 7546 -31635
rect 7466 -31765 7546 -31695
rect 7466 -31815 7476 -31765
rect 7020 -32127 7080 -31825
rect 7536 -31815 7546 -31765
rect 7922 -31695 7932 -31635
rect 7992 -31695 8002 -31635
rect 7922 -31765 8002 -31695
rect 7922 -31815 7932 -31765
rect 7476 -32127 7536 -31825
rect 7992 -31815 8002 -31765
rect 8396 -31695 8406 -31635
rect 8466 -31695 8476 -31635
rect 8396 -31765 8476 -31695
rect 8396 -31815 8406 -31765
rect 7932 -32127 7992 -31825
rect 8466 -31815 8476 -31765
rect 8852 -31695 8862 -31635
rect 8922 -31695 8932 -31635
rect 8852 -31765 8932 -31695
rect 8852 -31815 8862 -31765
rect 8406 -32127 8466 -31825
rect 8922 -31815 8932 -31765
rect 9310 -31695 9320 -31635
rect 9380 -31695 9390 -31635
rect 9310 -31765 9390 -31695
rect 9310 -31815 9320 -31765
rect 8862 -32127 8922 -31825
rect 9380 -31815 9390 -31765
rect 9766 -31695 9776 -31635
rect 9836 -31695 9846 -31635
rect 9766 -31765 9846 -31695
rect 9766 -31815 9776 -31765
rect 9320 -32127 9380 -31825
rect 9836 -31815 9846 -31765
rect 10222 -31695 10232 -31635
rect 10292 -31695 10302 -31635
rect 10222 -31765 10302 -31695
rect 10222 -31815 10232 -31765
rect 9776 -32127 9836 -31825
rect 10292 -31815 10302 -31765
rect 10680 -31695 10690 -31635
rect 10750 -31695 10760 -31635
rect 10680 -31765 10760 -31695
rect 10680 -31815 10690 -31765
rect 10232 -32127 10292 -31825
rect 10750 -31815 10760 -31765
rect 11136 -31695 11146 -31635
rect 11206 -31695 11216 -31635
rect 11136 -31765 11216 -31695
rect 11136 -31815 11146 -31765
rect 10690 -32127 10750 -31825
rect 11206 -31815 11216 -31765
rect 11592 -31695 11602 -31635
rect 11662 -31695 11672 -31635
rect 11592 -31765 11672 -31695
rect 11592 -31815 11602 -31765
rect 11146 -32127 11206 -31825
rect 11662 -31815 11672 -31765
rect 12050 -31695 12060 -31635
rect 12120 -31695 12130 -31635
rect 12050 -31765 12130 -31695
rect 12050 -31815 12060 -31765
rect 11602 -32127 11662 -31825
rect 12120 -31815 12130 -31765
rect 12506 -31695 12516 -31635
rect 12576 -31695 12586 -31635
rect 12506 -31765 12586 -31695
rect 12506 -31815 12516 -31765
rect 12060 -32127 12120 -31825
rect 12576 -31815 12586 -31765
rect 12962 -31695 12972 -31635
rect 13032 -31695 13042 -31635
rect 12962 -31765 13042 -31695
rect 12962 -31815 12972 -31765
rect 12516 -32127 12576 -31825
rect 13032 -31815 13042 -31765
rect 13420 -31695 13430 -31635
rect 13490 -31695 13500 -31635
rect 13420 -31765 13500 -31695
rect 13420 -31815 13430 -31765
rect 12972 -32127 13032 -31825
rect 13490 -31815 13500 -31765
rect 13876 -31695 13886 -31635
rect 13946 -31695 13956 -31635
rect 13876 -31765 13956 -31695
rect 13876 -31815 13886 -31765
rect 13430 -32127 13490 -31825
rect 13946 -31815 13956 -31765
rect 14332 -31695 14342 -31635
rect 14402 -31695 14412 -31635
rect 14332 -31765 14412 -31695
rect 14332 -31815 14342 -31765
rect 13886 -32127 13946 -31825
rect 14402 -31815 14412 -31765
rect 14790 -31695 14800 -31635
rect 14860 -31695 14870 -31635
rect 14790 -31765 14870 -31695
rect 14790 -31815 14800 -31765
rect 14342 -32127 14402 -31825
rect 14860 -31815 14870 -31765
rect 15246 -31695 15256 -31635
rect 15316 -31695 15326 -31635
rect 15246 -31765 15326 -31695
rect 15246 -31815 15256 -31765
rect 14800 -32127 14860 -31825
rect 15316 -31815 15326 -31765
rect 15256 -32127 15316 -31825
rect 160 -32187 170 -32127
rect 230 -32187 240 -32127
rect 160 -32257 240 -32187
rect 160 -32307 170 -32257
rect 230 -32307 240 -32257
rect 616 -32187 626 -32127
rect 686 -32187 696 -32127
rect 616 -32257 696 -32187
rect 616 -32307 626 -32257
rect 170 -32447 230 -32317
rect 686 -32307 696 -32257
rect 1072 -32187 1082 -32127
rect 1142 -32187 1152 -32127
rect 1072 -32257 1152 -32187
rect 1072 -32307 1082 -32257
rect 626 -32447 686 -32317
rect 1142 -32307 1152 -32257
rect 1530 -32187 1540 -32127
rect 1600 -32187 1610 -32127
rect 1530 -32257 1610 -32187
rect 1530 -32307 1540 -32257
rect 1082 -32447 1142 -32317
rect 1600 -32307 1610 -32257
rect 1986 -32187 1996 -32127
rect 2056 -32187 2066 -32127
rect 1986 -32257 2066 -32187
rect 1986 -32307 1996 -32257
rect 1540 -32447 1600 -32317
rect 2056 -32307 2066 -32257
rect 2442 -32187 2452 -32127
rect 2512 -32187 2522 -32127
rect 2442 -32257 2522 -32187
rect 2442 -32307 2452 -32257
rect 1996 -32447 2056 -32317
rect 2512 -32307 2522 -32257
rect 2900 -32187 2910 -32127
rect 2970 -32187 2980 -32127
rect 2900 -32257 2980 -32187
rect 2900 -32307 2910 -32257
rect 2452 -32447 2512 -32317
rect 2970 -32307 2980 -32257
rect 3356 -32187 3366 -32127
rect 3426 -32187 3436 -32127
rect 3356 -32257 3436 -32187
rect 3356 -32307 3366 -32257
rect 2910 -32447 2970 -32317
rect 3426 -32307 3436 -32257
rect 3812 -32187 3822 -32127
rect 3882 -32187 3892 -32127
rect 3812 -32257 3892 -32187
rect 3812 -32307 3822 -32257
rect 3366 -32447 3426 -32317
rect 3882 -32307 3892 -32257
rect 4270 -32187 4280 -32127
rect 4340 -32187 4350 -32127
rect 4270 -32257 4350 -32187
rect 4270 -32307 4280 -32257
rect 3822 -32447 3882 -32317
rect 4340 -32307 4350 -32257
rect 4726 -32187 4736 -32127
rect 4796 -32187 4806 -32127
rect 4726 -32257 4806 -32187
rect 4726 -32307 4736 -32257
rect 4280 -32447 4340 -32317
rect 4796 -32307 4806 -32257
rect 5182 -32187 5192 -32127
rect 5252 -32187 5262 -32127
rect 5182 -32257 5262 -32187
rect 5182 -32307 5192 -32257
rect 4736 -32447 4796 -32317
rect 5252 -32307 5262 -32257
rect 5640 -32187 5650 -32127
rect 5710 -32187 5720 -32127
rect 5640 -32257 5720 -32187
rect 5640 -32307 5650 -32257
rect 5192 -32447 5252 -32317
rect 5710 -32307 5720 -32257
rect 6096 -32187 6106 -32127
rect 6166 -32187 6176 -32127
rect 6096 -32257 6176 -32187
rect 6096 -32307 6106 -32257
rect 5650 -32447 5710 -32317
rect 6166 -32307 6176 -32257
rect 6552 -32187 6562 -32127
rect 6622 -32187 6632 -32127
rect 6552 -32257 6632 -32187
rect 6552 -32307 6562 -32257
rect 6106 -32447 6166 -32317
rect 6622 -32307 6632 -32257
rect 7010 -32187 7020 -32127
rect 7080 -32187 7090 -32127
rect 7010 -32257 7090 -32187
rect 7010 -32307 7020 -32257
rect 6562 -32447 6622 -32317
rect 7080 -32307 7090 -32257
rect 7466 -32187 7476 -32127
rect 7536 -32187 7546 -32127
rect 7466 -32257 7546 -32187
rect 7466 -32307 7476 -32257
rect 7020 -32447 7080 -32317
rect 7536 -32307 7546 -32257
rect 7922 -32187 7932 -32127
rect 7992 -32187 8002 -32127
rect 7922 -32257 8002 -32187
rect 7922 -32307 7932 -32257
rect 7476 -32447 7536 -32317
rect 7992 -32307 8002 -32257
rect 8396 -32187 8406 -32127
rect 8466 -32187 8476 -32127
rect 8396 -32257 8476 -32187
rect 8396 -32307 8406 -32257
rect 7932 -32447 7992 -32317
rect 8466 -32307 8476 -32257
rect 8852 -32187 8862 -32127
rect 8922 -32187 8932 -32127
rect 8852 -32257 8932 -32187
rect 8852 -32307 8862 -32257
rect 8406 -32447 8466 -32317
rect 8922 -32307 8932 -32257
rect 9310 -32187 9320 -32127
rect 9380 -32187 9390 -32127
rect 9310 -32257 9390 -32187
rect 9310 -32307 9320 -32257
rect 8862 -32447 8922 -32317
rect 9380 -32307 9390 -32257
rect 9766 -32187 9776 -32127
rect 9836 -32187 9846 -32127
rect 9766 -32257 9846 -32187
rect 9766 -32307 9776 -32257
rect 9320 -32447 9380 -32317
rect 9836 -32307 9846 -32257
rect 10222 -32187 10232 -32127
rect 10292 -32187 10302 -32127
rect 10222 -32257 10302 -32187
rect 10222 -32307 10232 -32257
rect 9776 -32447 9836 -32317
rect 10292 -32307 10302 -32257
rect 10680 -32187 10690 -32127
rect 10750 -32187 10760 -32127
rect 10680 -32257 10760 -32187
rect 10680 -32307 10690 -32257
rect 10232 -32447 10292 -32317
rect 10750 -32307 10760 -32257
rect 11136 -32187 11146 -32127
rect 11206 -32187 11216 -32127
rect 11136 -32257 11216 -32187
rect 11136 -32307 11146 -32257
rect 10690 -32447 10750 -32317
rect 11206 -32307 11216 -32257
rect 11592 -32187 11602 -32127
rect 11662 -32187 11672 -32127
rect 11592 -32257 11672 -32187
rect 11592 -32307 11602 -32257
rect 11146 -32447 11206 -32317
rect 11662 -32307 11672 -32257
rect 12050 -32187 12060 -32127
rect 12120 -32187 12130 -32127
rect 12050 -32257 12130 -32187
rect 12050 -32307 12060 -32257
rect 11602 -32447 11662 -32317
rect 12120 -32307 12130 -32257
rect 12506 -32187 12516 -32127
rect 12576 -32187 12586 -32127
rect 12506 -32257 12586 -32187
rect 12506 -32307 12516 -32257
rect 12060 -32447 12120 -32317
rect 12576 -32307 12586 -32257
rect 12962 -32187 12972 -32127
rect 13032 -32187 13042 -32127
rect 12962 -32257 13042 -32187
rect 12962 -32307 12972 -32257
rect 12516 -32447 12576 -32317
rect 13032 -32307 13042 -32257
rect 13420 -32187 13430 -32127
rect 13490 -32187 13500 -32127
rect 13420 -32257 13500 -32187
rect 13420 -32307 13430 -32257
rect 12972 -32447 13032 -32317
rect 13490 -32307 13500 -32257
rect 13876 -32187 13886 -32127
rect 13946 -32187 13956 -32127
rect 13876 -32257 13956 -32187
rect 13876 -32307 13886 -32257
rect 13430 -32447 13490 -32317
rect 13946 -32307 13956 -32257
rect 14332 -32187 14342 -32127
rect 14402 -32187 14412 -32127
rect 14332 -32257 14412 -32187
rect 14332 -32307 14342 -32257
rect 13886 -32447 13946 -32317
rect 14402 -32307 14412 -32257
rect 14790 -32187 14800 -32127
rect 14860 -32187 14870 -32127
rect 14790 -32257 14870 -32187
rect 14790 -32307 14800 -32257
rect 14342 -32447 14402 -32317
rect 14860 -32307 14870 -32257
rect 15246 -32187 15256 -32127
rect 15316 -32187 15326 -32127
rect 15246 -32257 15326 -32187
rect 15246 -32307 15256 -32257
rect 14800 -32447 14860 -32317
rect 15316 -32307 15326 -32257
rect 15256 -32447 15316 -32317
<< via4 >>
rect 15127 612 15200 622
rect 15127 611 15201 612
rect 15127 551 15201 611
rect 15357 611 15430 621
rect 15357 551 15358 611
rect 15358 551 15430 611
rect 15357 550 15430 551
rect 614 270 699 348
rect 1066 271 1154 350
rect 1527 330 1612 350
rect 1527 270 1540 330
rect 1540 270 1600 330
rect 1600 270 1612 330
rect 1982 330 2067 350
rect 1982 270 1996 330
rect 1996 270 2056 330
rect 2056 270 2067 330
rect 2438 330 2523 350
rect 2438 270 2452 330
rect 2452 270 2512 330
rect 2512 270 2523 330
rect 2897 330 2982 350
rect 2897 270 2910 330
rect 2910 270 2970 330
rect 2970 270 2982 330
rect 3355 330 3440 350
rect 3355 270 3366 330
rect 3366 270 3426 330
rect 3426 270 3440 330
rect 3807 330 3892 350
rect 3807 270 3822 330
rect 3822 270 3882 330
rect 3882 270 3892 330
rect 4267 330 4352 350
rect 4267 270 4280 330
rect 4280 270 4340 330
rect 4340 270 4352 330
rect 4721 330 4806 350
rect 4721 270 4736 330
rect 4736 270 4796 330
rect 4796 270 4806 330
rect 5180 330 5265 350
rect 5180 270 5192 330
rect 5192 270 5252 330
rect 5252 270 5265 330
rect 5636 330 5721 350
rect 5636 270 5650 330
rect 5650 270 5710 330
rect 5710 270 5721 330
rect 6094 330 6179 350
rect 6094 270 6106 330
rect 6106 270 6166 330
rect 6166 270 6179 330
rect 6548 330 6633 350
rect 6548 270 6562 330
rect 6562 270 6622 330
rect 6622 270 6633 330
rect 7008 330 7093 350
rect 7008 270 7020 330
rect 7020 270 7080 330
rect 7080 270 7093 330
rect 7464 330 7549 350
rect 7464 270 7476 330
rect 7476 270 7536 330
rect 7536 270 7549 330
rect 7917 330 8002 350
rect 7917 270 7932 330
rect 7932 270 7992 330
rect 7992 270 8002 330
rect 8394 330 8479 350
rect 8394 270 8406 330
rect 8406 270 8466 330
rect 8466 270 8479 330
rect 8848 330 8933 350
rect 8848 270 8862 330
rect 8862 270 8922 330
rect 8922 270 8933 330
rect 9306 330 9391 350
rect 9306 270 9320 330
rect 9320 270 9380 330
rect 9380 270 9391 330
rect 9763 330 9848 350
rect 9763 270 9776 330
rect 9776 270 9836 330
rect 9836 270 9848 330
rect 10219 330 10304 350
rect 10219 270 10232 330
rect 10232 270 10292 330
rect 10292 270 10304 330
rect 10678 330 10763 350
rect 10678 270 10690 330
rect 10690 270 10750 330
rect 10750 270 10763 330
rect 11134 330 11219 350
rect 11134 270 11146 330
rect 11146 270 11206 330
rect 11206 270 11219 330
rect 11588 330 11673 350
rect 11588 270 11602 330
rect 11602 270 11662 330
rect 11662 270 11673 330
rect 12048 330 12133 350
rect 12048 270 12060 330
rect 12060 270 12120 330
rect 12120 270 12133 330
rect 12505 330 12590 350
rect 12505 270 12516 330
rect 12516 270 12576 330
rect 12576 270 12590 330
rect 12959 330 13044 350
rect 12959 270 12972 330
rect 12972 270 13032 330
rect 13032 270 13044 330
rect 13419 330 13504 350
rect 13419 270 13430 330
rect 13430 270 13490 330
rect 13490 270 13504 330
rect 13872 330 13957 350
rect 13872 270 13886 330
rect 13886 270 13946 330
rect 13946 270 13957 330
rect 14330 330 14415 350
rect 14330 270 14342 330
rect 14342 270 14402 330
rect 14402 270 14415 330
rect 14790 330 14875 350
rect 14790 270 14800 330
rect 14800 270 14860 330
rect 14860 270 14875 330
<< metal5 >>
rect 15098 622 15461 637
rect 13399 620 13520 621
rect 599 530 14889 620
rect 15098 551 15127 622
rect 15200 621 15461 622
rect 15200 612 15357 621
rect 15201 551 15357 612
rect 15098 550 15357 551
rect 15430 550 15461 621
rect 15098 530 15461 550
rect 600 348 720 530
rect 600 270 614 348
rect 699 270 720 348
rect 600 261 720 270
rect 1050 529 14889 530
rect 1050 350 1170 529
rect 1050 271 1066 350
rect 1154 271 1170 350
rect 1050 262 1170 271
rect 1509 350 1630 529
rect 1509 270 1527 350
rect 1612 270 1630 350
rect 1509 261 1630 270
rect 1967 350 2088 529
rect 1967 270 1982 350
rect 2067 270 2088 350
rect 1967 261 2088 270
rect 2422 350 2543 529
rect 2422 270 2438 350
rect 2523 270 2543 350
rect 2422 261 2543 270
rect 2882 350 3003 529
rect 2882 270 2897 350
rect 2982 270 3003 350
rect 2882 261 3003 270
rect 3339 350 3460 529
rect 3339 270 3355 350
rect 3440 270 3460 350
rect 3339 261 3460 270
rect 3789 350 3910 529
rect 3789 270 3807 350
rect 3892 270 3910 350
rect 3789 261 3910 270
rect 4249 350 4370 529
rect 4249 270 4267 350
rect 4352 270 4370 350
rect 4249 261 4370 270
rect 4702 350 4823 529
rect 4702 270 4721 350
rect 4806 270 4823 350
rect 4702 261 4823 270
rect 5161 350 5282 529
rect 5161 270 5180 350
rect 5265 270 5282 350
rect 5161 261 5282 270
rect 5618 350 5739 529
rect 5618 270 5636 350
rect 5721 270 5739 350
rect 5618 261 5739 270
rect 6078 350 6199 529
rect 6078 270 6094 350
rect 6179 270 6199 350
rect 6078 261 6199 270
rect 6532 350 6653 529
rect 6532 270 6548 350
rect 6633 270 6653 350
rect 6532 261 6653 270
rect 6989 350 7110 529
rect 6989 270 7008 350
rect 7093 270 7110 350
rect 6989 261 7110 270
rect 7444 350 7565 529
rect 7444 270 7464 350
rect 7549 270 7565 350
rect 7444 261 7565 270
rect 7894 350 8015 529
rect 7894 270 7917 350
rect 8002 270 8015 350
rect 7894 261 8015 270
rect 8379 350 8500 529
rect 8379 270 8394 350
rect 8479 270 8500 350
rect 8379 261 8500 270
rect 8830 350 8951 529
rect 8830 270 8848 350
rect 8933 270 8951 350
rect 8830 261 8951 270
rect 9289 350 9410 529
rect 9289 270 9306 350
rect 9391 270 9410 350
rect 9289 261 9410 270
rect 9742 350 9863 529
rect 9742 270 9763 350
rect 9848 270 9863 350
rect 9742 261 9863 270
rect 10199 350 10320 529
rect 10199 270 10219 350
rect 10304 270 10320 350
rect 10199 261 10320 270
rect 10660 350 10781 529
rect 10660 270 10678 350
rect 10763 270 10781 350
rect 10660 261 10781 270
rect 11116 350 11237 529
rect 11116 270 11134 350
rect 11219 270 11237 350
rect 11116 261 11237 270
rect 11570 350 11691 529
rect 11570 270 11588 350
rect 11673 270 11691 350
rect 11570 261 11691 270
rect 12030 350 12151 529
rect 12030 270 12048 350
rect 12133 270 12151 350
rect 12030 261 12151 270
rect 12486 350 12607 529
rect 12486 270 12505 350
rect 12590 270 12607 350
rect 12486 261 12607 270
rect 12943 350 13064 529
rect 12943 270 12959 350
rect 13044 270 13064 350
rect 12943 261 13064 270
rect 13399 350 13520 529
rect 13399 270 13419 350
rect 13504 270 13520 350
rect 13399 262 13520 270
rect 13855 350 13976 529
rect 13855 270 13872 350
rect 13957 270 13976 350
rect 13855 261 13976 270
rect 14310 350 14431 529
rect 14310 270 14330 350
rect 14415 270 14431 350
rect 14310 261 14431 270
rect 14768 350 14889 529
rect 14768 270 14790 350
rect 14875 270 14889 350
rect 14768 261 14889 270
use unit_Cap  unit_Cap_0
timestamp 1756801411
transform 1 0 0 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_1
timestamp 1756801411
transform 1 0 456 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_2
timestamp 1756801411
transform 1 0 912 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_3
timestamp 1756801411
transform 1 0 2282 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_4
timestamp 1756801411
transform 1 0 1826 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_5
timestamp 1756801411
transform 1 0 1370 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_6
timestamp 1756801411
transform 1 0 4110 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_7
timestamp 1756801411
transform 1 0 4566 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_8
timestamp 1756801411
transform 1 0 5022 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_9
timestamp 1756801411
transform 1 0 3652 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_10
timestamp 1756801411
transform 1 0 3196 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_11
timestamp 1756801411
transform 1 0 2740 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_12
timestamp 1756801411
transform 1 0 6850 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_13
timestamp 1756801411
transform 1 0 7306 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_14
timestamp 1756801411
transform 1 0 7762 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_15
timestamp 1756801411
transform 1 0 6392 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_16
timestamp 1756801411
transform 1 0 5936 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_17
timestamp 1756801411
transform 1 0 5480 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_18
timestamp 1756801411
transform 1 0 15086 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_19
timestamp 1756801411
transform 1 0 15086 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_20
timestamp 1756801411
transform 1 0 14630 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_21
timestamp 1756801411
transform 1 0 14172 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_22
timestamp 1756801411
transform 1 0 13716 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_23
timestamp 1756801411
transform 1 0 13260 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_24
timestamp 1756801411
transform 1 0 12802 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_25
timestamp 1756801411
transform 1 0 12346 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_26
timestamp 1756801411
transform 1 0 11890 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_27
timestamp 1756801411
transform 1 0 11432 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_28
timestamp 1756801411
transform 1 0 10976 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_29
timestamp 1756801411
transform 1 0 10520 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_30
timestamp 1756801411
transform 1 0 10062 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_31
timestamp 1756801411
transform 1 0 9606 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_32
timestamp 1756801411
transform 1 0 9150 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_33
timestamp 1756801411
transform 1 0 8692 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_34
timestamp 1756801411
transform 1 0 8236 0 1 20
box 0 -20 400 440
use unit_Cap  unit_Cap_35
timestamp 1756801411
transform 1 0 14630 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_36
timestamp 1756801411
transform 1 0 14172 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_37
timestamp 1756801411
transform 1 0 13716 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_38
timestamp 1756801411
transform 1 0 13260 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_39
timestamp 1756801411
transform 1 0 12802 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_40
timestamp 1756801411
transform 1 0 12346 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_41
timestamp 1756801411
transform 1 0 11890 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_42
timestamp 1756801411
transform 1 0 11432 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_43
timestamp 1756801411
transform 1 0 10976 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_44
timestamp 1756801411
transform 1 0 10520 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_45
timestamp 1756801411
transform 1 0 10062 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_46
timestamp 1756801411
transform 1 0 9606 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_47
timestamp 1756801411
transform 1 0 9150 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_48
timestamp 1756801411
transform 1 0 8692 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_49
timestamp 1756801411
transform 1 0 8236 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_50
timestamp 1756801411
transform 1 0 7762 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_51
timestamp 1756801411
transform 1 0 7306 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_52
timestamp 1756801411
transform 1 0 6850 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_53
timestamp 1756801411
transform 1 0 6392 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_54
timestamp 1756801411
transform 1 0 5936 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_55
timestamp 1756801411
transform 1 0 5480 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_56
timestamp 1756801411
transform 1 0 5022 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_57
timestamp 1756801411
transform 1 0 4110 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_58
timestamp 1756801411
transform 1 0 4566 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_59
timestamp 1756801411
transform 1 0 3196 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_60
timestamp 1756801411
transform 1 0 3652 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_61
timestamp 1756801411
transform 1 0 2282 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_62
timestamp 1756801411
transform 1 0 2740 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_63
timestamp 1756801411
transform 1 0 1370 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_64
timestamp 1756801411
transform 1 0 1826 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_65
timestamp 1756801411
transform 1 0 456 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_66
timestamp 1756801411
transform 1 0 912 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_67
timestamp 1756801411
transform 1 0 0 0 1 -472
box 0 -20 400 440
use unit_Cap  unit_Cap_68
timestamp 1756801411
transform 1 0 14630 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_69
timestamp 1756801411
transform 1 0 15086 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_70
timestamp 1756801411
transform 1 0 13716 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_71
timestamp 1756801411
transform 1 0 14172 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_72
timestamp 1756801411
transform 1 0 12802 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_73
timestamp 1756801411
transform 1 0 13260 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_74
timestamp 1756801411
transform 1 0 11890 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_75
timestamp 1756801411
transform 1 0 12346 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_76
timestamp 1756801411
transform 1 0 10976 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_77
timestamp 1756801411
transform 1 0 11432 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_78
timestamp 1756801411
transform 1 0 10062 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_79
timestamp 1756801411
transform 1 0 10520 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_80
timestamp 1756801411
transform 1 0 9150 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_81
timestamp 1756801411
transform 1 0 9606 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_82
timestamp 1756801411
transform 1 0 8236 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_83
timestamp 1756801411
transform 1 0 8692 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_84
timestamp 1756801411
transform 1 0 7306 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_85
timestamp 1756801411
transform 1 0 7762 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_86
timestamp 1756801411
transform 1 0 6392 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_87
timestamp 1756801411
transform 1 0 6850 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_88
timestamp 1756801411
transform 1 0 5480 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_89
timestamp 1756801411
transform 1 0 5936 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_90
timestamp 1756801411
transform 1 0 4566 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_91
timestamp 1756801411
transform 1 0 5022 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_92
timestamp 1756801411
transform 1 0 3652 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_93
timestamp 1756801411
transform 1 0 4110 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_94
timestamp 1756801411
transform 1 0 2740 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_95
timestamp 1756801411
transform 1 0 3196 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_96
timestamp 1756801411
transform 1 0 1826 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_97
timestamp 1756801411
transform 1 0 2282 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_98
timestamp 1756801411
transform 1 0 912 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_99
timestamp 1756801411
transform 1 0 1370 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_100
timestamp 1756801411
transform 1 0 0 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_101
timestamp 1756801411
transform 1 0 456 0 1 -974
box 0 -20 400 440
use unit_Cap  unit_Cap_102
timestamp 1756801411
transform 1 0 14630 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_103
timestamp 1756801411
transform 1 0 15086 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_104
timestamp 1756801411
transform 1 0 13716 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_105
timestamp 1756801411
transform 1 0 14172 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_106
timestamp 1756801411
transform 1 0 12802 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_107
timestamp 1756801411
transform 1 0 13260 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_108
timestamp 1756801411
transform 1 0 11890 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_109
timestamp 1756801411
transform 1 0 12346 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_110
timestamp 1756801411
transform 1 0 10976 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_111
timestamp 1756801411
transform 1 0 11432 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_112
timestamp 1756801411
transform 1 0 10062 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_113
timestamp 1756801411
transform 1 0 10520 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_114
timestamp 1756801411
transform 1 0 9150 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_115
timestamp 1756801411
transform 1 0 9606 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_116
timestamp 1756801411
transform 1 0 8236 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_117
timestamp 1756801411
transform 1 0 8692 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_118
timestamp 1756801411
transform 1 0 7306 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_119
timestamp 1756801411
transform 1 0 7762 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_120
timestamp 1756801411
transform 1 0 6392 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_121
timestamp 1756801411
transform 1 0 6850 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_122
timestamp 1756801411
transform 1 0 5480 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_123
timestamp 1756801411
transform 1 0 5936 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_124
timestamp 1756801411
transform 1 0 4566 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_125
timestamp 1756801411
transform 1 0 5022 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_126
timestamp 1756801411
transform 1 0 3652 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_127
timestamp 1756801411
transform 1 0 4110 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_128
timestamp 1756801411
transform 1 0 2740 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_129
timestamp 1756801411
transform 1 0 3196 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_130
timestamp 1756801411
transform 1 0 1826 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_131
timestamp 1756801411
transform 1 0 2282 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_132
timestamp 1756801411
transform 1 0 912 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_133
timestamp 1756801411
transform 1 0 1370 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_134
timestamp 1756801411
transform 1 0 0 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_135
timestamp 1756801411
transform 1 0 456 0 1 -1466
box 0 -20 400 440
use unit_Cap  unit_Cap_136
timestamp 1756801411
transform 1 0 15086 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_137
timestamp 1756801411
transform 1 0 15086 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_138
timestamp 1756801411
transform 1 0 14172 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_139
timestamp 1756801411
transform 1 0 14630 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_140
timestamp 1756801411
transform 1 0 14630 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_141
timestamp 1756801411
transform 1 0 14172 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_142
timestamp 1756801411
transform 1 0 13260 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_143
timestamp 1756801411
transform 1 0 13716 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_144
timestamp 1756801411
transform 1 0 13716 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_145
timestamp 1756801411
transform 1 0 13260 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_146
timestamp 1756801411
transform 1 0 12346 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_147
timestamp 1756801411
transform 1 0 12802 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_148
timestamp 1756801411
transform 1 0 12802 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_149
timestamp 1756801411
transform 1 0 12346 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_150
timestamp 1756801411
transform 1 0 11432 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_151
timestamp 1756801411
transform 1 0 11890 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_152
timestamp 1756801411
transform 1 0 11890 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_153
timestamp 1756801411
transform 1 0 11432 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_154
timestamp 1756801411
transform 1 0 10520 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_155
timestamp 1756801411
transform 1 0 10976 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_156
timestamp 1756801411
transform 1 0 10976 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_157
timestamp 1756801411
transform 1 0 10520 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_158
timestamp 1756801411
transform 1 0 9606 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_159
timestamp 1756801411
transform 1 0 10062 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_160
timestamp 1756801411
transform 1 0 10062 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_161
timestamp 1756801411
transform 1 0 9606 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_162
timestamp 1756801411
transform 1 0 8236 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_163
timestamp 1756801411
transform 1 0 8692 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_164
timestamp 1756801411
transform 1 0 9150 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_165
timestamp 1756801411
transform 1 0 9150 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_166
timestamp 1756801411
transform 1 0 8692 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_167
timestamp 1756801411
transform 1 0 8236 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_168
timestamp 1756801411
transform 1 0 7306 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_169
timestamp 1756801411
transform 1 0 7762 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_170
timestamp 1756801411
transform 1 0 7762 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_171
timestamp 1756801411
transform 1 0 7306 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_172
timestamp 1756801411
transform 1 0 6392 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_173
timestamp 1756801411
transform 1 0 6850 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_174
timestamp 1756801411
transform 1 0 6850 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_175
timestamp 1756801411
transform 1 0 6392 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_176
timestamp 1756801411
transform 1 0 5480 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_177
timestamp 1756801411
transform 1 0 5936 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_178
timestamp 1756801411
transform 1 0 5936 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_179
timestamp 1756801411
transform 1 0 5480 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_180
timestamp 1756801411
transform 1 0 4566 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_181
timestamp 1756801411
transform 1 0 5022 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_182
timestamp 1756801411
transform 1 0 4566 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_183
timestamp 1756801411
transform 1 0 5022 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_184
timestamp 1756801411
transform 1 0 3652 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_185
timestamp 1756801411
transform 1 0 4110 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_186
timestamp 1756801411
transform 1 0 3652 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_187
timestamp 1756801411
transform 1 0 4110 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_188
timestamp 1756801411
transform 1 0 2740 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_189
timestamp 1756801411
transform 1 0 3196 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_190
timestamp 1756801411
transform 1 0 2740 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_191
timestamp 1756801411
transform 1 0 3196 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_192
timestamp 1756801411
transform 1 0 1826 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_193
timestamp 1756801411
transform 1 0 2282 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_194
timestamp 1756801411
transform 1 0 2282 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_195
timestamp 1756801411
transform 1 0 1826 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_196
timestamp 1756801411
transform 1 0 912 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_197
timestamp 1756801411
transform 1 0 1370 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_198
timestamp 1756801411
transform 1 0 1370 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_199
timestamp 1756801411
transform 1 0 912 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_200
timestamp 1756801411
transform 1 0 0 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_201
timestamp 1756801411
transform 1 0 456 0 1 -1982
box 0 -20 400 440
use unit_Cap  unit_Cap_202
timestamp 1756801411
transform 1 0 456 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_203
timestamp 1756801411
transform 1 0 0 0 1 -2484
box 0 -20 400 440
use unit_Cap  unit_Cap_204
timestamp 1756801411
transform 1 0 15086 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_205
timestamp 1756801411
transform 1 0 14630 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_206
timestamp 1756801411
transform 1 0 14172 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_207
timestamp 1756801411
transform 1 0 13716 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_208
timestamp 1756801411
transform 1 0 13260 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_209
timestamp 1756801411
transform 1 0 12802 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_210
timestamp 1756801411
transform 1 0 12346 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_211
timestamp 1756801411
transform 1 0 11890 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_212
timestamp 1756801411
transform 1 0 11432 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_213
timestamp 1756801411
transform 1 0 10976 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_214
timestamp 1756801411
transform 1 0 10520 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_215
timestamp 1756801411
transform 1 0 10062 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_216
timestamp 1756801411
transform 1 0 9606 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_217
timestamp 1756801411
transform 1 0 9150 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_218
timestamp 1756801411
transform 1 0 8692 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_219
timestamp 1756801411
transform 1 0 8236 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_220
timestamp 1756801411
transform 1 0 7762 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_221
timestamp 1756801411
transform 1 0 7306 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_222
timestamp 1756801411
transform 1 0 6850 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_223
timestamp 1756801411
transform 1 0 6392 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_224
timestamp 1756801411
transform 1 0 5936 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_225
timestamp 1756801411
transform 1 0 5480 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_226
timestamp 1756801411
transform 1 0 4566 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_227
timestamp 1756801411
transform 1 0 5022 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_228
timestamp 1756801411
transform 1 0 3652 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_229
timestamp 1756801411
transform 1 0 4110 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_230
timestamp 1756801411
transform 1 0 2740 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_231
timestamp 1756801411
transform 1 0 3196 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_232
timestamp 1756801411
transform 1 0 2282 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_233
timestamp 1756801411
transform 1 0 1826 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_234
timestamp 1756801411
transform 1 0 1370 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_235
timestamp 1756801411
transform 1 0 912 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_236
timestamp 1756801411
transform 1 0 456 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_237
timestamp 1756801411
transform 1 0 0 0 1 -2976
box 0 -20 400 440
use unit_Cap  unit_Cap_238
timestamp 1756801411
transform 1 0 0 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_239
timestamp 1756801411
transform 1 0 456 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_240
timestamp 1756801411
transform 1 0 0 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_241
timestamp 1756801411
transform 1 0 456 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_242
timestamp 1756801411
transform 1 0 912 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_243
timestamp 1756801411
transform 1 0 1370 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_244
timestamp 1756801411
transform 1 0 912 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_245
timestamp 1756801411
transform 1 0 1370 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_246
timestamp 1756801411
transform 1 0 1826 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_247
timestamp 1756801411
transform 1 0 2282 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_248
timestamp 1756801411
transform 1 0 1826 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_249
timestamp 1756801411
transform 1 0 2282 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_250
timestamp 1756801411
transform 1 0 3652 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_251
timestamp 1756801411
transform 1 0 3652 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_252
timestamp 1756801411
transform 1 0 2740 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_253
timestamp 1756801411
transform 1 0 3196 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_254
timestamp 1756801411
transform 1 0 2740 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_255
timestamp 1756801411
transform 1 0 3196 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_256
timestamp 1756801411
transform 1 0 4110 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_257
timestamp 1756801411
transform 1 0 4566 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_258
timestamp 1756801411
transform 1 0 4110 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_259
timestamp 1756801411
transform 1 0 4566 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_260
timestamp 1756801411
transform 1 0 5022 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_261
timestamp 1756801411
transform 1 0 5480 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_262
timestamp 1756801411
transform 1 0 5022 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_263
timestamp 1756801411
transform 1 0 5480 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_264
timestamp 1756801411
transform 1 0 5936 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_265
timestamp 1756801411
transform 1 0 6392 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_266
timestamp 1756801411
transform 1 0 5936 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_267
timestamp 1756801411
transform 1 0 6392 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_268
timestamp 1756801411
transform 1 0 6850 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_269
timestamp 1756801411
transform 1 0 7306 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_270
timestamp 1756801411
transform 1 0 6850 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_271
timestamp 1756801411
transform 1 0 7306 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_272
timestamp 1756801411
transform 1 0 7762 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_273
timestamp 1756801411
transform 1 0 8236 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_274
timestamp 1756801411
transform 1 0 7762 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_275
timestamp 1756801411
transform 1 0 8236 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_276
timestamp 1756801411
transform 1 0 9150 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_277
timestamp 1756801411
transform 1 0 8692 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_278
timestamp 1756801411
transform 1 0 9150 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_279
timestamp 1756801411
transform 1 0 8692 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_280
timestamp 1756801411
transform 1 0 10062 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_281
timestamp 1756801411
transform 1 0 9606 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_282
timestamp 1756801411
transform 1 0 10062 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_283
timestamp 1756801411
transform 1 0 9606 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_284
timestamp 1756801411
transform 1 0 10976 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_285
timestamp 1756801411
transform 1 0 10520 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_286
timestamp 1756801411
transform 1 0 10976 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_287
timestamp 1756801411
transform 1 0 10520 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_288
timestamp 1756801411
transform 1 0 11890 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_289
timestamp 1756801411
transform 1 0 11432 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_290
timestamp 1756801411
transform 1 0 11890 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_291
timestamp 1756801411
transform 1 0 11432 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_292
timestamp 1756801411
transform 1 0 12346 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_293
timestamp 1756801411
transform 1 0 12802 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_294
timestamp 1756801411
transform 1 0 12346 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_295
timestamp 1756801411
transform 1 0 12802 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_296
timestamp 1756801411
transform 1 0 13260 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_297
timestamp 1756801411
transform 1 0 13716 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_298
timestamp 1756801411
transform 1 0 13260 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_299
timestamp 1756801411
transform 1 0 13716 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_300
timestamp 1756801411
transform 1 0 14172 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_301
timestamp 1756801411
transform 1 0 14630 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_302
timestamp 1756801411
transform 1 0 14172 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_303
timestamp 1756801411
transform 1 0 14630 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_304
timestamp 1756801411
transform 1 0 15086 0 1 -4464
box 0 -20 400 440
use unit_Cap  unit_Cap_305
timestamp 1756801411
transform 1 0 15086 0 1 -3972
box 0 -20 400 440
use unit_Cap  unit_Cap_306
timestamp 1756801411
transform 1 0 0 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_307
timestamp 1756801411
transform 1 0 456 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_308
timestamp 1756801411
transform 1 0 912 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_309
timestamp 1756801411
transform 1 0 1370 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_310
timestamp 1756801411
transform 1 0 1826 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_311
timestamp 1756801411
transform 1 0 2282 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_312
timestamp 1756801411
transform 1 0 3652 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_313
timestamp 1756801411
transform 1 0 2740 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_314
timestamp 1756801411
transform 1 0 3196 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_315
timestamp 1756801411
transform 1 0 4110 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_316
timestamp 1756801411
transform 1 0 4566 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_317
timestamp 1756801411
transform 1 0 5022 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_318
timestamp 1756801411
transform 1 0 5480 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_319
timestamp 1756801411
transform 1 0 5936 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_320
timestamp 1756801411
transform 1 0 6392 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_321
timestamp 1756801411
transform 1 0 6850 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_322
timestamp 1756801411
transform 1 0 7306 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_323
timestamp 1756801411
transform 1 0 7762 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_324
timestamp 1756801411
transform 1 0 8236 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_325
timestamp 1756801411
transform 1 0 8692 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_326
timestamp 1756801411
transform 1 0 9150 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_327
timestamp 1756801411
transform 1 0 9606 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_328
timestamp 1756801411
transform 1 0 10062 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_329
timestamp 1756801411
transform 1 0 10520 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_330
timestamp 1756801411
transform 1 0 10976 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_331
timestamp 1756801411
transform 1 0 11432 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_332
timestamp 1756801411
transform 1 0 11890 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_333
timestamp 1756801411
transform 1 0 12346 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_334
timestamp 1756801411
transform 1 0 12802 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_335
timestamp 1756801411
transform 1 0 13260 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_336
timestamp 1756801411
transform 1 0 13716 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_337
timestamp 1756801411
transform 1 0 14172 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_338
timestamp 1756801411
transform 1 0 14630 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_339
timestamp 1756801411
transform 1 0 15086 0 1 -3470
box 0 -20 400 440
use unit_Cap  unit_Cap_340
timestamp 1756801411
transform 1 0 15086 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_341
timestamp 1756801411
transform 1 0 15086 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_342
timestamp 1756801411
transform 1 0 14172 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_343
timestamp 1756801411
transform 1 0 14630 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_344
timestamp 1756801411
transform 1 0 14172 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_345
timestamp 1756801411
transform 1 0 14630 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_346
timestamp 1756801411
transform 1 0 13716 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_347
timestamp 1756801411
transform 1 0 13260 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_348
timestamp 1756801411
transform 1 0 13260 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_349
timestamp 1756801411
transform 1 0 13716 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_350
timestamp 1756801411
transform 1 0 12802 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_351
timestamp 1756801411
transform 1 0 12346 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_352
timestamp 1756801411
transform 1 0 12346 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_353
timestamp 1756801411
transform 1 0 12802 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_354
timestamp 1756801411
transform 1 0 11890 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_355
timestamp 1756801411
transform 1 0 11432 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_356
timestamp 1756801411
transform 1 0 11432 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_357
timestamp 1756801411
transform 1 0 11890 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_358
timestamp 1756801411
transform 1 0 10976 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_359
timestamp 1756801411
transform 1 0 10520 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_360
timestamp 1756801411
transform 1 0 10520 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_361
timestamp 1756801411
transform 1 0 10976 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_362
timestamp 1756801411
transform 1 0 10062 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_363
timestamp 1756801411
transform 1 0 9606 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_364
timestamp 1756801411
transform 1 0 9606 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_365
timestamp 1756801411
transform 1 0 10062 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_366
timestamp 1756801411
transform 1 0 9150 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_367
timestamp 1756801411
transform 1 0 8692 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_368
timestamp 1756801411
transform 1 0 8692 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_369
timestamp 1756801411
transform 1 0 9150 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_370
timestamp 1756801411
transform 1 0 8236 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_371
timestamp 1756801411
transform 1 0 7762 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_372
timestamp 1756801411
transform 1 0 8236 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_373
timestamp 1756801411
transform 1 0 7762 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_374
timestamp 1756801411
transform 1 0 7306 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_375
timestamp 1756801411
transform 1 0 6850 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_376
timestamp 1756801411
transform 1 0 7306 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_377
timestamp 1756801411
transform 1 0 6850 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_378
timestamp 1756801411
transform 1 0 6392 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_379
timestamp 1756801411
transform 1 0 5936 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_380
timestamp 1756801411
transform 1 0 6392 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_381
timestamp 1756801411
transform 1 0 5936 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_382
timestamp 1756801411
transform 1 0 5480 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_383
timestamp 1756801411
transform 1 0 5022 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_384
timestamp 1756801411
transform 1 0 5480 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_385
timestamp 1756801411
transform 1 0 5022 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_386
timestamp 1756801411
transform 1 0 4566 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_387
timestamp 1756801411
transform 1 0 4110 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_388
timestamp 1756801411
transform 1 0 4566 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_389
timestamp 1756801411
transform 1 0 4110 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_390
timestamp 1756801411
transform 1 0 3652 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_391
timestamp 1756801411
transform 1 0 3652 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_392
timestamp 1756801411
transform 1 0 3196 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_393
timestamp 1756801411
transform 1 0 2740 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_394
timestamp 1756801411
transform 1 0 3196 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_395
timestamp 1756801411
transform 1 0 2740 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_396
timestamp 1756801411
transform 1 0 1826 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_397
timestamp 1756801411
transform 1 0 2282 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_398
timestamp 1756801411
transform 1 0 1826 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_399
timestamp 1756801411
transform 1 0 2282 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_400
timestamp 1756801411
transform 1 0 912 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_401
timestamp 1756801411
transform 1 0 1370 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_402
timestamp 1756801411
transform 1 0 912 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_403
timestamp 1756801411
transform 1 0 1370 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_404
timestamp 1756801411
transform 1 0 0 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_405
timestamp 1756801411
transform 1 0 456 0 1 -4980
box 0 -20 400 440
use unit_Cap  unit_Cap_406
timestamp 1756801411
transform 1 0 0 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_407
timestamp 1756801411
transform 1 0 456 0 1 -5482
box 0 -20 400 440
use unit_Cap  unit_Cap_408
timestamp 1756801411
transform 1 0 15086 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_409
timestamp 1756801411
transform 1 0 14172 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_410
timestamp 1756801411
transform 1 0 14630 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_411
timestamp 1756801411
transform 1 0 13260 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_412
timestamp 1756801411
transform 1 0 13716 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_413
timestamp 1756801411
transform 1 0 12346 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_414
timestamp 1756801411
transform 1 0 12802 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_415
timestamp 1756801411
transform 1 0 11432 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_416
timestamp 1756801411
transform 1 0 11890 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_417
timestamp 1756801411
transform 1 0 10520 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_418
timestamp 1756801411
transform 1 0 10976 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_419
timestamp 1756801411
transform 1 0 9606 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_420
timestamp 1756801411
transform 1 0 10062 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_421
timestamp 1756801411
transform 1 0 8692 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_422
timestamp 1756801411
transform 1 0 9150 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_423
timestamp 1756801411
transform 1 0 8236 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_424
timestamp 1756801411
transform 1 0 7762 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_425
timestamp 1756801411
transform 1 0 7306 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_426
timestamp 1756801411
transform 1 0 6850 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_427
timestamp 1756801411
transform 1 0 6392 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_428
timestamp 1756801411
transform 1 0 5936 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_429
timestamp 1756801411
transform 1 0 5480 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_430
timestamp 1756801411
transform 1 0 5022 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_431
timestamp 1756801411
transform 1 0 4566 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_432
timestamp 1756801411
transform 1 0 4110 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_433
timestamp 1756801411
transform 1 0 3652 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_434
timestamp 1756801411
transform 1 0 3196 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_435
timestamp 1756801411
transform 1 0 2740 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_436
timestamp 1756801411
transform 1 0 1826 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_437
timestamp 1756801411
transform 1 0 2282 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_438
timestamp 1756801411
transform 1 0 912 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_439
timestamp 1756801411
transform 1 0 1370 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_440
timestamp 1756801411
transform 1 0 0 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_441
timestamp 1756801411
transform 1 0 456 0 1 -5974
box 0 -20 400 440
use unit_Cap  unit_Cap_442
timestamp 1756801411
transform 1 0 1 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_443
timestamp 1756801411
transform 1 0 457 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_444
timestamp 1756801411
transform 1 0 913 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_445
timestamp 1756801411
transform 1 0 1371 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_446
timestamp 1756801411
transform 1 0 1827 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_447
timestamp 1756801411
transform 1 0 2283 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_448
timestamp 1756801411
transform 1 0 2741 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_449
timestamp 1756801411
transform 1 0 3197 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_450
timestamp 1756801411
transform 1 0 4111 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_451
timestamp 1756801411
transform 1 0 4567 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_452
timestamp 1756801411
transform 1 0 3653 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_453
timestamp 1756801411
transform 1 0 5023 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_454
timestamp 1756801411
transform 1 0 5481 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_455
timestamp 1756801411
transform 1 0 5937 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_456
timestamp 1756801411
transform 1 0 6393 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_457
timestamp 1756801411
transform 1 0 6851 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_458
timestamp 1756801411
transform 1 0 7307 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_459
timestamp 1756801411
transform 1 0 7763 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_460
timestamp 1756801411
transform 1 0 8237 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_461
timestamp 1756801411
transform 1 0 9151 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_462
timestamp 1756801411
transform 1 0 8693 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_463
timestamp 1756801411
transform 1 0 10063 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_464
timestamp 1756801411
transform 1 0 9607 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_465
timestamp 1756801411
transform 1 0 10521 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_466
timestamp 1756801411
transform 1 0 10977 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_467
timestamp 1756801411
transform 1 0 11433 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_468
timestamp 1756801411
transform 1 0 11891 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_469
timestamp 1756801411
transform 1 0 12347 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_470
timestamp 1756801411
transform 1 0 12803 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_471
timestamp 1756801411
transform 1 0 13261 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_472
timestamp 1756801411
transform 1 0 13717 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_473
timestamp 1756801411
transform 1 0 14173 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_474
timestamp 1756801411
transform 1 0 14631 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_475
timestamp 1756801411
transform 1 0 15087 0 1 -6471
box 0 -20 400 440
use unit_Cap  unit_Cap_476
timestamp 1756801411
transform 1 0 15087 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_477
timestamp 1756801411
transform 1 0 15087 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_478
timestamp 1756801411
transform 1 0 14173 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_479
timestamp 1756801411
transform 1 0 14173 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_480
timestamp 1756801411
transform 1 0 14631 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_481
timestamp 1756801411
transform 1 0 14631 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_482
timestamp 1756801411
transform 1 0 13717 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_483
timestamp 1756801411
transform 1 0 13261 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_484
timestamp 1756801411
transform 1 0 13261 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_485
timestamp 1756801411
transform 1 0 13717 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_486
timestamp 1756801411
transform 1 0 12347 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_487
timestamp 1756801411
transform 1 0 12347 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_488
timestamp 1756801411
transform 1 0 12803 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_489
timestamp 1756801411
transform 1 0 12803 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_490
timestamp 1756801411
transform 1 0 11433 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_491
timestamp 1756801411
transform 1 0 11433 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_492
timestamp 1756801411
transform 1 0 11891 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_493
timestamp 1756801411
transform 1 0 11891 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_494
timestamp 1756801411
transform 1 0 10521 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_495
timestamp 1756801411
transform 1 0 10521 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_496
timestamp 1756801411
transform 1 0 10977 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_497
timestamp 1756801411
transform 1 0 10977 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_498
timestamp 1756801411
transform 1 0 10063 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_499
timestamp 1756801411
transform 1 0 9607 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_500
timestamp 1756801411
transform 1 0 10063 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_501
timestamp 1756801411
transform 1 0 9607 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_502
timestamp 1756801411
transform 1 0 9151 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_503
timestamp 1756801411
transform 1 0 8693 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_504
timestamp 1756801411
transform 1 0 9151 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_505
timestamp 1756801411
transform 1 0 8693 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_506
timestamp 1756801411
transform 1 0 7763 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_507
timestamp 1756801411
transform 1 0 7763 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_508
timestamp 1756801411
transform 1 0 8237 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_509
timestamp 1756801411
transform 1 0 8237 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_510
timestamp 1756801411
transform 1 0 6851 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_511
timestamp 1756801411
transform 1 0 6851 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_512
timestamp 1756801411
transform 1 0 7307 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_513
timestamp 1756801411
transform 1 0 7307 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_514
timestamp 1756801411
transform 1 0 5937 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_515
timestamp 1756801411
transform 1 0 5937 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_516
timestamp 1756801411
transform 1 0 6393 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_517
timestamp 1756801411
transform 1 0 6393 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_518
timestamp 1756801411
transform 1 0 5023 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_519
timestamp 1756801411
transform 1 0 5023 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_520
timestamp 1756801411
transform 1 0 5481 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_521
timestamp 1756801411
transform 1 0 5481 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_522
timestamp 1756801411
transform 1 0 4111 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_523
timestamp 1756801411
transform 1 0 4111 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_524
timestamp 1756801411
transform 1 0 4567 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_525
timestamp 1756801411
transform 1 0 4567 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_526
timestamp 1756801411
transform 1 0 2741 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_527
timestamp 1756801411
transform 1 0 2741 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_528
timestamp 1756801411
transform 1 0 3197 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_529
timestamp 1756801411
transform 1 0 3197 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_530
timestamp 1756801411
transform 1 0 3653 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_531
timestamp 1756801411
transform 1 0 3653 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_532
timestamp 1756801411
transform 1 0 1827 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_533
timestamp 1756801411
transform 1 0 1827 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_534
timestamp 1756801411
transform 1 0 2283 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_535
timestamp 1756801411
transform 1 0 2283 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_536
timestamp 1756801411
transform 1 0 913 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_537
timestamp 1756801411
transform 1 0 913 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_538
timestamp 1756801411
transform 1 0 1371 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_539
timestamp 1756801411
transform 1 0 1371 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_540
timestamp 1756801411
transform 1 0 1 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_541
timestamp 1756801411
transform 1 0 1 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_542
timestamp 1756801411
transform 1 0 457 0 1 -7479
box 0 -20 400 440
use unit_Cap  unit_Cap_543
timestamp 1756801411
transform 1 0 457 0 1 -6963
box 0 -20 400 440
use unit_Cap  unit_Cap_544
timestamp 1756801411
transform 1 0 15087 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_545
timestamp 1756801411
transform 1 0 15087 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_546
timestamp 1756801411
transform 1 0 14173 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_547
timestamp 1756801411
transform 1 0 14173 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_548
timestamp 1756801411
transform 1 0 14631 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_549
timestamp 1756801411
transform 1 0 14631 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_550
timestamp 1756801411
transform 1 0 13717 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_551
timestamp 1756801411
transform 1 0 13261 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_552
timestamp 1756801411
transform 1 0 13717 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_553
timestamp 1756801411
transform 1 0 13261 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_554
timestamp 1756801411
transform 1 0 12347 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_555
timestamp 1756801411
transform 1 0 12347 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_556
timestamp 1756801411
transform 1 0 12803 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_557
timestamp 1756801411
transform 1 0 12803 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_558
timestamp 1756801411
transform 1 0 11433 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_559
timestamp 1756801411
transform 1 0 11433 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_560
timestamp 1756801411
transform 1 0 11891 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_561
timestamp 1756801411
transform 1 0 11891 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_562
timestamp 1756801411
transform 1 0 10521 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_563
timestamp 1756801411
transform 1 0 10521 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_564
timestamp 1756801411
transform 1 0 10977 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_565
timestamp 1756801411
transform 1 0 10977 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_566
timestamp 1756801411
transform 1 0 10063 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_567
timestamp 1756801411
transform 1 0 9607 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_568
timestamp 1756801411
transform 1 0 10063 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_569
timestamp 1756801411
transform 1 0 9607 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_570
timestamp 1756801411
transform 1 0 9151 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_571
timestamp 1756801411
transform 1 0 8693 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_572
timestamp 1756801411
transform 1 0 9151 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_573
timestamp 1756801411
transform 1 0 8693 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_574
timestamp 1756801411
transform 1 0 7763 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_575
timestamp 1756801411
transform 1 0 7763 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_576
timestamp 1756801411
transform 1 0 8237 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_577
timestamp 1756801411
transform 1 0 8237 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_578
timestamp 1756801411
transform 1 0 6851 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_579
timestamp 1756801411
transform 1 0 6851 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_580
timestamp 1756801411
transform 1 0 7307 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_581
timestamp 1756801411
transform 1 0 7307 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_582
timestamp 1756801411
transform 1 0 5937 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_583
timestamp 1756801411
transform 1 0 5937 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_584
timestamp 1756801411
transform 1 0 6393 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_585
timestamp 1756801411
transform 1 0 6393 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_586
timestamp 1756801411
transform 1 0 5023 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_587
timestamp 1756801411
transform 1 0 5023 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_588
timestamp 1756801411
transform 1 0 5481 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_589
timestamp 1756801411
transform 1 0 5481 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_590
timestamp 1756801411
transform 1 0 4111 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_591
timestamp 1756801411
transform 1 0 4111 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_592
timestamp 1756801411
transform 1 0 4567 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_593
timestamp 1756801411
transform 1 0 4567 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_594
timestamp 1756801411
transform 1 0 2741 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_595
timestamp 1756801411
transform 1 0 2741 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_596
timestamp 1756801411
transform 1 0 3197 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_597
timestamp 1756801411
transform 1 0 3197 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_598
timestamp 1756801411
transform 1 0 3653 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_599
timestamp 1756801411
transform 1 0 3653 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_600
timestamp 1756801411
transform 1 0 1827 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_601
timestamp 1756801411
transform 1 0 1827 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_602
timestamp 1756801411
transform 1 0 2283 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_603
timestamp 1756801411
transform 1 0 2283 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_604
timestamp 1756801411
transform 1 0 913 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_605
timestamp 1756801411
transform 1 0 913 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_606
timestamp 1756801411
transform 1 0 1371 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_607
timestamp 1756801411
transform 1 0 1371 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_608
timestamp 1756801411
transform 1 0 1 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_609
timestamp 1756801411
transform 1 0 1 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_610
timestamp 1756801411
transform 1 0 457 0 1 -8473
box 0 -20 400 440
use unit_Cap  unit_Cap_611
timestamp 1756801411
transform 1 0 457 0 1 -7981
box 0 -20 400 440
use unit_Cap  unit_Cap_612
timestamp 1756801411
transform 1 0 15087 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_613
timestamp 1756801411
transform 1 0 15087 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_614
timestamp 1756801411
transform 1 0 14631 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_615
timestamp 1756801411
transform 1 0 14173 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_616
timestamp 1756801411
transform 1 0 14631 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_617
timestamp 1756801411
transform 1 0 14173 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_618
timestamp 1756801411
transform 1 0 13717 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_619
timestamp 1756801411
transform 1 0 13261 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_620
timestamp 1756801411
transform 1 0 13717 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_621
timestamp 1756801411
transform 1 0 13261 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_622
timestamp 1756801411
transform 1 0 12347 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_623
timestamp 1756801411
transform 1 0 12347 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_624
timestamp 1756801411
transform 1 0 12803 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_625
timestamp 1756801411
transform 1 0 12803 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_626
timestamp 1756801411
transform 1 0 11433 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_627
timestamp 1756801411
transform 1 0 11433 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_628
timestamp 1756801411
transform 1 0 11891 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_629
timestamp 1756801411
transform 1 0 11891 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_630
timestamp 1756801411
transform 1 0 10521 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_631
timestamp 1756801411
transform 1 0 10521 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_632
timestamp 1756801411
transform 1 0 10977 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_633
timestamp 1756801411
transform 1 0 10977 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_634
timestamp 1756801411
transform 1 0 10063 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_635
timestamp 1756801411
transform 1 0 9607 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_636
timestamp 1756801411
transform 1 0 9607 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_637
timestamp 1756801411
transform 1 0 10063 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_638
timestamp 1756801411
transform 1 0 9151 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_639
timestamp 1756801411
transform 1 0 8693 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_640
timestamp 1756801411
transform 1 0 8693 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_641
timestamp 1756801411
transform 1 0 9151 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_642
timestamp 1756801411
transform 1 0 8237 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_643
timestamp 1756801411
transform 1 0 7763 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_644
timestamp 1756801411
transform 1 0 8237 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_645
timestamp 1756801411
transform 1 0 7763 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_646
timestamp 1756801411
transform 1 0 6851 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_647
timestamp 1756801411
transform 1 0 6851 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_648
timestamp 1756801411
transform 1 0 7307 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_649
timestamp 1756801411
transform 1 0 7307 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_650
timestamp 1756801411
transform 1 0 5937 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_651
timestamp 1756801411
transform 1 0 5937 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_652
timestamp 1756801411
transform 1 0 6393 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_653
timestamp 1756801411
transform 1 0 6393 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_654
timestamp 1756801411
transform 1 0 5023 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_655
timestamp 1756801411
transform 1 0 5023 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_656
timestamp 1756801411
transform 1 0 5481 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_657
timestamp 1756801411
transform 1 0 5481 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_658
timestamp 1756801411
transform 1 0 4567 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_659
timestamp 1756801411
transform 1 0 4111 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_660
timestamp 1756801411
transform 1 0 4567 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_661
timestamp 1756801411
transform 1 0 4111 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_662
timestamp 1756801411
transform 1 0 2741 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_663
timestamp 1756801411
transform 1 0 2741 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_664
timestamp 1756801411
transform 1 0 3653 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_665
timestamp 1756801411
transform 1 0 3197 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_666
timestamp 1756801411
transform 1 0 3653 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_667
timestamp 1756801411
transform 1 0 3197 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_668
timestamp 1756801411
transform 1 0 1827 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_669
timestamp 1756801411
transform 1 0 1827 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_670
timestamp 1756801411
transform 1 0 2283 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_671
timestamp 1756801411
transform 1 0 2283 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_672
timestamp 1756801411
transform 1 0 1371 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_673
timestamp 1756801411
transform 1 0 913 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_674
timestamp 1756801411
transform 1 0 1371 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_675
timestamp 1756801411
transform 1 0 913 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_676
timestamp 1756801411
transform 1 0 457 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_677
timestamp 1756801411
transform 1 0 1 0 1 -8967
box 0 -20 400 440
use unit_Cap  unit_Cap_678
timestamp 1756801411
transform 1 0 457 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_679
timestamp 1756801411
transform 1 0 1 0 1 -9469
box 0 -20 400 440
use unit_Cap  unit_Cap_680
timestamp 1756801411
transform 1 0 15087 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_681
timestamp 1756801411
transform 1 0 15087 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_682
timestamp 1756801411
transform 1 0 14631 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_683
timestamp 1756801411
transform 1 0 14173 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_684
timestamp 1756801411
transform 1 0 14631 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_685
timestamp 1756801411
transform 1 0 14173 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_686
timestamp 1756801411
transform 1 0 13717 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_687
timestamp 1756801411
transform 1 0 13261 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_688
timestamp 1756801411
transform 1 0 13717 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_689
timestamp 1756801411
transform 1 0 13261 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_690
timestamp 1756801411
transform 1 0 12347 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_691
timestamp 1756801411
transform 1 0 12347 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_692
timestamp 1756801411
transform 1 0 12803 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_693
timestamp 1756801411
transform 1 0 12803 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_694
timestamp 1756801411
transform 1 0 11433 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_695
timestamp 1756801411
transform 1 0 11433 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_696
timestamp 1756801411
transform 1 0 11891 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_697
timestamp 1756801411
transform 1 0 11891 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_698
timestamp 1756801411
transform 1 0 10521 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_699
timestamp 1756801411
transform 1 0 10521 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_700
timestamp 1756801411
transform 1 0 10977 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_701
timestamp 1756801411
transform 1 0 10977 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_702
timestamp 1756801411
transform 1 0 9607 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_703
timestamp 1756801411
transform 1 0 10063 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_704
timestamp 1756801411
transform 1 0 10063 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_705
timestamp 1756801411
transform 1 0 9607 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_706
timestamp 1756801411
transform 1 0 8693 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_707
timestamp 1756801411
transform 1 0 9151 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_708
timestamp 1756801411
transform 1 0 9151 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_709
timestamp 1756801411
transform 1 0 8693 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_710
timestamp 1756801411
transform 1 0 8237 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_711
timestamp 1756801411
transform 1 0 7763 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_712
timestamp 1756801411
transform 1 0 8237 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_713
timestamp 1756801411
transform 1 0 7763 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_714
timestamp 1756801411
transform 1 0 6851 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_715
timestamp 1756801411
transform 1 0 6851 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_716
timestamp 1756801411
transform 1 0 7307 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_717
timestamp 1756801411
transform 1 0 7307 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_718
timestamp 1756801411
transform 1 0 5937 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_719
timestamp 1756801411
transform 1 0 5937 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_720
timestamp 1756801411
transform 1 0 6393 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_721
timestamp 1756801411
transform 1 0 6393 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_722
timestamp 1756801411
transform 1 0 5023 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_723
timestamp 1756801411
transform 1 0 5023 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_724
timestamp 1756801411
transform 1 0 5481 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_725
timestamp 1756801411
transform 1 0 5481 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_726
timestamp 1756801411
transform 1 0 4567 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_727
timestamp 1756801411
transform 1 0 4111 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_728
timestamp 1756801411
transform 1 0 4111 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_729
timestamp 1756801411
transform 1 0 4567 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_730
timestamp 1756801411
transform 1 0 2741 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_731
timestamp 1756801411
transform 1 0 2741 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_732
timestamp 1756801411
transform 1 0 3653 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_733
timestamp 1756801411
transform 1 0 3197 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_734
timestamp 1756801411
transform 1 0 3653 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_735
timestamp 1756801411
transform 1 0 3197 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_736
timestamp 1756801411
transform 1 0 1827 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_737
timestamp 1756801411
transform 1 0 1827 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_738
timestamp 1756801411
transform 1 0 2283 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_739
timestamp 1756801411
transform 1 0 2283 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_740
timestamp 1756801411
transform 1 0 1371 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_741
timestamp 1756801411
transform 1 0 913 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_742
timestamp 1756801411
transform 1 0 1371 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_743
timestamp 1756801411
transform 1 0 913 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_744
timestamp 1756801411
transform 1 0 457 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_745
timestamp 1756801411
transform 1 0 1 0 1 -9961
box 0 -20 400 440
use unit_Cap  unit_Cap_746
timestamp 1756801411
transform 1 0 457 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_747
timestamp 1756801411
transform 1 0 1 0 1 -10477
box 0 -20 400 440
use unit_Cap  unit_Cap_748
timestamp 1756801411
transform 1 0 15087 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_749
timestamp 1756801411
transform 1 0 15087 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_750
timestamp 1756801411
transform 1 0 14631 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_751
timestamp 1756801411
transform 1 0 14173 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_752
timestamp 1756801411
transform 1 0 14631 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_753
timestamp 1756801411
transform 1 0 14173 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_754
timestamp 1756801411
transform 1 0 13717 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_755
timestamp 1756801411
transform 1 0 13261 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_756
timestamp 1756801411
transform 1 0 13717 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_757
timestamp 1756801411
transform 1 0 13261 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_758
timestamp 1756801411
transform 1 0 12347 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_759
timestamp 1756801411
transform 1 0 12347 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_760
timestamp 1756801411
transform 1 0 12803 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_761
timestamp 1756801411
transform 1 0 12803 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_762
timestamp 1756801411
transform 1 0 11433 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_763
timestamp 1756801411
transform 1 0 11433 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_764
timestamp 1756801411
transform 1 0 11891 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_765
timestamp 1756801411
transform 1 0 11891 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_766
timestamp 1756801411
transform 1 0 10521 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_767
timestamp 1756801411
transform 1 0 10521 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_768
timestamp 1756801411
transform 1 0 10977 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_769
timestamp 1756801411
transform 1 0 10977 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_770
timestamp 1756801411
transform 1 0 10063 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_771
timestamp 1756801411
transform 1 0 9607 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_772
timestamp 1756801411
transform 1 0 10063 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_773
timestamp 1756801411
transform 1 0 9607 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_774
timestamp 1756801411
transform 1 0 9151 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_775
timestamp 1756801411
transform 1 0 8693 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_776
timestamp 1756801411
transform 1 0 9151 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_777
timestamp 1756801411
transform 1 0 8693 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_778
timestamp 1756801411
transform 1 0 8237 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_779
timestamp 1756801411
transform 1 0 7763 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_780
timestamp 1756801411
transform 1 0 8237 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_781
timestamp 1756801411
transform 1 0 7763 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_782
timestamp 1756801411
transform 1 0 6851 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_783
timestamp 1756801411
transform 1 0 6851 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_784
timestamp 1756801411
transform 1 0 7307 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_785
timestamp 1756801411
transform 1 0 7307 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_786
timestamp 1756801411
transform 1 0 5937 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_787
timestamp 1756801411
transform 1 0 5937 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_788
timestamp 1756801411
transform 1 0 6393 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_789
timestamp 1756801411
transform 1 0 6393 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_790
timestamp 1756801411
transform 1 0 5023 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_791
timestamp 1756801411
transform 1 0 5023 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_792
timestamp 1756801411
transform 1 0 5481 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_793
timestamp 1756801411
transform 1 0 5481 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_794
timestamp 1756801411
transform 1 0 4111 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_795
timestamp 1756801411
transform 1 0 4567 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_796
timestamp 1756801411
transform 1 0 4111 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_797
timestamp 1756801411
transform 1 0 4567 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_798
timestamp 1756801411
transform 1 0 2741 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_799
timestamp 1756801411
transform 1 0 2741 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_800
timestamp 1756801411
transform 1 0 3653 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_801
timestamp 1756801411
transform 1 0 3197 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_802
timestamp 1756801411
transform 1 0 3653 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_803
timestamp 1756801411
transform 1 0 3197 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_804
timestamp 1756801411
transform 1 0 1827 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_805
timestamp 1756801411
transform 1 0 1827 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_806
timestamp 1756801411
transform 1 0 2283 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_807
timestamp 1756801411
transform 1 0 2283 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_808
timestamp 1756801411
transform 1 0 1371 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_809
timestamp 1756801411
transform 1 0 913 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_810
timestamp 1756801411
transform 1 0 1371 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_811
timestamp 1756801411
transform 1 0 913 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_812
timestamp 1756801411
transform 1 0 457 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_813
timestamp 1756801411
transform 1 0 1 0 1 -10979
box 0 -20 400 440
use unit_Cap  unit_Cap_814
timestamp 1756801411
transform 1 0 457 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_815
timestamp 1756801411
transform 1 0 1 0 1 -11471
box 0 -20 400 440
use unit_Cap  unit_Cap_816
timestamp 1756801411
transform 1 0 1 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_817
timestamp 1756801411
transform 1 0 457 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_818
timestamp 1756801411
transform 1 0 913 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_819
timestamp 1756801411
transform 1 0 1371 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_820
timestamp 1756801411
transform 1 0 1827 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_821
timestamp 1756801411
transform 1 0 2283 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_822
timestamp 1756801411
transform 1 0 2741 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_823
timestamp 1756801411
transform 1 0 3653 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_824
timestamp 1756801411
transform 1 0 3197 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_825
timestamp 1756801411
transform 1 0 4111 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_826
timestamp 1756801411
transform 1 0 4567 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_827
timestamp 1756801411
transform 1 0 5023 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_828
timestamp 1756801411
transform 1 0 5481 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_829
timestamp 1756801411
transform 1 0 5937 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_830
timestamp 1756801411
transform 1 0 6393 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_831
timestamp 1756801411
transform 1 0 6851 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_832
timestamp 1756801411
transform 1 0 7307 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_833
timestamp 1756801411
transform 1 0 7763 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_834
timestamp 1756801411
transform 1 0 8237 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_835
timestamp 1756801411
transform 1 0 8693 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_836
timestamp 1756801411
transform 1 0 9151 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_837
timestamp 1756801411
transform 1 0 9607 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_838
timestamp 1756801411
transform 1 0 10063 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_839
timestamp 1756801411
transform 1 0 10521 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_840
timestamp 1756801411
transform 1 0 10977 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_841
timestamp 1756801411
transform 1 0 11433 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_842
timestamp 1756801411
transform 1 0 11891 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_843
timestamp 1756801411
transform 1 0 12347 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_844
timestamp 1756801411
transform 1 0 12803 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_845
timestamp 1756801411
transform 1 0 13717 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_846
timestamp 1756801411
transform 1 0 13261 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_847
timestamp 1756801411
transform 1 0 15087 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_848
timestamp 1756801411
transform 1 0 14631 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_849
timestamp 1756801411
transform 1 0 14173 0 1 -22461
box 0 -20 400 440
use unit_Cap  unit_Cap_850
timestamp 1756801411
transform 1 0 1 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_851
timestamp 1756801411
transform 1 0 457 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_852
timestamp 1756801411
transform 1 0 1 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_853
timestamp 1756801411
transform 1 0 457 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_854
timestamp 1756801411
transform 1 0 913 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_855
timestamp 1756801411
transform 1 0 1371 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_856
timestamp 1756801411
transform 1 0 913 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_857
timestamp 1756801411
transform 1 0 1371 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_858
timestamp 1756801411
transform 1 0 1827 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_859
timestamp 1756801411
transform 1 0 2283 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_860
timestamp 1756801411
transform 1 0 1827 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_861
timestamp 1756801411
transform 1 0 2283 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_862
timestamp 1756801411
transform 1 0 2741 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_863
timestamp 1756801411
transform 1 0 3653 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_864
timestamp 1756801411
transform 1 0 3197 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_865
timestamp 1756801411
transform 1 0 2741 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_866
timestamp 1756801411
transform 1 0 3653 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_867
timestamp 1756801411
transform 1 0 3197 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_868
timestamp 1756801411
transform 1 0 4111 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_869
timestamp 1756801411
transform 1 0 4567 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_870
timestamp 1756801411
transform 1 0 4111 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_871
timestamp 1756801411
transform 1 0 4567 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_872
timestamp 1756801411
transform 1 0 5023 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_873
timestamp 1756801411
transform 1 0 5481 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_874
timestamp 1756801411
transform 1 0 5023 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_875
timestamp 1756801411
transform 1 0 5481 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_876
timestamp 1756801411
transform 1 0 5937 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_877
timestamp 1756801411
transform 1 0 6393 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_878
timestamp 1756801411
transform 1 0 5937 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_879
timestamp 1756801411
transform 1 0 6393 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_880
timestamp 1756801411
transform 1 0 6851 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_881
timestamp 1756801411
transform 1 0 7307 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_882
timestamp 1756801411
transform 1 0 6851 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_883
timestamp 1756801411
transform 1 0 7307 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_884
timestamp 1756801411
transform 1 0 7763 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_885
timestamp 1756801411
transform 1 0 8237 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_886
timestamp 1756801411
transform 1 0 7763 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_887
timestamp 1756801411
transform 1 0 8237 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_888
timestamp 1756801411
transform 1 0 8693 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_889
timestamp 1756801411
transform 1 0 9151 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_890
timestamp 1756801411
transform 1 0 8693 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_891
timestamp 1756801411
transform 1 0 9151 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_892
timestamp 1756801411
transform 1 0 9607 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_893
timestamp 1756801411
transform 1 0 10063 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_894
timestamp 1756801411
transform 1 0 9607 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_895
timestamp 1756801411
transform 1 0 10063 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_896
timestamp 1756801411
transform 1 0 10521 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_897
timestamp 1756801411
transform 1 0 10977 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_898
timestamp 1756801411
transform 1 0 10521 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_899
timestamp 1756801411
transform 1 0 10977 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_900
timestamp 1756801411
transform 1 0 11433 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_901
timestamp 1756801411
transform 1 0 11891 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_902
timestamp 1756801411
transform 1 0 11433 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_903
timestamp 1756801411
transform 1 0 11891 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_904
timestamp 1756801411
transform 1 0 12347 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_905
timestamp 1756801411
transform 1 0 12803 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_906
timestamp 1756801411
transform 1 0 12347 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_907
timestamp 1756801411
transform 1 0 12803 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_908
timestamp 1756801411
transform 1 0 13717 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_909
timestamp 1756801411
transform 1 0 13261 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_910
timestamp 1756801411
transform 1 0 13717 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_911
timestamp 1756801411
transform 1 0 13261 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_912
timestamp 1756801411
transform 1 0 15087 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_913
timestamp 1756801411
transform 1 0 14631 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_914
timestamp 1756801411
transform 1 0 14173 0 1 -21467
box 0 -20 400 440
use unit_Cap  unit_Cap_915
timestamp 1756801411
transform 1 0 15087 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_916
timestamp 1756801411
transform 1 0 14631 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_917
timestamp 1756801411
transform 1 0 14173 0 1 -21969
box 0 -20 400 440
use unit_Cap  unit_Cap_918
timestamp 1756801411
transform 1 0 1 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_919
timestamp 1756801411
transform 1 0 457 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_920
timestamp 1756801411
transform 1 0 1 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_921
timestamp 1756801411
transform 1 0 457 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_922
timestamp 1756801411
transform 1 0 913 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_923
timestamp 1756801411
transform 1 0 1371 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_924
timestamp 1756801411
transform 1 0 913 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_925
timestamp 1756801411
transform 1 0 1371 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_926
timestamp 1756801411
transform 1 0 1827 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_927
timestamp 1756801411
transform 1 0 2283 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_928
timestamp 1756801411
transform 1 0 1827 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_929
timestamp 1756801411
transform 1 0 2283 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_930
timestamp 1756801411
transform 1 0 2741 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_931
timestamp 1756801411
transform 1 0 3653 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_932
timestamp 1756801411
transform 1 0 3197 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_933
timestamp 1756801411
transform 1 0 2741 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_934
timestamp 1756801411
transform 1 0 3653 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_935
timestamp 1756801411
transform 1 0 3197 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_936
timestamp 1756801411
transform 1 0 4111 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_937
timestamp 1756801411
transform 1 0 4567 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_938
timestamp 1756801411
transform 1 0 4111 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_939
timestamp 1756801411
transform 1 0 4567 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_940
timestamp 1756801411
transform 1 0 5023 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_941
timestamp 1756801411
transform 1 0 5481 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_942
timestamp 1756801411
transform 1 0 5023 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_943
timestamp 1756801411
transform 1 0 5481 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_944
timestamp 1756801411
transform 1 0 5937 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_945
timestamp 1756801411
transform 1 0 6393 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_946
timestamp 1756801411
transform 1 0 5937 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_947
timestamp 1756801411
transform 1 0 6393 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_948
timestamp 1756801411
transform 1 0 6851 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_949
timestamp 1756801411
transform 1 0 7307 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_950
timestamp 1756801411
transform 1 0 6851 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_951
timestamp 1756801411
transform 1 0 7307 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_952
timestamp 1756801411
transform 1 0 7763 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_953
timestamp 1756801411
transform 1 0 8237 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_954
timestamp 1756801411
transform 1 0 7763 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_955
timestamp 1756801411
transform 1 0 8237 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_956
timestamp 1756801411
transform 1 0 8693 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_957
timestamp 1756801411
transform 1 0 9151 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_958
timestamp 1756801411
transform 1 0 8693 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_959
timestamp 1756801411
transform 1 0 9151 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_960
timestamp 1756801411
transform 1 0 9607 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_961
timestamp 1756801411
transform 1 0 10063 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_962
timestamp 1756801411
transform 1 0 9607 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_963
timestamp 1756801411
transform 1 0 10063 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_964
timestamp 1756801411
transform 1 0 10521 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_965
timestamp 1756801411
transform 1 0 10977 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_966
timestamp 1756801411
transform 1 0 10521 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_967
timestamp 1756801411
transform 1 0 10977 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_968
timestamp 1756801411
transform 1 0 11433 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_969
timestamp 1756801411
transform 1 0 11891 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_970
timestamp 1756801411
transform 1 0 11433 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_971
timestamp 1756801411
transform 1 0 11891 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_972
timestamp 1756801411
transform 1 0 12347 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_973
timestamp 1756801411
transform 1 0 12803 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_974
timestamp 1756801411
transform 1 0 12347 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_975
timestamp 1756801411
transform 1 0 12803 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_976
timestamp 1756801411
transform 1 0 13717 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_977
timestamp 1756801411
transform 1 0 13261 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_978
timestamp 1756801411
transform 1 0 13717 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_979
timestamp 1756801411
transform 1 0 13261 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_980
timestamp 1756801411
transform 1 0 15087 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_981
timestamp 1756801411
transform 1 0 15087 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_982
timestamp 1756801411
transform 1 0 14631 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_983
timestamp 1756801411
transform 1 0 14173 0 1 -20951
box 0 -20 400 440
use unit_Cap  unit_Cap_984
timestamp 1756801411
transform 1 0 14631 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_985
timestamp 1756801411
transform 1 0 14173 0 1 -20459
box 0 -20 400 440
use unit_Cap  unit_Cap_986
timestamp 1756801411
transform 1 0 1 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_987
timestamp 1756801411
transform 1 0 457 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_988
timestamp 1756801411
transform 1 0 1 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_989
timestamp 1756801411
transform 1 0 457 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_990
timestamp 1756801411
transform 1 0 913 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_991
timestamp 1756801411
transform 1 0 1371 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_992
timestamp 1756801411
transform 1 0 913 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_993
timestamp 1756801411
transform 1 0 1371 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_994
timestamp 1756801411
transform 1 0 1827 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_995
timestamp 1756801411
transform 1 0 2283 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_996
timestamp 1756801411
transform 1 0 1827 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_997
timestamp 1756801411
transform 1 0 2283 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_998
timestamp 1756801411
transform 1 0 2741 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_999
timestamp 1756801411
transform 1 0 3197 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_1000
timestamp 1756801411
transform 1 0 3653 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_1001
timestamp 1756801411
transform 1 0 2741 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_1002
timestamp 1756801411
transform 1 0 3653 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_1003
timestamp 1756801411
transform 1 0 3197 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_1004
timestamp 1756801411
transform 1 0 4111 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_1005
timestamp 1756801411
transform 1 0 4567 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_1006
timestamp 1756801411
transform 1 0 4111 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_1007
timestamp 1756801411
transform 1 0 4567 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_1008
timestamp 1756801411
transform 1 0 5023 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_1009
timestamp 1756801411
transform 1 0 5481 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_1010
timestamp 1756801411
transform 1 0 5023 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_1011
timestamp 1756801411
transform 1 0 5481 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_1012
timestamp 1756801411
transform 1 0 5937 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_1013
timestamp 1756801411
transform 1 0 6393 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_1014
timestamp 1756801411
transform 1 0 5937 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_1015
timestamp 1756801411
transform 1 0 6393 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_1016
timestamp 1756801411
transform 1 0 6851 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_1017
timestamp 1756801411
transform 1 0 7307 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_1018
timestamp 1756801411
transform 1 0 6851 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_1019
timestamp 1756801411
transform 1 0 7307 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_1020
timestamp 1756801411
transform 1 0 7763 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_1021
timestamp 1756801411
transform 1 0 8237 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_1022
timestamp 1756801411
transform 1 0 7763 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_1023
timestamp 1756801411
transform 1 0 8237 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_1024
timestamp 1756801411
transform 1 0 8693 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_1025
timestamp 1756801411
transform 1 0 9151 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_1026
timestamp 1756801411
transform 1 0 8693 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_1027
timestamp 1756801411
transform 1 0 9151 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_1028
timestamp 1756801411
transform 1 0 9607 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_1029
timestamp 1756801411
transform 1 0 10063 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_1030
timestamp 1756801411
transform 1 0 9607 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_1031
timestamp 1756801411
transform 1 0 10063 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_1032
timestamp 1756801411
transform 1 0 10521 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_1033
timestamp 1756801411
transform 1 0 10977 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_1034
timestamp 1756801411
transform 1 0 10521 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_1035
timestamp 1756801411
transform 1 0 10977 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_1036
timestamp 1756801411
transform 1 0 11433 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_1037
timestamp 1756801411
transform 1 0 11891 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_1038
timestamp 1756801411
transform 1 0 11433 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_1039
timestamp 1756801411
transform 1 0 11891 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_1040
timestamp 1756801411
transform 1 0 12347 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_1041
timestamp 1756801411
transform 1 0 12803 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_1042
timestamp 1756801411
transform 1 0 12347 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_1043
timestamp 1756801411
transform 1 0 12803 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_1044
timestamp 1756801411
transform 1 0 13717 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_1045
timestamp 1756801411
transform 1 0 13261 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_1046
timestamp 1756801411
transform 1 0 13717 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_1047
timestamp 1756801411
transform 1 0 13261 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_1048
timestamp 1756801411
transform 1 0 15087 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_1049
timestamp 1756801411
transform 1 0 14173 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_1050
timestamp 1756801411
transform 1 0 14631 0 1 -19463
box 0 -20 400 440
use unit_Cap  unit_Cap_1051
timestamp 1756801411
transform 1 0 15087 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_1052
timestamp 1756801411
transform 1 0 14631 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_1053
timestamp 1756801411
transform 1 0 14173 0 1 -19957
box 0 -20 400 440
use unit_Cap  unit_Cap_1054
timestamp 1756801411
transform 1 0 1 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1055
timestamp 1756801411
transform 1 0 457 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1056
timestamp 1756801411
transform 1 0 1 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1057
timestamp 1756801411
transform 1 0 457 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1058
timestamp 1756801411
transform 1 0 913 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1059
timestamp 1756801411
transform 1 0 1371 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1060
timestamp 1756801411
transform 1 0 913 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1061
timestamp 1756801411
transform 1 0 1371 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1062
timestamp 1756801411
transform 1 0 1827 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1063
timestamp 1756801411
transform 1 0 2283 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1064
timestamp 1756801411
transform 1 0 1827 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1065
timestamp 1756801411
transform 1 0 2283 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1066
timestamp 1756801411
transform 1 0 2741 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1067
timestamp 1756801411
transform 1 0 3197 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1068
timestamp 1756801411
transform 1 0 3653 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1069
timestamp 1756801411
transform 1 0 2741 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1070
timestamp 1756801411
transform 1 0 3197 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1071
timestamp 1756801411
transform 1 0 3653 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1072
timestamp 1756801411
transform 1 0 4111 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1073
timestamp 1756801411
transform 1 0 4567 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1074
timestamp 1756801411
transform 1 0 4111 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1075
timestamp 1756801411
transform 1 0 4567 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1076
timestamp 1756801411
transform 1 0 5023 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1077
timestamp 1756801411
transform 1 0 5481 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1078
timestamp 1756801411
transform 1 0 5023 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1079
timestamp 1756801411
transform 1 0 5481 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1080
timestamp 1756801411
transform 1 0 5937 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1081
timestamp 1756801411
transform 1 0 6393 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1082
timestamp 1756801411
transform 1 0 5937 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1083
timestamp 1756801411
transform 1 0 6393 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1084
timestamp 1756801411
transform 1 0 6851 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1085
timestamp 1756801411
transform 1 0 7307 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1086
timestamp 1756801411
transform 1 0 6851 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1087
timestamp 1756801411
transform 1 0 7307 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1088
timestamp 1756801411
transform 1 0 7763 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1089
timestamp 1756801411
transform 1 0 8237 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1090
timestamp 1756801411
transform 1 0 7763 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1091
timestamp 1756801411
transform 1 0 8237 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1092
timestamp 1756801411
transform 1 0 8693 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1093
timestamp 1756801411
transform 1 0 9151 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1094
timestamp 1756801411
transform 1 0 8693 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1095
timestamp 1756801411
transform 1 0 9151 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1096
timestamp 1756801411
transform 1 0 9607 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1097
timestamp 1756801411
transform 1 0 10063 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1098
timestamp 1756801411
transform 1 0 9607 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1099
timestamp 1756801411
transform 1 0 10063 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1100
timestamp 1756801411
transform 1 0 10521 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1101
timestamp 1756801411
transform 1 0 10977 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1102
timestamp 1756801411
transform 1 0 10521 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1103
timestamp 1756801411
transform 1 0 10977 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1104
timestamp 1756801411
transform 1 0 11433 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1105
timestamp 1756801411
transform 1 0 11891 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1106
timestamp 1756801411
transform 1 0 11433 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1107
timestamp 1756801411
transform 1 0 11891 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1108
timestamp 1756801411
transform 1 0 12347 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1109
timestamp 1756801411
transform 1 0 12803 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1110
timestamp 1756801411
transform 1 0 12347 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1111
timestamp 1756801411
transform 1 0 12803 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1112
timestamp 1756801411
transform 1 0 13717 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1113
timestamp 1756801411
transform 1 0 13261 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1114
timestamp 1756801411
transform 1 0 13717 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1115
timestamp 1756801411
transform 1 0 13261 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1116
timestamp 1756801411
transform 1 0 15087 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1117
timestamp 1756801411
transform 1 0 14173 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1118
timestamp 1756801411
transform 1 0 14631 0 1 -18469
box 0 -20 400 440
use unit_Cap  unit_Cap_1119
timestamp 1756801411
transform 1 0 15087 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1120
timestamp 1756801411
transform 1 0 14173 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1121
timestamp 1756801411
transform 1 0 14631 0 1 -18971
box 0 -20 400 440
use unit_Cap  unit_Cap_1122
timestamp 1756801411
transform 1 0 1 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1123
timestamp 1756801411
transform 1 0 457 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1124
timestamp 1756801411
transform 1 0 1 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1125
timestamp 1756801411
transform 1 0 457 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1126
timestamp 1756801411
transform 1 0 913 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1127
timestamp 1756801411
transform 1 0 1371 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1128
timestamp 1756801411
transform 1 0 913 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1129
timestamp 1756801411
transform 1 0 1371 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1130
timestamp 1756801411
transform 1 0 1827 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1131
timestamp 1756801411
transform 1 0 2283 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1132
timestamp 1756801411
transform 1 0 1827 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1133
timestamp 1756801411
transform 1 0 2283 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1134
timestamp 1756801411
transform 1 0 2741 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1135
timestamp 1756801411
transform 1 0 3197 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1136
timestamp 1756801411
transform 1 0 3653 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1137
timestamp 1756801411
transform 1 0 2741 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1138
timestamp 1756801411
transform 1 0 3197 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1139
timestamp 1756801411
transform 1 0 3653 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1140
timestamp 1756801411
transform 1 0 4111 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1141
timestamp 1756801411
transform 1 0 4567 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1142
timestamp 1756801411
transform 1 0 4111 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1143
timestamp 1756801411
transform 1 0 4567 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1144
timestamp 1756801411
transform 1 0 5023 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1145
timestamp 1756801411
transform 1 0 5481 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1146
timestamp 1756801411
transform 1 0 5023 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1147
timestamp 1756801411
transform 1 0 5481 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1148
timestamp 1756801411
transform 1 0 5937 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1149
timestamp 1756801411
transform 1 0 6393 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1150
timestamp 1756801411
transform 1 0 5937 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1151
timestamp 1756801411
transform 1 0 6393 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1152
timestamp 1756801411
transform 1 0 6851 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1153
timestamp 1756801411
transform 1 0 7307 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1154
timestamp 1756801411
transform 1 0 6851 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1155
timestamp 1756801411
transform 1 0 7307 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1156
timestamp 1756801411
transform 1 0 7763 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1157
timestamp 1756801411
transform 1 0 8237 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1158
timestamp 1756801411
transform 1 0 7763 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1159
timestamp 1756801411
transform 1 0 8237 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1160
timestamp 1756801411
transform 1 0 8693 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1161
timestamp 1756801411
transform 1 0 9151 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1162
timestamp 1756801411
transform 1 0 8693 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1163
timestamp 1756801411
transform 1 0 9151 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1164
timestamp 1756801411
transform 1 0 9607 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1165
timestamp 1756801411
transform 1 0 10063 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1166
timestamp 1756801411
transform 1 0 9607 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1167
timestamp 1756801411
transform 1 0 10063 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1168
timestamp 1756801411
transform 1 0 10521 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1169
timestamp 1756801411
transform 1 0 10977 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1170
timestamp 1756801411
transform 1 0 10521 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1171
timestamp 1756801411
transform 1 0 10977 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1172
timestamp 1756801411
transform 1 0 11433 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1173
timestamp 1756801411
transform 1 0 11891 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1174
timestamp 1756801411
transform 1 0 11433 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1175
timestamp 1756801411
transform 1 0 11891 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1176
timestamp 1756801411
transform 1 0 12347 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1177
timestamp 1756801411
transform 1 0 12803 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1178
timestamp 1756801411
transform 1 0 12347 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1179
timestamp 1756801411
transform 1 0 12803 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1180
timestamp 1756801411
transform 1 0 13261 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1181
timestamp 1756801411
transform 1 0 13717 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1182
timestamp 1756801411
transform 1 0 13261 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1183
timestamp 1756801411
transform 1 0 13717 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1184
timestamp 1756801411
transform 1 0 15087 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1185
timestamp 1756801411
transform 1 0 14173 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1186
timestamp 1756801411
transform 1 0 14631 0 1 -17461
box 0 -20 400 440
use unit_Cap  unit_Cap_1187
timestamp 1756801411
transform 1 0 15087 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1188
timestamp 1756801411
transform 1 0 14173 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1189
timestamp 1756801411
transform 1 0 14631 0 1 -17953
box 0 -20 400 440
use unit_Cap  unit_Cap_1190
timestamp 1756801411
transform 1 0 0 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1191
timestamp 1756801411
transform 1 0 456 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1192
timestamp 1756801411
transform 1 0 0 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1193
timestamp 1756801411
transform 1 0 456 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1194
timestamp 1756801411
transform 1 0 912 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1195
timestamp 1756801411
transform 1 0 1370 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1196
timestamp 1756801411
transform 1 0 912 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1197
timestamp 1756801411
transform 1 0 1370 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1198
timestamp 1756801411
transform 1 0 1826 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1199
timestamp 1756801411
transform 1 0 2282 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1200
timestamp 1756801411
transform 1 0 1826 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1201
timestamp 1756801411
transform 1 0 2282 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1202
timestamp 1756801411
transform 1 0 2740 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1203
timestamp 1756801411
transform 1 0 3652 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1204
timestamp 1756801411
transform 1 0 3196 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1205
timestamp 1756801411
transform 1 0 2740 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1206
timestamp 1756801411
transform 1 0 3652 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1207
timestamp 1756801411
transform 1 0 3196 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1208
timestamp 1756801411
transform 1 0 4110 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1209
timestamp 1756801411
transform 1 0 4566 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1210
timestamp 1756801411
transform 1 0 4110 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1211
timestamp 1756801411
transform 1 0 4566 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1212
timestamp 1756801411
transform 1 0 5022 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1213
timestamp 1756801411
transform 1 0 5480 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1214
timestamp 1756801411
transform 1 0 5022 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1215
timestamp 1756801411
transform 1 0 5480 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1216
timestamp 1756801411
transform 1 0 5936 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1217
timestamp 1756801411
transform 1 0 6392 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1218
timestamp 1756801411
transform 1 0 5936 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1219
timestamp 1756801411
transform 1 0 6392 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1220
timestamp 1756801411
transform 1 0 6850 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1221
timestamp 1756801411
transform 1 0 7306 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1222
timestamp 1756801411
transform 1 0 6850 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1223
timestamp 1756801411
transform 1 0 7306 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1224
timestamp 1756801411
transform 1 0 7762 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1225
timestamp 1756801411
transform 1 0 8236 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1226
timestamp 1756801411
transform 1 0 7762 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1227
timestamp 1756801411
transform 1 0 8236 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1228
timestamp 1756801411
transform 1 0 8692 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1229
timestamp 1756801411
transform 1 0 9150 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1230
timestamp 1756801411
transform 1 0 8692 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1231
timestamp 1756801411
transform 1 0 9150 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1232
timestamp 1756801411
transform 1 0 9606 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1233
timestamp 1756801411
transform 1 0 10062 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1234
timestamp 1756801411
transform 1 0 9606 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1235
timestamp 1756801411
transform 1 0 10062 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1236
timestamp 1756801411
transform 1 0 10520 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1237
timestamp 1756801411
transform 1 0 10976 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1238
timestamp 1756801411
transform 1 0 10520 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1239
timestamp 1756801411
transform 1 0 10976 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1240
timestamp 1756801411
transform 1 0 11432 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1241
timestamp 1756801411
transform 1 0 11890 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1242
timestamp 1756801411
transform 1 0 11432 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1243
timestamp 1756801411
transform 1 0 11890 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1244
timestamp 1756801411
transform 1 0 12346 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1245
timestamp 1756801411
transform 1 0 12802 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1246
timestamp 1756801411
transform 1 0 12346 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1247
timestamp 1756801411
transform 1 0 12802 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1248
timestamp 1756801411
transform 1 0 13716 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1249
timestamp 1756801411
transform 1 0 13260 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1250
timestamp 1756801411
transform 1 0 13716 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1251
timestamp 1756801411
transform 1 0 13260 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1252
timestamp 1756801411
transform 1 0 15086 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1253
timestamp 1756801411
transform 1 0 14630 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1254
timestamp 1756801411
transform 1 0 14172 0 1 -16472
box 0 -20 400 440
use unit_Cap  unit_Cap_1255
timestamp 1756801411
transform 1 0 15086 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1256
timestamp 1756801411
transform 1 0 14630 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1257
timestamp 1756801411
transform 1 0 14172 0 1 -16964
box 0 -20 400 440
use unit_Cap  unit_Cap_1258
timestamp 1756801411
transform 1 0 0 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1259
timestamp 1756801411
transform 1 0 456 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1260
timestamp 1756801411
transform 1 0 912 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1261
timestamp 1756801411
transform 1 0 1370 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1262
timestamp 1756801411
transform 1 0 1826 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1263
timestamp 1756801411
transform 1 0 2282 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1264
timestamp 1756801411
transform 1 0 2740 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1265
timestamp 1756801411
transform 1 0 3652 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1266
timestamp 1756801411
transform 1 0 3196 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1267
timestamp 1756801411
transform 1 0 4110 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1268
timestamp 1756801411
transform 1 0 4566 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1269
timestamp 1756801411
transform 1 0 5022 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1270
timestamp 1756801411
transform 1 0 5480 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1271
timestamp 1756801411
transform 1 0 5936 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1272
timestamp 1756801411
transform 1 0 6392 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1273
timestamp 1756801411
transform 1 0 6850 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1274
timestamp 1756801411
transform 1 0 7306 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1275
timestamp 1756801411
transform 1 0 7762 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1276
timestamp 1756801411
transform 1 0 8236 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1277
timestamp 1756801411
transform 1 0 8692 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1278
timestamp 1756801411
transform 1 0 9150 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1279
timestamp 1756801411
transform 1 0 9606 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1280
timestamp 1756801411
transform 1 0 10062 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1281
timestamp 1756801411
transform 1 0 10520 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1282
timestamp 1756801411
transform 1 0 10976 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1283
timestamp 1756801411
transform 1 0 11432 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1284
timestamp 1756801411
transform 1 0 11890 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1285
timestamp 1756801411
transform 1 0 12346 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1286
timestamp 1756801411
transform 1 0 12802 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1287
timestamp 1756801411
transform 1 0 13716 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1288
timestamp 1756801411
transform 1 0 13260 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1289
timestamp 1756801411
transform 1 0 15086 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1290
timestamp 1756801411
transform 1 0 14630 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1291
timestamp 1756801411
transform 1 0 14172 0 1 -15970
box 0 -20 400 440
use unit_Cap  unit_Cap_1292
timestamp 1756801411
transform 1 0 0 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1293
timestamp 1756801411
transform 1 0 456 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1294
timestamp 1756801411
transform 1 0 0 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1295
timestamp 1756801411
transform 1 0 456 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1296
timestamp 1756801411
transform 1 0 912 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1297
timestamp 1756801411
transform 1 0 1370 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1298
timestamp 1756801411
transform 1 0 912 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1299
timestamp 1756801411
transform 1 0 1370 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1300
timestamp 1756801411
transform 1 0 1826 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1301
timestamp 1756801411
transform 1 0 2282 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1302
timestamp 1756801411
transform 1 0 1826 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1303
timestamp 1756801411
transform 1 0 2282 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1304
timestamp 1756801411
transform 1 0 2740 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1305
timestamp 1756801411
transform 1 0 3652 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1306
timestamp 1756801411
transform 1 0 3196 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1307
timestamp 1756801411
transform 1 0 2740 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1308
timestamp 1756801411
transform 1 0 3652 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1309
timestamp 1756801411
transform 1 0 3196 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1310
timestamp 1756801411
transform 1 0 4110 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1311
timestamp 1756801411
transform 1 0 4566 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1312
timestamp 1756801411
transform 1 0 4110 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1313
timestamp 1756801411
transform 1 0 4566 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1314
timestamp 1756801411
transform 1 0 5022 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1315
timestamp 1756801411
transform 1 0 5480 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1316
timestamp 1756801411
transform 1 0 5022 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1317
timestamp 1756801411
transform 1 0 5480 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1318
timestamp 1756801411
transform 1 0 5936 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1319
timestamp 1756801411
transform 1 0 6392 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1320
timestamp 1756801411
transform 1 0 5936 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1321
timestamp 1756801411
transform 1 0 6392 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1322
timestamp 1756801411
transform 1 0 6850 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1323
timestamp 1756801411
transform 1 0 7306 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1324
timestamp 1756801411
transform 1 0 6850 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1325
timestamp 1756801411
transform 1 0 7306 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1326
timestamp 1756801411
transform 1 0 7762 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1327
timestamp 1756801411
transform 1 0 8236 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1328
timestamp 1756801411
transform 1 0 7762 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1329
timestamp 1756801411
transform 1 0 8236 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1330
timestamp 1756801411
transform 1 0 8692 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1331
timestamp 1756801411
transform 1 0 9150 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1332
timestamp 1756801411
transform 1 0 8692 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1333
timestamp 1756801411
transform 1 0 9150 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1334
timestamp 1756801411
transform 1 0 9606 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1335
timestamp 1756801411
transform 1 0 10062 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1336
timestamp 1756801411
transform 1 0 9606 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1337
timestamp 1756801411
transform 1 0 10062 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1338
timestamp 1756801411
transform 1 0 10520 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1339
timestamp 1756801411
transform 1 0 10976 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1340
timestamp 1756801411
transform 1 0 10520 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1341
timestamp 1756801411
transform 1 0 10976 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1342
timestamp 1756801411
transform 1 0 11432 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1343
timestamp 1756801411
transform 1 0 11890 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1344
timestamp 1756801411
transform 1 0 11432 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1345
timestamp 1756801411
transform 1 0 11890 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1346
timestamp 1756801411
transform 1 0 12346 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1347
timestamp 1756801411
transform 1 0 12802 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1348
timestamp 1756801411
transform 1 0 12346 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1349
timestamp 1756801411
transform 1 0 12802 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1350
timestamp 1756801411
transform 1 0 13716 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1351
timestamp 1756801411
transform 1 0 13260 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1352
timestamp 1756801411
transform 1 0 13716 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1353
timestamp 1756801411
transform 1 0 13260 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1354
timestamp 1756801411
transform 1 0 14630 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1355
timestamp 1756801411
transform 1 0 14172 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1356
timestamp 1756801411
transform 1 0 15086 0 1 -14962
box 0 -20 400 440
use unit_Cap  unit_Cap_1357
timestamp 1756801411
transform 1 0 14630 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1358
timestamp 1756801411
transform 1 0 14172 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1359
timestamp 1756801411
transform 1 0 15086 0 1 -15454
box 0 -20 400 440
use unit_Cap  unit_Cap_1360
timestamp 1756801411
transform 1 0 0 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1361
timestamp 1756801411
transform 1 0 456 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1362
timestamp 1756801411
transform 1 0 0 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1363
timestamp 1756801411
transform 1 0 456 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1364
timestamp 1756801411
transform 1 0 912 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1365
timestamp 1756801411
transform 1 0 1370 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1366
timestamp 1756801411
transform 1 0 912 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1367
timestamp 1756801411
transform 1 0 1370 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1368
timestamp 1756801411
transform 1 0 1826 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1369
timestamp 1756801411
transform 1 0 2282 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1370
timestamp 1756801411
transform 1 0 1826 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1371
timestamp 1756801411
transform 1 0 2282 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1372
timestamp 1756801411
transform 1 0 2740 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1373
timestamp 1756801411
transform 1 0 3196 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1374
timestamp 1756801411
transform 1 0 3652 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1375
timestamp 1756801411
transform 1 0 2740 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1376
timestamp 1756801411
transform 1 0 3652 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1377
timestamp 1756801411
transform 1 0 3196 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1378
timestamp 1756801411
transform 1 0 4110 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1379
timestamp 1756801411
transform 1 0 4566 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1380
timestamp 1756801411
transform 1 0 4110 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1381
timestamp 1756801411
transform 1 0 4566 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1382
timestamp 1756801411
transform 1 0 5022 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1383
timestamp 1756801411
transform 1 0 5480 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1384
timestamp 1756801411
transform 1 0 5022 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1385
timestamp 1756801411
transform 1 0 5480 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1386
timestamp 1756801411
transform 1 0 5936 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1387
timestamp 1756801411
transform 1 0 6392 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1388
timestamp 1756801411
transform 1 0 5936 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1389
timestamp 1756801411
transform 1 0 6392 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1390
timestamp 1756801411
transform 1 0 6850 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1391
timestamp 1756801411
transform 1 0 7306 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1392
timestamp 1756801411
transform 1 0 6850 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1393
timestamp 1756801411
transform 1 0 7306 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1394
timestamp 1756801411
transform 1 0 7762 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1395
timestamp 1756801411
transform 1 0 8236 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1396
timestamp 1756801411
transform 1 0 7762 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1397
timestamp 1756801411
transform 1 0 8236 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1398
timestamp 1756801411
transform 1 0 8692 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1399
timestamp 1756801411
transform 1 0 9150 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1400
timestamp 1756801411
transform 1 0 8692 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1401
timestamp 1756801411
transform 1 0 9150 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1402
timestamp 1756801411
transform 1 0 9606 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1403
timestamp 1756801411
transform 1 0 10062 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1404
timestamp 1756801411
transform 1 0 9606 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1405
timestamp 1756801411
transform 1 0 10062 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1406
timestamp 1756801411
transform 1 0 10520 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1407
timestamp 1756801411
transform 1 0 10976 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1408
timestamp 1756801411
transform 1 0 10520 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1409
timestamp 1756801411
transform 1 0 10976 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1410
timestamp 1756801411
transform 1 0 11432 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1411
timestamp 1756801411
transform 1 0 11890 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1412
timestamp 1756801411
transform 1 0 11432 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1413
timestamp 1756801411
transform 1 0 11890 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1414
timestamp 1756801411
transform 1 0 12346 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1415
timestamp 1756801411
transform 1 0 12802 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1416
timestamp 1756801411
transform 1 0 12346 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1417
timestamp 1756801411
transform 1 0 12802 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1418
timestamp 1756801411
transform 1 0 13716 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1419
timestamp 1756801411
transform 1 0 13260 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1420
timestamp 1756801411
transform 1 0 13716 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1421
timestamp 1756801411
transform 1 0 13260 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1422
timestamp 1756801411
transform 1 0 14172 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1423
timestamp 1756801411
transform 1 0 14630 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1424
timestamp 1756801411
transform 1 0 15086 0 1 -13966
box 0 -20 400 440
use unit_Cap  unit_Cap_1425
timestamp 1756801411
transform 1 0 14630 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1426
timestamp 1756801411
transform 1 0 14172 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1427
timestamp 1756801411
transform 1 0 15086 0 1 -14460
box 0 -20 400 440
use unit_Cap  unit_Cap_1428
timestamp 1756801411
transform 1 0 0 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1429
timestamp 1756801411
transform 1 0 456 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1430
timestamp 1756801411
transform 1 0 0 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1431
timestamp 1756801411
transform 1 0 456 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1432
timestamp 1756801411
transform 1 0 912 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1433
timestamp 1756801411
transform 1 0 1370 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1434
timestamp 1756801411
transform 1 0 912 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1435
timestamp 1756801411
transform 1 0 1370 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1436
timestamp 1756801411
transform 1 0 1826 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1437
timestamp 1756801411
transform 1 0 2282 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1438
timestamp 1756801411
transform 1 0 1826 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1439
timestamp 1756801411
transform 1 0 2282 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1440
timestamp 1756801411
transform 1 0 2740 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1441
timestamp 1756801411
transform 1 0 3196 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1442
timestamp 1756801411
transform 1 0 3652 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1443
timestamp 1756801411
transform 1 0 2740 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1444
timestamp 1756801411
transform 1 0 3196 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1445
timestamp 1756801411
transform 1 0 3652 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1446
timestamp 1756801411
transform 1 0 4110 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1447
timestamp 1756801411
transform 1 0 4566 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1448
timestamp 1756801411
transform 1 0 4110 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1449
timestamp 1756801411
transform 1 0 4566 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1450
timestamp 1756801411
transform 1 0 5022 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1451
timestamp 1756801411
transform 1 0 5480 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1452
timestamp 1756801411
transform 1 0 5022 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1453
timestamp 1756801411
transform 1 0 5480 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1454
timestamp 1756801411
transform 1 0 5936 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1455
timestamp 1756801411
transform 1 0 6392 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1456
timestamp 1756801411
transform 1 0 5936 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1457
timestamp 1756801411
transform 1 0 6392 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1458
timestamp 1756801411
transform 1 0 6850 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1459
timestamp 1756801411
transform 1 0 7306 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1460
timestamp 1756801411
transform 1 0 6850 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1461
timestamp 1756801411
transform 1 0 7306 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1462
timestamp 1756801411
transform 1 0 7762 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1463
timestamp 1756801411
transform 1 0 8236 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1464
timestamp 1756801411
transform 1 0 7762 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1465
timestamp 1756801411
transform 1 0 8236 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1466
timestamp 1756801411
transform 1 0 8692 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1467
timestamp 1756801411
transform 1 0 9150 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1468
timestamp 1756801411
transform 1 0 8692 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1469
timestamp 1756801411
transform 1 0 9150 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1470
timestamp 1756801411
transform 1 0 9606 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1471
timestamp 1756801411
transform 1 0 10062 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1472
timestamp 1756801411
transform 1 0 9606 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1473
timestamp 1756801411
transform 1 0 10062 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1474
timestamp 1756801411
transform 1 0 10520 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1475
timestamp 1756801411
transform 1 0 10976 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1476
timestamp 1756801411
transform 1 0 10520 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1477
timestamp 1756801411
transform 1 0 10976 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1478
timestamp 1756801411
transform 1 0 11432 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1479
timestamp 1756801411
transform 1 0 11890 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1480
timestamp 1756801411
transform 1 0 11432 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1481
timestamp 1756801411
transform 1 0 11890 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1482
timestamp 1756801411
transform 1 0 12346 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1483
timestamp 1756801411
transform 1 0 12802 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1484
timestamp 1756801411
transform 1 0 12346 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1485
timestamp 1756801411
transform 1 0 12802 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1486
timestamp 1756801411
transform 1 0 13716 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1487
timestamp 1756801411
transform 1 0 13260 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1488
timestamp 1756801411
transform 1 0 13716 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1489
timestamp 1756801411
transform 1 0 13260 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1490
timestamp 1756801411
transform 1 0 14172 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1491
timestamp 1756801411
transform 1 0 14630 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1492
timestamp 1756801411
transform 1 0 15086 0 1 -13474
box 0 -20 400 440
use unit_Cap  unit_Cap_1493
timestamp 1756801411
transform 1 0 14172 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1494
timestamp 1756801411
transform 1 0 14630 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1495
timestamp 1756801411
transform 1 0 15086 0 1 -12972
box 0 -20 400 440
use unit_Cap  unit_Cap_1496
timestamp 1756801411
transform 1 0 0 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1497
timestamp 1756801411
transform 1 0 456 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1498
timestamp 1756801411
transform 1 0 0 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1499
timestamp 1756801411
transform 1 0 456 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1500
timestamp 1756801411
transform 1 0 912 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1501
timestamp 1756801411
transform 1 0 1370 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1502
timestamp 1756801411
transform 1 0 912 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1503
timestamp 1756801411
transform 1 0 1370 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1504
timestamp 1756801411
transform 1 0 1826 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1505
timestamp 1756801411
transform 1 0 2282 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1506
timestamp 1756801411
transform 1 0 1826 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1507
timestamp 1756801411
transform 1 0 2282 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1508
timestamp 1756801411
transform 1 0 2740 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1509
timestamp 1756801411
transform 1 0 3196 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1510
timestamp 1756801411
transform 1 0 3652 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1511
timestamp 1756801411
transform 1 0 2740 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1512
timestamp 1756801411
transform 1 0 3196 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1513
timestamp 1756801411
transform 1 0 3652 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1514
timestamp 1756801411
transform 1 0 4110 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1515
timestamp 1756801411
transform 1 0 4566 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1516
timestamp 1756801411
transform 1 0 4110 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1517
timestamp 1756801411
transform 1 0 4566 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1518
timestamp 1756801411
transform 1 0 5022 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1519
timestamp 1756801411
transform 1 0 5480 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1520
timestamp 1756801411
transform 1 0 5022 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1521
timestamp 1756801411
transform 1 0 5480 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1522
timestamp 1756801411
transform 1 0 5936 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1523
timestamp 1756801411
transform 1 0 6392 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1524
timestamp 1756801411
transform 1 0 5936 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1525
timestamp 1756801411
transform 1 0 6392 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1526
timestamp 1756801411
transform 1 0 6850 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1527
timestamp 1756801411
transform 1 0 7306 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1528
timestamp 1756801411
transform 1 0 6850 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1529
timestamp 1756801411
transform 1 0 7306 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1530
timestamp 1756801411
transform 1 0 7762 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1531
timestamp 1756801411
transform 1 0 8236 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1532
timestamp 1756801411
transform 1 0 7762 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1533
timestamp 1756801411
transform 1 0 8236 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1534
timestamp 1756801411
transform 1 0 8692 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1535
timestamp 1756801411
transform 1 0 9150 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1536
timestamp 1756801411
transform 1 0 8692 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1537
timestamp 1756801411
transform 1 0 9150 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1538
timestamp 1756801411
transform 1 0 9606 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1539
timestamp 1756801411
transform 1 0 10062 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1540
timestamp 1756801411
transform 1 0 9606 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1541
timestamp 1756801411
transform 1 0 10062 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1542
timestamp 1756801411
transform 1 0 10520 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1543
timestamp 1756801411
transform 1 0 10976 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1544
timestamp 1756801411
transform 1 0 10520 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1545
timestamp 1756801411
transform 1 0 10976 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1546
timestamp 1756801411
transform 1 0 11432 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1547
timestamp 1756801411
transform 1 0 11890 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1548
timestamp 1756801411
transform 1 0 11432 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1549
timestamp 1756801411
transform 1 0 11890 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1550
timestamp 1756801411
transform 1 0 12346 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1551
timestamp 1756801411
transform 1 0 12802 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1552
timestamp 1756801411
transform 1 0 12346 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1553
timestamp 1756801411
transform 1 0 12802 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1554
timestamp 1756801411
transform 1 0 13260 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1555
timestamp 1756801411
transform 1 0 13716 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1556
timestamp 1756801411
transform 1 0 13260 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1557
timestamp 1756801411
transform 1 0 13716 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1558
timestamp 1756801411
transform 1 0 14172 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1559
timestamp 1756801411
transform 1 0 14630 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1560
timestamp 1756801411
transform 1 0 15086 0 1 -12456
box 0 -20 400 440
use unit_Cap  unit_Cap_1561
timestamp 1756801411
transform 1 0 14172 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1562
timestamp 1756801411
transform 1 0 14630 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1563
timestamp 1756801411
transform 1 0 15086 0 1 -11964
box 0 -20 400 440
use unit_Cap  unit_Cap_1564
timestamp 1756801411
transform 1 0 1 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_1565
timestamp 1756801411
transform 1 0 913 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_1566
timestamp 1756801411
transform 1 0 457 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_1567
timestamp 1756801411
transform 1 0 1827 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_1568
timestamp 1756801411
transform 1 0 1371 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_1569
timestamp 1756801411
transform 1 0 2741 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_1570
timestamp 1756801411
transform 1 0 2283 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_1571
timestamp 1756801411
transform 1 0 1 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_1572
timestamp 1756801411
transform 1 0 1 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_1573
timestamp 1756801411
transform 1 0 913 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_1574
timestamp 1756801411
transform 1 0 457 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_1575
timestamp 1756801411
transform 1 0 913 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_1576
timestamp 1756801411
transform 1 0 457 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_1577
timestamp 1756801411
transform 1 0 1827 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_1578
timestamp 1756801411
transform 1 0 1371 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_1579
timestamp 1756801411
transform 1 0 1827 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_1580
timestamp 1756801411
transform 1 0 1371 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_1581
timestamp 1756801411
transform 1 0 2741 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_1582
timestamp 1756801411
transform 1 0 2283 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_1583
timestamp 1756801411
transform 1 0 2741 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_1584
timestamp 1756801411
transform 1 0 2283 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_1585
timestamp 1756801411
transform 1 0 1 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_1586
timestamp 1756801411
transform 1 0 913 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_1587
timestamp 1756801411
transform 1 0 457 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_1588
timestamp 1756801411
transform 1 0 1827 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_1589
timestamp 1756801411
transform 1 0 1371 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_1590
timestamp 1756801411
transform 1 0 2741 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_1591
timestamp 1756801411
transform 1 0 2283 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_1592
timestamp 1756801411
transform 1 0 1 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_1593
timestamp 1756801411
transform 1 0 1 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_1594
timestamp 1756801411
transform 1 0 913 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_1595
timestamp 1756801411
transform 1 0 913 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_1596
timestamp 1756801411
transform 1 0 457 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_1597
timestamp 1756801411
transform 1 0 457 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_1598
timestamp 1756801411
transform 1 0 1827 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_1599
timestamp 1756801411
transform 1 0 1827 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_1600
timestamp 1756801411
transform 1 0 1371 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_1601
timestamp 1756801411
transform 1 0 1371 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_1602
timestamp 1756801411
transform 1 0 2741 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_1603
timestamp 1756801411
transform 1 0 2741 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_1604
timestamp 1756801411
transform 1 0 2283 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_1605
timestamp 1756801411
transform 1 0 2283 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_1606
timestamp 1756801411
transform 1 0 1 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_1607
timestamp 1756801411
transform 1 0 0 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_1608
timestamp 1756801411
transform 1 0 913 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_1609
timestamp 1756801411
transform 1 0 912 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_1610
timestamp 1756801411
transform 1 0 457 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_1611
timestamp 1756801411
transform 1 0 456 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_1612
timestamp 1756801411
transform 1 0 1827 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_1613
timestamp 1756801411
transform 1 0 1826 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_1614
timestamp 1756801411
transform 1 0 1371 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_1615
timestamp 1756801411
transform 1 0 1370 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_1616
timestamp 1756801411
transform 1 0 2741 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_1617
timestamp 1756801411
transform 1 0 2740 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_1618
timestamp 1756801411
transform 1 0 2283 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_1619
timestamp 1756801411
transform 1 0 2282 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_1620
timestamp 1756801411
transform 1 0 0 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_1621
timestamp 1756801411
transform 1 0 0 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_1622
timestamp 1756801411
transform 1 0 912 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_1623
timestamp 1756801411
transform 1 0 912 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_1624
timestamp 1756801411
transform 1 0 456 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_1625
timestamp 1756801411
transform 1 0 456 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_1626
timestamp 1756801411
transform 1 0 1826 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_1627
timestamp 1756801411
transform 1 0 1826 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_1628
timestamp 1756801411
transform 1 0 1370 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_1629
timestamp 1756801411
transform 1 0 1370 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_1630
timestamp 1756801411
transform 1 0 2740 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_1631
timestamp 1756801411
transform 1 0 2740 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_1632
timestamp 1756801411
transform 1 0 2282 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_1633
timestamp 1756801411
transform 1 0 2282 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_1634
timestamp 1756801411
transform 1 0 0 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1635
timestamp 1756801411
transform 1 0 0 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1636
timestamp 1756801411
transform 1 0 912 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1637
timestamp 1756801411
transform 1 0 456 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1638
timestamp 1756801411
transform 1 0 912 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1639
timestamp 1756801411
transform 1 0 456 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1640
timestamp 1756801411
transform 1 0 1826 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1641
timestamp 1756801411
transform 1 0 1370 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1642
timestamp 1756801411
transform 1 0 1826 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1643
timestamp 1756801411
transform 1 0 1370 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1644
timestamp 1756801411
transform 1 0 2740 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1645
timestamp 1756801411
transform 1 0 2282 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1646
timestamp 1756801411
transform 1 0 2740 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1647
timestamp 1756801411
transform 1 0 2282 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1648
timestamp 1756801411
transform 1 0 0 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1649
timestamp 1756801411
transform 1 0 0 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1650
timestamp 1756801411
transform 1 0 912 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1651
timestamp 1756801411
transform 1 0 456 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1652
timestamp 1756801411
transform 1 0 912 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1653
timestamp 1756801411
transform 1 0 456 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1654
timestamp 1756801411
transform 1 0 1826 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1655
timestamp 1756801411
transform 1 0 1370 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1656
timestamp 1756801411
transform 1 0 1826 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1657
timestamp 1756801411
transform 1 0 1370 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1658
timestamp 1756801411
transform 1 0 2740 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1659
timestamp 1756801411
transform 1 0 2282 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1660
timestamp 1756801411
transform 1 0 2740 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1661
timestamp 1756801411
transform 1 0 2282 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1662
timestamp 1756801411
transform 1 0 0 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1663
timestamp 1756801411
transform 1 0 0 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1664
timestamp 1756801411
transform 1 0 912 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1665
timestamp 1756801411
transform 1 0 456 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1666
timestamp 1756801411
transform 1 0 912 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1667
timestamp 1756801411
transform 1 0 456 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1668
timestamp 1756801411
transform 1 0 1826 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1669
timestamp 1756801411
transform 1 0 1370 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1670
timestamp 1756801411
transform 1 0 1826 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1671
timestamp 1756801411
transform 1 0 1370 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1672
timestamp 1756801411
transform 1 0 2740 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1673
timestamp 1756801411
transform 1 0 2282 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1674
timestamp 1756801411
transform 1 0 2740 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1675
timestamp 1756801411
transform 1 0 2282 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1676
timestamp 1756801411
transform 1 0 0 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1677
timestamp 1756801411
transform 1 0 0 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1678
timestamp 1756801411
transform 1 0 912 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1679
timestamp 1756801411
transform 1 0 456 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1680
timestamp 1756801411
transform 1 0 912 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1681
timestamp 1756801411
transform 1 0 456 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1682
timestamp 1756801411
transform 1 0 1826 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1683
timestamp 1756801411
transform 1 0 1370 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1684
timestamp 1756801411
transform 1 0 1826 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1685
timestamp 1756801411
transform 1 0 1370 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1686
timestamp 1756801411
transform 1 0 2740 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1687
timestamp 1756801411
transform 1 0 2282 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1688
timestamp 1756801411
transform 1 0 2740 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1689
timestamp 1756801411
transform 1 0 2282 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1690
timestamp 1756801411
transform 1 0 0 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1691
timestamp 1756801411
transform 1 0 0 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1692
timestamp 1756801411
transform 1 0 912 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1693
timestamp 1756801411
transform 1 0 456 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1694
timestamp 1756801411
transform 1 0 912 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1695
timestamp 1756801411
transform 1 0 456 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1696
timestamp 1756801411
transform 1 0 1826 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1697
timestamp 1756801411
transform 1 0 1370 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1698
timestamp 1756801411
transform 1 0 1826 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1699
timestamp 1756801411
transform 1 0 1370 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1700
timestamp 1756801411
transform 1 0 2740 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1701
timestamp 1756801411
transform 1 0 2282 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1702
timestamp 1756801411
transform 1 0 2740 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1703
timestamp 1756801411
transform 1 0 2282 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1704
timestamp 1756801411
transform 1 0 15086 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1705
timestamp 1756801411
transform 1 0 14172 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1706
timestamp 1756801411
transform 1 0 14630 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1707
timestamp 1756801411
transform 1 0 13260 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1708
timestamp 1756801411
transform 1 0 13716 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1709
timestamp 1756801411
transform 1 0 12346 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1710
timestamp 1756801411
transform 1 0 12802 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1711
timestamp 1756801411
transform 1 0 11432 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1712
timestamp 1756801411
transform 1 0 11890 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1713
timestamp 1756801411
transform 1 0 10520 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1714
timestamp 1756801411
transform 1 0 10976 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1715
timestamp 1756801411
transform 1 0 9606 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1716
timestamp 1756801411
transform 1 0 10062 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1717
timestamp 1756801411
transform 1 0 8692 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1718
timestamp 1756801411
transform 1 0 9150 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1719
timestamp 1756801411
transform 1 0 7762 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1720
timestamp 1756801411
transform 1 0 8236 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1721
timestamp 1756801411
transform 1 0 6850 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1722
timestamp 1756801411
transform 1 0 7306 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1723
timestamp 1756801411
transform 1 0 5936 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1724
timestamp 1756801411
transform 1 0 6392 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1725
timestamp 1756801411
transform 1 0 5022 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1726
timestamp 1756801411
transform 1 0 5480 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1727
timestamp 1756801411
transform 1 0 4110 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1728
timestamp 1756801411
transform 1 0 4566 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1729
timestamp 1756801411
transform 1 0 3196 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1730
timestamp 1756801411
transform 1 0 3652 0 -1 -32007
box 0 -20 400 440
use unit_Cap  unit_Cap_1731
timestamp 1756801411
transform 1 0 15086 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1732
timestamp 1756801411
transform 1 0 15086 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1733
timestamp 1756801411
transform 1 0 14172 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1734
timestamp 1756801411
transform 1 0 14172 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1735
timestamp 1756801411
transform 1 0 14630 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1736
timestamp 1756801411
transform 1 0 14630 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1737
timestamp 1756801411
transform 1 0 13260 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1738
timestamp 1756801411
transform 1 0 13260 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1739
timestamp 1756801411
transform 1 0 13716 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1740
timestamp 1756801411
transform 1 0 13716 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1741
timestamp 1756801411
transform 1 0 12346 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1742
timestamp 1756801411
transform 1 0 12346 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1743
timestamp 1756801411
transform 1 0 12802 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1744
timestamp 1756801411
transform 1 0 12802 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1745
timestamp 1756801411
transform 1 0 11432 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1746
timestamp 1756801411
transform 1 0 11432 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1747
timestamp 1756801411
transform 1 0 11890 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1748
timestamp 1756801411
transform 1 0 11890 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1749
timestamp 1756801411
transform 1 0 10520 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1750
timestamp 1756801411
transform 1 0 10520 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1751
timestamp 1756801411
transform 1 0 10976 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1752
timestamp 1756801411
transform 1 0 10976 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1753
timestamp 1756801411
transform 1 0 9606 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1754
timestamp 1756801411
transform 1 0 9606 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1755
timestamp 1756801411
transform 1 0 10062 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1756
timestamp 1756801411
transform 1 0 10062 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1757
timestamp 1756801411
transform 1 0 8692 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1758
timestamp 1756801411
transform 1 0 8692 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1759
timestamp 1756801411
transform 1 0 9150 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1760
timestamp 1756801411
transform 1 0 9150 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1761
timestamp 1756801411
transform 1 0 7762 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1762
timestamp 1756801411
transform 1 0 7762 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1763
timestamp 1756801411
transform 1 0 8236 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1764
timestamp 1756801411
transform 1 0 8236 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1765
timestamp 1756801411
transform 1 0 6850 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1766
timestamp 1756801411
transform 1 0 6850 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1767
timestamp 1756801411
transform 1 0 7306 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1768
timestamp 1756801411
transform 1 0 7306 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1769
timestamp 1756801411
transform 1 0 5936 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1770
timestamp 1756801411
transform 1 0 5936 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1771
timestamp 1756801411
transform 1 0 6392 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1772
timestamp 1756801411
transform 1 0 6392 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1773
timestamp 1756801411
transform 1 0 5022 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1774
timestamp 1756801411
transform 1 0 5022 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1775
timestamp 1756801411
transform 1 0 5480 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1776
timestamp 1756801411
transform 1 0 5480 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1777
timestamp 1756801411
transform 1 0 4110 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1778
timestamp 1756801411
transform 1 0 4110 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1779
timestamp 1756801411
transform 1 0 4566 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1780
timestamp 1756801411
transform 1 0 4566 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1781
timestamp 1756801411
transform 1 0 3196 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1782
timestamp 1756801411
transform 1 0 3196 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1783
timestamp 1756801411
transform 1 0 3652 0 -1 -31013
box 0 -20 400 440
use unit_Cap  unit_Cap_1784
timestamp 1756801411
transform 1 0 3652 0 -1 -31515
box 0 -20 400 440
use unit_Cap  unit_Cap_1785
timestamp 1756801411
transform 1 0 15086 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1786
timestamp 1756801411
transform 1 0 15086 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1787
timestamp 1756801411
transform 1 0 14172 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1788
timestamp 1756801411
transform 1 0 14172 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1789
timestamp 1756801411
transform 1 0 14630 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1790
timestamp 1756801411
transform 1 0 14630 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1791
timestamp 1756801411
transform 1 0 13260 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1792
timestamp 1756801411
transform 1 0 13260 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1793
timestamp 1756801411
transform 1 0 13716 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1794
timestamp 1756801411
transform 1 0 13716 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1795
timestamp 1756801411
transform 1 0 12346 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1796
timestamp 1756801411
transform 1 0 12346 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1797
timestamp 1756801411
transform 1 0 12802 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1798
timestamp 1756801411
transform 1 0 12802 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1799
timestamp 1756801411
transform 1 0 11432 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1800
timestamp 1756801411
transform 1 0 11432 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1801
timestamp 1756801411
transform 1 0 11890 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1802
timestamp 1756801411
transform 1 0 11890 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1803
timestamp 1756801411
transform 1 0 10520 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1804
timestamp 1756801411
transform 1 0 10520 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1805
timestamp 1756801411
transform 1 0 10976 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1806
timestamp 1756801411
transform 1 0 10976 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1807
timestamp 1756801411
transform 1 0 9606 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1808
timestamp 1756801411
transform 1 0 9606 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1809
timestamp 1756801411
transform 1 0 10062 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1810
timestamp 1756801411
transform 1 0 10062 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1811
timestamp 1756801411
transform 1 0 8692 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1812
timestamp 1756801411
transform 1 0 8692 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1813
timestamp 1756801411
transform 1 0 9150 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1814
timestamp 1756801411
transform 1 0 9150 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1815
timestamp 1756801411
transform 1 0 7762 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1816
timestamp 1756801411
transform 1 0 7762 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1817
timestamp 1756801411
transform 1 0 8236 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1818
timestamp 1756801411
transform 1 0 8236 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1819
timestamp 1756801411
transform 1 0 6850 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1820
timestamp 1756801411
transform 1 0 6850 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1821
timestamp 1756801411
transform 1 0 7306 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1822
timestamp 1756801411
transform 1 0 7306 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1823
timestamp 1756801411
transform 1 0 5936 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1824
timestamp 1756801411
transform 1 0 5936 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1825
timestamp 1756801411
transform 1 0 6392 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1826
timestamp 1756801411
transform 1 0 6392 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1827
timestamp 1756801411
transform 1 0 5022 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1828
timestamp 1756801411
transform 1 0 5022 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1829
timestamp 1756801411
transform 1 0 5480 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1830
timestamp 1756801411
transform 1 0 5480 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1831
timestamp 1756801411
transform 1 0 4110 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1832
timestamp 1756801411
transform 1 0 4110 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1833
timestamp 1756801411
transform 1 0 4566 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1834
timestamp 1756801411
transform 1 0 4566 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1835
timestamp 1756801411
transform 1 0 3196 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1836
timestamp 1756801411
transform 1 0 3196 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1837
timestamp 1756801411
transform 1 0 3652 0 -1 -30005
box 0 -20 400 440
use unit_Cap  unit_Cap_1838
timestamp 1756801411
transform 1 0 3652 0 -1 -30521
box 0 -20 400 440
use unit_Cap  unit_Cap_1839
timestamp 1756801411
transform 1 0 15086 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1840
timestamp 1756801411
transform 1 0 15086 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1841
timestamp 1756801411
transform 1 0 14172 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1842
timestamp 1756801411
transform 1 0 14630 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1843
timestamp 1756801411
transform 1 0 14172 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1844
timestamp 1756801411
transform 1 0 14630 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1845
timestamp 1756801411
transform 1 0 13260 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1846
timestamp 1756801411
transform 1 0 13716 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1847
timestamp 1756801411
transform 1 0 13260 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1848
timestamp 1756801411
transform 1 0 13716 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1849
timestamp 1756801411
transform 1 0 12346 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1850
timestamp 1756801411
transform 1 0 12802 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1851
timestamp 1756801411
transform 1 0 12346 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1852
timestamp 1756801411
transform 1 0 12802 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1853
timestamp 1756801411
transform 1 0 11432 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1854
timestamp 1756801411
transform 1 0 11890 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1855
timestamp 1756801411
transform 1 0 11432 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1856
timestamp 1756801411
transform 1 0 11890 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1857
timestamp 1756801411
transform 1 0 10520 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1858
timestamp 1756801411
transform 1 0 10976 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1859
timestamp 1756801411
transform 1 0 10520 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1860
timestamp 1756801411
transform 1 0 10976 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1861
timestamp 1756801411
transform 1 0 9606 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1862
timestamp 1756801411
transform 1 0 10062 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1863
timestamp 1756801411
transform 1 0 9606 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1864
timestamp 1756801411
transform 1 0 10062 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1865
timestamp 1756801411
transform 1 0 8692 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1866
timestamp 1756801411
transform 1 0 9150 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1867
timestamp 1756801411
transform 1 0 8692 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1868
timestamp 1756801411
transform 1 0 9150 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1869
timestamp 1756801411
transform 1 0 7762 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1870
timestamp 1756801411
transform 1 0 8236 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1871
timestamp 1756801411
transform 1 0 7762 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1872
timestamp 1756801411
transform 1 0 8236 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1873
timestamp 1756801411
transform 1 0 6850 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1874
timestamp 1756801411
transform 1 0 7306 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1875
timestamp 1756801411
transform 1 0 6850 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1876
timestamp 1756801411
transform 1 0 7306 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1877
timestamp 1756801411
transform 1 0 5936 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1878
timestamp 1756801411
transform 1 0 6392 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1879
timestamp 1756801411
transform 1 0 5936 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1880
timestamp 1756801411
transform 1 0 6392 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1881
timestamp 1756801411
transform 1 0 5022 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1882
timestamp 1756801411
transform 1 0 5480 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1883
timestamp 1756801411
transform 1 0 5022 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1884
timestamp 1756801411
transform 1 0 5480 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1885
timestamp 1756801411
transform 1 0 4110 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1886
timestamp 1756801411
transform 1 0 4566 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1887
timestamp 1756801411
transform 1 0 4110 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1888
timestamp 1756801411
transform 1 0 4566 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1889
timestamp 1756801411
transform 1 0 3196 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1890
timestamp 1756801411
transform 1 0 3652 0 -1 -29011
box 0 -20 400 440
use unit_Cap  unit_Cap_1891
timestamp 1756801411
transform 1 0 3196 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1892
timestamp 1756801411
transform 1 0 3652 0 -1 -29503
box 0 -20 400 440
use unit_Cap  unit_Cap_1893
timestamp 1756801411
transform 1 0 15086 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1894
timestamp 1756801411
transform 1 0 15086 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1895
timestamp 1756801411
transform 1 0 14172 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1896
timestamp 1756801411
transform 1 0 14630 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1897
timestamp 1756801411
transform 1 0 14172 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1898
timestamp 1756801411
transform 1 0 14630 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1899
timestamp 1756801411
transform 1 0 13260 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1900
timestamp 1756801411
transform 1 0 13716 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1901
timestamp 1756801411
transform 1 0 13260 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1902
timestamp 1756801411
transform 1 0 13716 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1903
timestamp 1756801411
transform 1 0 12346 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1904
timestamp 1756801411
transform 1 0 12802 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1905
timestamp 1756801411
transform 1 0 12346 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1906
timestamp 1756801411
transform 1 0 12802 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1907
timestamp 1756801411
transform 1 0 11432 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1908
timestamp 1756801411
transform 1 0 11890 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1909
timestamp 1756801411
transform 1 0 11432 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1910
timestamp 1756801411
transform 1 0 11890 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1911
timestamp 1756801411
transform 1 0 10520 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1912
timestamp 1756801411
transform 1 0 10976 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1913
timestamp 1756801411
transform 1 0 10520 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1914
timestamp 1756801411
transform 1 0 10976 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1915
timestamp 1756801411
transform 1 0 9606 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1916
timestamp 1756801411
transform 1 0 10062 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1917
timestamp 1756801411
transform 1 0 9606 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1918
timestamp 1756801411
transform 1 0 10062 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1919
timestamp 1756801411
transform 1 0 8692 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1920
timestamp 1756801411
transform 1 0 9150 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1921
timestamp 1756801411
transform 1 0 8692 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1922
timestamp 1756801411
transform 1 0 9150 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1923
timestamp 1756801411
transform 1 0 7762 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1924
timestamp 1756801411
transform 1 0 8236 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1925
timestamp 1756801411
transform 1 0 7762 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1926
timestamp 1756801411
transform 1 0 8236 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1927
timestamp 1756801411
transform 1 0 6850 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1928
timestamp 1756801411
transform 1 0 7306 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1929
timestamp 1756801411
transform 1 0 6850 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1930
timestamp 1756801411
transform 1 0 7306 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1931
timestamp 1756801411
transform 1 0 5936 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1932
timestamp 1756801411
transform 1 0 6392 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1933
timestamp 1756801411
transform 1 0 5936 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1934
timestamp 1756801411
transform 1 0 6392 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1935
timestamp 1756801411
transform 1 0 5022 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1936
timestamp 1756801411
transform 1 0 5480 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1937
timestamp 1756801411
transform 1 0 5022 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1938
timestamp 1756801411
transform 1 0 5480 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1939
timestamp 1756801411
transform 1 0 4110 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1940
timestamp 1756801411
transform 1 0 4566 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1941
timestamp 1756801411
transform 1 0 4110 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1942
timestamp 1756801411
transform 1 0 4566 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1943
timestamp 1756801411
transform 1 0 3196 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1944
timestamp 1756801411
transform 1 0 3652 0 -1 -28015
box 0 -20 400 440
use unit_Cap  unit_Cap_1945
timestamp 1756801411
transform 1 0 3196 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1946
timestamp 1756801411
transform 1 0 3652 0 -1 -28517
box 0 -20 400 440
use unit_Cap  unit_Cap_1947
timestamp 1756801411
transform 1 0 15086 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1948
timestamp 1756801411
transform 1 0 14172 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1949
timestamp 1756801411
transform 1 0 14630 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1950
timestamp 1756801411
transform 1 0 13260 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1951
timestamp 1756801411
transform 1 0 13716 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1952
timestamp 1756801411
transform 1 0 12346 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1953
timestamp 1756801411
transform 1 0 12802 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1954
timestamp 1756801411
transform 1 0 11432 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1955
timestamp 1756801411
transform 1 0 11890 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1956
timestamp 1756801411
transform 1 0 10520 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1957
timestamp 1756801411
transform 1 0 10976 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1958
timestamp 1756801411
transform 1 0 9606 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1959
timestamp 1756801411
transform 1 0 10062 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1960
timestamp 1756801411
transform 1 0 8692 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1961
timestamp 1756801411
transform 1 0 9150 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1962
timestamp 1756801411
transform 1 0 7762 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1963
timestamp 1756801411
transform 1 0 8236 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1964
timestamp 1756801411
transform 1 0 6850 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1965
timestamp 1756801411
transform 1 0 7306 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1966
timestamp 1756801411
transform 1 0 5936 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1967
timestamp 1756801411
transform 1 0 6392 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1968
timestamp 1756801411
transform 1 0 5022 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1969
timestamp 1756801411
transform 1 0 5480 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1970
timestamp 1756801411
transform 1 0 4110 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1971
timestamp 1756801411
transform 1 0 4566 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1972
timestamp 1756801411
transform 1 0 3196 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1973
timestamp 1756801411
transform 1 0 3652 0 -1 -27523
box 0 -20 400 440
use unit_Cap  unit_Cap_1974
timestamp 1756801411
transform 1 0 15086 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_1975
timestamp 1756801411
transform 1 0 15086 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_1976
timestamp 1756801411
transform 1 0 14172 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_1977
timestamp 1756801411
transform 1 0 14172 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_1978
timestamp 1756801411
transform 1 0 14630 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_1979
timestamp 1756801411
transform 1 0 14630 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_1980
timestamp 1756801411
transform 1 0 13260 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_1981
timestamp 1756801411
transform 1 0 13260 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_1982
timestamp 1756801411
transform 1 0 13716 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_1983
timestamp 1756801411
transform 1 0 13716 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_1984
timestamp 1756801411
transform 1 0 12346 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_1985
timestamp 1756801411
transform 1 0 12346 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_1986
timestamp 1756801411
transform 1 0 12802 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_1987
timestamp 1756801411
transform 1 0 12802 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_1988
timestamp 1756801411
transform 1 0 11432 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_1989
timestamp 1756801411
transform 1 0 11432 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_1990
timestamp 1756801411
transform 1 0 11890 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_1991
timestamp 1756801411
transform 1 0 11890 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_1992
timestamp 1756801411
transform 1 0 10520 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_1993
timestamp 1756801411
transform 1 0 10520 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_1994
timestamp 1756801411
transform 1 0 10976 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_1995
timestamp 1756801411
transform 1 0 10976 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_1996
timestamp 1756801411
transform 1 0 9606 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_1997
timestamp 1756801411
transform 1 0 9606 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_1998
timestamp 1756801411
transform 1 0 10062 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_1999
timestamp 1756801411
transform 1 0 10062 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_2000
timestamp 1756801411
transform 1 0 8692 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_2001
timestamp 1756801411
transform 1 0 8692 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_2002
timestamp 1756801411
transform 1 0 9150 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_2003
timestamp 1756801411
transform 1 0 9150 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_2004
timestamp 1756801411
transform 1 0 7762 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_2005
timestamp 1756801411
transform 1 0 7762 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_2006
timestamp 1756801411
transform 1 0 8236 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_2007
timestamp 1756801411
transform 1 0 8236 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_2008
timestamp 1756801411
transform 1 0 6850 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_2009
timestamp 1756801411
transform 1 0 6850 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_2010
timestamp 1756801411
transform 1 0 7306 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_2011
timestamp 1756801411
transform 1 0 7306 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_2012
timestamp 1756801411
transform 1 0 5936 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_2013
timestamp 1756801411
transform 1 0 5936 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_2014
timestamp 1756801411
transform 1 0 6392 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_2015
timestamp 1756801411
transform 1 0 6392 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_2016
timestamp 1756801411
transform 1 0 5022 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_2017
timestamp 1756801411
transform 1 0 5022 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_2018
timestamp 1756801411
transform 1 0 5480 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_2019
timestamp 1756801411
transform 1 0 5480 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_2020
timestamp 1756801411
transform 1 0 4110 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_2021
timestamp 1756801411
transform 1 0 4110 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_2022
timestamp 1756801411
transform 1 0 4566 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_2023
timestamp 1756801411
transform 1 0 4566 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_2024
timestamp 1756801411
transform 1 0 3196 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_2025
timestamp 1756801411
transform 1 0 3196 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_2026
timestamp 1756801411
transform 1 0 3652 0 -1 -26505
box 0 -20 400 440
use unit_Cap  unit_Cap_2027
timestamp 1756801411
transform 1 0 3652 0 -1 -27007
box 0 -20 400 440
use unit_Cap  unit_Cap_2028
timestamp 1756801411
transform 1 0 15087 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_2029
timestamp 1756801411
transform 1 0 15086 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_2030
timestamp 1756801411
transform 1 0 14173 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_2031
timestamp 1756801411
transform 1 0 14172 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_2032
timestamp 1756801411
transform 1 0 14631 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_2033
timestamp 1756801411
transform 1 0 14630 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_2034
timestamp 1756801411
transform 1 0 13261 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_2035
timestamp 1756801411
transform 1 0 13260 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_2036
timestamp 1756801411
transform 1 0 13717 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_2037
timestamp 1756801411
transform 1 0 13716 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_2038
timestamp 1756801411
transform 1 0 12347 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_2039
timestamp 1756801411
transform 1 0 12346 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_2040
timestamp 1756801411
transform 1 0 12803 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_2041
timestamp 1756801411
transform 1 0 12802 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_2042
timestamp 1756801411
transform 1 0 11433 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_2043
timestamp 1756801411
transform 1 0 11432 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_2044
timestamp 1756801411
transform 1 0 11891 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_2045
timestamp 1756801411
transform 1 0 11890 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_2046
timestamp 1756801411
transform 1 0 10521 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_2047
timestamp 1756801411
transform 1 0 10520 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_2048
timestamp 1756801411
transform 1 0 10977 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_2049
timestamp 1756801411
transform 1 0 10976 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_2050
timestamp 1756801411
transform 1 0 9607 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_2051
timestamp 1756801411
transform 1 0 9606 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_2052
timestamp 1756801411
transform 1 0 10063 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_2053
timestamp 1756801411
transform 1 0 10062 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_2054
timestamp 1756801411
transform 1 0 8693 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_2055
timestamp 1756801411
transform 1 0 8692 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_2056
timestamp 1756801411
transform 1 0 9151 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_2057
timestamp 1756801411
transform 1 0 9150 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_2058
timestamp 1756801411
transform 1 0 7763 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_2059
timestamp 1756801411
transform 1 0 7762 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_2060
timestamp 1756801411
transform 1 0 8237 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_2061
timestamp 1756801411
transform 1 0 8236 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_2062
timestamp 1756801411
transform 1 0 6851 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_2063
timestamp 1756801411
transform 1 0 6850 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_2064
timestamp 1756801411
transform 1 0 7307 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_2065
timestamp 1756801411
transform 1 0 7306 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_2066
timestamp 1756801411
transform 1 0 5937 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_2067
timestamp 1756801411
transform 1 0 5936 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_2068
timestamp 1756801411
transform 1 0 6393 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_2069
timestamp 1756801411
transform 1 0 6392 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_2070
timestamp 1756801411
transform 1 0 5023 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_2071
timestamp 1756801411
transform 1 0 5022 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_2072
timestamp 1756801411
transform 1 0 5481 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_2073
timestamp 1756801411
transform 1 0 5480 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_2074
timestamp 1756801411
transform 1 0 4111 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_2075
timestamp 1756801411
transform 1 0 4110 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_2076
timestamp 1756801411
transform 1 0 4567 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_2077
timestamp 1756801411
transform 1 0 4566 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_2078
timestamp 1756801411
transform 1 0 3197 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_2079
timestamp 1756801411
transform 1 0 3196 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_2080
timestamp 1756801411
transform 1 0 3653 0 -1 -25516
box 0 -20 400 440
use unit_Cap  unit_Cap_2081
timestamp 1756801411
transform 1 0 3652 0 -1 -26013
box 0 -20 400 440
use unit_Cap  unit_Cap_2082
timestamp 1756801411
transform 1 0 15087 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_2083
timestamp 1756801411
transform 1 0 15087 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_2084
timestamp 1756801411
transform 1 0 14173 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_2085
timestamp 1756801411
transform 1 0 14173 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_2086
timestamp 1756801411
transform 1 0 14631 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_2087
timestamp 1756801411
transform 1 0 14631 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_2088
timestamp 1756801411
transform 1 0 13261 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_2089
timestamp 1756801411
transform 1 0 13261 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_2090
timestamp 1756801411
transform 1 0 13717 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_2091
timestamp 1756801411
transform 1 0 13717 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_2092
timestamp 1756801411
transform 1 0 12347 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_2093
timestamp 1756801411
transform 1 0 12347 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_2094
timestamp 1756801411
transform 1 0 12803 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_2095
timestamp 1756801411
transform 1 0 12803 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_2096
timestamp 1756801411
transform 1 0 11433 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_2097
timestamp 1756801411
transform 1 0 11433 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_2098
timestamp 1756801411
transform 1 0 11891 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_2099
timestamp 1756801411
transform 1 0 11891 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_2100
timestamp 1756801411
transform 1 0 10521 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_2101
timestamp 1756801411
transform 1 0 10521 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_2102
timestamp 1756801411
transform 1 0 10977 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_2103
timestamp 1756801411
transform 1 0 10977 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_2104
timestamp 1756801411
transform 1 0 9607 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_2105
timestamp 1756801411
transform 1 0 9607 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_2106
timestamp 1756801411
transform 1 0 10063 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_2107
timestamp 1756801411
transform 1 0 10063 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_2108
timestamp 1756801411
transform 1 0 8693 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_2109
timestamp 1756801411
transform 1 0 8693 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_2110
timestamp 1756801411
transform 1 0 9151 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_2111
timestamp 1756801411
transform 1 0 9151 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_2112
timestamp 1756801411
transform 1 0 7763 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_2113
timestamp 1756801411
transform 1 0 7763 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_2114
timestamp 1756801411
transform 1 0 8237 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_2115
timestamp 1756801411
transform 1 0 8237 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_2116
timestamp 1756801411
transform 1 0 6851 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_2117
timestamp 1756801411
transform 1 0 6851 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_2118
timestamp 1756801411
transform 1 0 7307 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_2119
timestamp 1756801411
transform 1 0 7307 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_2120
timestamp 1756801411
transform 1 0 5937 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_2121
timestamp 1756801411
transform 1 0 5937 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_2122
timestamp 1756801411
transform 1 0 6393 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_2123
timestamp 1756801411
transform 1 0 6393 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_2124
timestamp 1756801411
transform 1 0 5023 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_2125
timestamp 1756801411
transform 1 0 5023 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_2126
timestamp 1756801411
transform 1 0 5481 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_2127
timestamp 1756801411
transform 1 0 5481 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_2128
timestamp 1756801411
transform 1 0 4111 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_2129
timestamp 1756801411
transform 1 0 4111 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_2130
timestamp 1756801411
transform 1 0 4567 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_2131
timestamp 1756801411
transform 1 0 4567 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_2132
timestamp 1756801411
transform 1 0 3197 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_2133
timestamp 1756801411
transform 1 0 3197 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_2134
timestamp 1756801411
transform 1 0 3653 0 -1 -24508
box 0 -20 400 440
use unit_Cap  unit_Cap_2135
timestamp 1756801411
transform 1 0 3653 0 -1 -25024
box 0 -20 400 440
use unit_Cap  unit_Cap_2136
timestamp 1756801411
transform 1 0 15087 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_2137
timestamp 1756801411
transform 1 0 15087 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_2138
timestamp 1756801411
transform 1 0 14173 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_2139
timestamp 1756801411
transform 1 0 14631 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_2140
timestamp 1756801411
transform 1 0 14173 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_2141
timestamp 1756801411
transform 1 0 14631 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_2142
timestamp 1756801411
transform 1 0 13261 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_2143
timestamp 1756801411
transform 1 0 13717 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_2144
timestamp 1756801411
transform 1 0 13261 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_2145
timestamp 1756801411
transform 1 0 13717 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_2146
timestamp 1756801411
transform 1 0 12347 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_2147
timestamp 1756801411
transform 1 0 12803 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_2148
timestamp 1756801411
transform 1 0 12347 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_2149
timestamp 1756801411
transform 1 0 12803 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_2150
timestamp 1756801411
transform 1 0 11433 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_2151
timestamp 1756801411
transform 1 0 11891 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_2152
timestamp 1756801411
transform 1 0 11433 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_2153
timestamp 1756801411
transform 1 0 11891 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_2154
timestamp 1756801411
transform 1 0 10521 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_2155
timestamp 1756801411
transform 1 0 10977 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_2156
timestamp 1756801411
transform 1 0 10521 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_2157
timestamp 1756801411
transform 1 0 10977 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_2158
timestamp 1756801411
transform 1 0 9607 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_2159
timestamp 1756801411
transform 1 0 10063 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_2160
timestamp 1756801411
transform 1 0 9607 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_2161
timestamp 1756801411
transform 1 0 10063 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_2162
timestamp 1756801411
transform 1 0 8693 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_2163
timestamp 1756801411
transform 1 0 9151 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_2164
timestamp 1756801411
transform 1 0 8693 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_2165
timestamp 1756801411
transform 1 0 9151 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_2166
timestamp 1756801411
transform 1 0 7763 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_2167
timestamp 1756801411
transform 1 0 8237 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_2168
timestamp 1756801411
transform 1 0 7763 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_2169
timestamp 1756801411
transform 1 0 8237 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_2170
timestamp 1756801411
transform 1 0 6851 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_2171
timestamp 1756801411
transform 1 0 7307 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_2172
timestamp 1756801411
transform 1 0 6851 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_2173
timestamp 1756801411
transform 1 0 7307 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_2174
timestamp 1756801411
transform 1 0 5937 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_2175
timestamp 1756801411
transform 1 0 6393 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_2176
timestamp 1756801411
transform 1 0 5937 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_2177
timestamp 1756801411
transform 1 0 6393 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_2178
timestamp 1756801411
transform 1 0 5023 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_2179
timestamp 1756801411
transform 1 0 5481 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_2180
timestamp 1756801411
transform 1 0 5023 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_2181
timestamp 1756801411
transform 1 0 5481 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_2182
timestamp 1756801411
transform 1 0 4111 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_2183
timestamp 1756801411
transform 1 0 4567 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_2184
timestamp 1756801411
transform 1 0 4111 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_2185
timestamp 1756801411
transform 1 0 4567 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_2186
timestamp 1756801411
transform 1 0 3197 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_2187
timestamp 1756801411
transform 1 0 3653 0 -1 -24006
box 0 -20 400 440
use unit_Cap  unit_Cap_2188
timestamp 1756801411
transform 1 0 3197 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_2189
timestamp 1756801411
transform 1 0 3653 0 -1 -23514
box 0 -20 400 440
use unit_Cap  unit_Cap_2190
timestamp 1756801411
transform 1 0 15087 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_2191
timestamp 1756801411
transform 1 0 15087 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_2192
timestamp 1756801411
transform 1 0 14173 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_2193
timestamp 1756801411
transform 1 0 14631 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_2194
timestamp 1756801411
transform 1 0 14173 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_2195
timestamp 1756801411
transform 1 0 14631 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_2196
timestamp 1756801411
transform 1 0 13261 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_2197
timestamp 1756801411
transform 1 0 13717 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_2198
timestamp 1756801411
transform 1 0 13261 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_2199
timestamp 1756801411
transform 1 0 13717 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_2200
timestamp 1756801411
transform 1 0 12347 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_2201
timestamp 1756801411
transform 1 0 12803 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_2202
timestamp 1756801411
transform 1 0 12347 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_2203
timestamp 1756801411
transform 1 0 12803 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_2204
timestamp 1756801411
transform 1 0 11433 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_2205
timestamp 1756801411
transform 1 0 11891 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_2206
timestamp 1756801411
transform 1 0 11433 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_2207
timestamp 1756801411
transform 1 0 11891 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_2208
timestamp 1756801411
transform 1 0 10521 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_2209
timestamp 1756801411
transform 1 0 10977 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_2210
timestamp 1756801411
transform 1 0 10521 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_2211
timestamp 1756801411
transform 1 0 10977 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_2212
timestamp 1756801411
transform 1 0 9607 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_2213
timestamp 1756801411
transform 1 0 10063 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_2214
timestamp 1756801411
transform 1 0 9607 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_2215
timestamp 1756801411
transform 1 0 10063 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_2216
timestamp 1756801411
transform 1 0 8693 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_2217
timestamp 1756801411
transform 1 0 9151 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_2218
timestamp 1756801411
transform 1 0 8693 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_2219
timestamp 1756801411
transform 1 0 9151 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_2220
timestamp 1756801411
transform 1 0 7763 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_2221
timestamp 1756801411
transform 1 0 8237 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_2222
timestamp 1756801411
transform 1 0 7763 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_2223
timestamp 1756801411
transform 1 0 8237 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_2224
timestamp 1756801411
transform 1 0 6851 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_2225
timestamp 1756801411
transform 1 0 7307 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_2226
timestamp 1756801411
transform 1 0 6851 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_2227
timestamp 1756801411
transform 1 0 7307 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_2228
timestamp 1756801411
transform 1 0 5937 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_2229
timestamp 1756801411
transform 1 0 6393 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_2230
timestamp 1756801411
transform 1 0 5937 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_2231
timestamp 1756801411
transform 1 0 6393 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_2232
timestamp 1756801411
transform 1 0 5023 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_2233
timestamp 1756801411
transform 1 0 5481 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_2234
timestamp 1756801411
transform 1 0 5023 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_2235
timestamp 1756801411
transform 1 0 5481 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_2236
timestamp 1756801411
transform 1 0 4111 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_2237
timestamp 1756801411
transform 1 0 4567 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_2238
timestamp 1756801411
transform 1 0 4111 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_2239
timestamp 1756801411
transform 1 0 4567 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_2240
timestamp 1756801411
transform 1 0 3197 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_2241
timestamp 1756801411
transform 1 0 3653 0 -1 -23020
box 0 -20 400 440
use unit_Cap  unit_Cap_2242
timestamp 1756801411
transform 1 0 3197 0 -1 -22518
box 0 -20 400 440
use unit_Cap  unit_Cap_2243
timestamp 1756801411
transform 1 0 3653 0 -1 -22518
box 0 -20 400 440
<< labels >>
flabel metal2 15666 -14777 15716 -14714 0 FreeSans 160 0 0 0 C3
port 5 nsew
flabel metal2 15649 -15273 15719 -15208 0 FreeSans 160 0 0 0 C1
port 3 nsew
flabel metal2 15646 -15786 15714 -15726 0 FreeSans 160 0 0 0 C0
port 2 nsew
flabel metal2 15650 -16288 15718 -16228 0 FreeSans 160 0 0 0 C0_dummy
port 1 nsew
flabel metal2 15649 -16781 15714 -16717 0 FreeSans 160 0 0 0 C2
port 4 nsew
flabel metal2 15645 -17278 15717 -17215 0 FreeSans 160 0 0 0 C4
port 6 nsew
flabel metal2 15646 -18288 15713 -18224 0 FreeSans 160 0 0 0 C5
port 7 nsew
flabel metal2 15643 -18786 15715 -18725 0 FreeSans 160 0 0 0 C6
port 8 nsew
flabel metal2 15647 -19776 15715 -19713 0 FreeSans 160 0 0 0 C7
port 9 nsew
flabel metal2 15635 -21286 15717 -21221 0 FreeSans 160 0 0 0 C8
port 10 nsew
flabel metal2 15633 -23761 15717 -23699 0 FreeSans 160 0 0 0 C9
port 11 nsew
flabel metal2 15642 -26755 15716 -26692 0 FreeSans 160 0 0 0 C10
port 12 nsew
flabel metal5 14340 540 14530 610 0 FreeSans 320 0 0 0 Ctop
port 13 nsew
flabel metal5 15110 540 15460 630 0 FreeSans 320 0 0 0 VSS
port 14 nsew
<< end >>
