magic
tech gf180mcuD
magscale 1 10
timestamp 1757840551
<< pwell >>
rect -1736 -2658 1736 2658
<< psubdiff >>
rect -1712 2562 1712 2634
rect -1712 2518 -1640 2562
rect -1712 -2518 -1699 2518
rect -1653 -2518 -1640 2518
rect 1640 2518 1712 2562
rect -1712 -2562 -1640 -2518
rect 1640 -2518 1653 2518
rect 1699 -2518 1712 2518
rect 1640 -2562 1712 -2518
rect -1712 -2634 1712 -2562
<< psubdiffcont >>
rect -1699 -2518 -1653 2518
rect 1653 -2518 1699 2518
<< polysilicon >>
rect -1500 2409 -1300 2422
rect -1500 2363 -1487 2409
rect -1313 2363 -1300 2409
rect -1500 2300 -1300 2363
rect -1500 -2363 -1300 -2300
rect -1500 -2409 -1487 -2363
rect -1313 -2409 -1300 -2363
rect -1500 -2422 -1300 -2409
rect -1220 2409 -1020 2422
rect -1220 2363 -1207 2409
rect -1033 2363 -1020 2409
rect -1220 2300 -1020 2363
rect -1220 -2363 -1020 -2300
rect -1220 -2409 -1207 -2363
rect -1033 -2409 -1020 -2363
rect -1220 -2422 -1020 -2409
rect -940 2409 -740 2422
rect -940 2363 -927 2409
rect -753 2363 -740 2409
rect -940 2300 -740 2363
rect -940 -2363 -740 -2300
rect -940 -2409 -927 -2363
rect -753 -2409 -740 -2363
rect -940 -2422 -740 -2409
rect -660 2409 -460 2422
rect -660 2363 -647 2409
rect -473 2363 -460 2409
rect -660 2300 -460 2363
rect -660 -2363 -460 -2300
rect -660 -2409 -647 -2363
rect -473 -2409 -460 -2363
rect -660 -2422 -460 -2409
rect -380 2409 -180 2422
rect -380 2363 -367 2409
rect -193 2363 -180 2409
rect -380 2300 -180 2363
rect -380 -2363 -180 -2300
rect -380 -2409 -367 -2363
rect -193 -2409 -180 -2363
rect -380 -2422 -180 -2409
rect -100 2409 100 2422
rect -100 2363 -87 2409
rect 87 2363 100 2409
rect -100 2300 100 2363
rect -100 -2363 100 -2300
rect -100 -2409 -87 -2363
rect 87 -2409 100 -2363
rect -100 -2422 100 -2409
rect 180 2409 380 2422
rect 180 2363 193 2409
rect 367 2363 380 2409
rect 180 2300 380 2363
rect 180 -2363 380 -2300
rect 180 -2409 193 -2363
rect 367 -2409 380 -2363
rect 180 -2422 380 -2409
rect 460 2409 660 2422
rect 460 2363 473 2409
rect 647 2363 660 2409
rect 460 2300 660 2363
rect 460 -2363 660 -2300
rect 460 -2409 473 -2363
rect 647 -2409 660 -2363
rect 460 -2422 660 -2409
rect 740 2409 940 2422
rect 740 2363 753 2409
rect 927 2363 940 2409
rect 740 2300 940 2363
rect 740 -2363 940 -2300
rect 740 -2409 753 -2363
rect 927 -2409 940 -2363
rect 740 -2422 940 -2409
rect 1020 2409 1220 2422
rect 1020 2363 1033 2409
rect 1207 2363 1220 2409
rect 1020 2300 1220 2363
rect 1020 -2363 1220 -2300
rect 1020 -2409 1033 -2363
rect 1207 -2409 1220 -2363
rect 1020 -2422 1220 -2409
rect 1300 2409 1500 2422
rect 1300 2363 1313 2409
rect 1487 2363 1500 2409
rect 1300 2300 1500 2363
rect 1300 -2363 1500 -2300
rect 1300 -2409 1313 -2363
rect 1487 -2409 1500 -2363
rect 1300 -2422 1500 -2409
<< polycontact >>
rect -1487 2363 -1313 2409
rect -1487 -2409 -1313 -2363
rect -1207 2363 -1033 2409
rect -1207 -2409 -1033 -2363
rect -927 2363 -753 2409
rect -927 -2409 -753 -2363
rect -647 2363 -473 2409
rect -647 -2409 -473 -2363
rect -367 2363 -193 2409
rect -367 -2409 -193 -2363
rect -87 2363 87 2409
rect -87 -2409 87 -2363
rect 193 2363 367 2409
rect 193 -2409 367 -2363
rect 473 2363 647 2409
rect 473 -2409 647 -2363
rect 753 2363 927 2409
rect 753 -2409 927 -2363
rect 1033 2363 1207 2409
rect 1033 -2409 1207 -2363
rect 1313 2363 1487 2409
rect 1313 -2409 1487 -2363
<< nhighres >>
rect -1500 -2300 -1300 2300
rect -1220 -2300 -1020 2300
rect -940 -2300 -740 2300
rect -660 -2300 -460 2300
rect -380 -2300 -180 2300
rect -100 -2300 100 2300
rect 180 -2300 380 2300
rect 460 -2300 660 2300
rect 740 -2300 940 2300
rect 1020 -2300 1220 2300
rect 1300 -2300 1500 2300
<< metal1 >>
rect -1699 2575 1699 2621
rect -1699 2518 -1653 2575
rect 1653 2518 1699 2575
rect -1498 2363 -1487 2409
rect -1313 2363 -1302 2409
rect -1218 2363 -1207 2409
rect -1033 2363 -1022 2409
rect -938 2363 -927 2409
rect -753 2363 -742 2409
rect -658 2363 -647 2409
rect -473 2363 -462 2409
rect -378 2363 -367 2409
rect -193 2363 -182 2409
rect -98 2363 -87 2409
rect 87 2363 98 2409
rect 182 2363 193 2409
rect 367 2363 378 2409
rect 462 2363 473 2409
rect 647 2363 658 2409
rect 742 2363 753 2409
rect 927 2363 938 2409
rect 1022 2363 1033 2409
rect 1207 2363 1218 2409
rect 1302 2363 1313 2409
rect 1487 2363 1498 2409
rect -1498 -2409 -1487 -2363
rect -1313 -2409 -1302 -2363
rect -1218 -2409 -1207 -2363
rect -1033 -2409 -1022 -2363
rect -938 -2409 -927 -2363
rect -753 -2409 -742 -2363
rect -658 -2409 -647 -2363
rect -473 -2409 -462 -2363
rect -378 -2409 -367 -2363
rect -193 -2409 -182 -2363
rect -98 -2409 -87 -2363
rect 87 -2409 98 -2363
rect 182 -2409 193 -2363
rect 367 -2409 378 -2363
rect 462 -2409 473 -2363
rect 647 -2409 658 -2363
rect 742 -2409 753 -2363
rect 927 -2409 938 -2363
rect 1022 -2409 1033 -2363
rect 1207 -2409 1218 -2363
rect 1302 -2409 1313 -2363
rect 1487 -2409 1498 -2363
rect -1699 -2575 -1653 -2518
rect 1653 -2575 1699 -2518
rect -1699 -2621 1699 -2575
<< properties >>
string FIXED_BBOX -1676 -2598 1676 2598
string gencell ppolyf_u_1k
string library gf180mcu
string parameters w 1.000 l 23.000 m 1 nx 11 wmin 1.000 lmin 1.000 class resistor rho 1000 val 23.0k dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 1 grc 1 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 1 compatible {ppolyf_u_1k ppolyf_u_1k_6p0}
<< end >>
