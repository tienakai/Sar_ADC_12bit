magic
tech gf180mcuD
magscale 1 10
timestamp 1757239713
<< nwell >>
rect -442 -930 442 930
<< pmos >>
rect -268 -800 -212 800
rect -108 -800 -52 800
rect 52 -800 108 800
rect 212 -800 268 800
<< pdiff >>
rect -356 787 -268 800
rect -356 -787 -343 787
rect -297 -787 -268 787
rect -356 -800 -268 -787
rect -212 787 -108 800
rect -212 -787 -183 787
rect -137 -787 -108 787
rect -212 -800 -108 -787
rect -52 787 52 800
rect -52 -787 -23 787
rect 23 -787 52 787
rect -52 -800 52 -787
rect 108 787 212 800
rect 108 -787 137 787
rect 183 -787 212 787
rect 108 -800 212 -787
rect 268 787 356 800
rect 268 -787 297 787
rect 343 -787 356 787
rect 268 -800 356 -787
<< pdiffc >>
rect -343 -787 -297 787
rect -183 -787 -137 787
rect -23 -787 23 787
rect 137 -787 183 787
rect 297 -787 343 787
<< polysilicon >>
rect -268 800 -212 844
rect -108 800 -52 844
rect 52 800 108 844
rect 212 800 268 844
rect -268 -844 -212 -800
rect -108 -844 -52 -800
rect 52 -844 108 -800
rect 212 -844 268 -800
<< metal1 >>
rect -343 787 -297 798
rect -343 -798 -297 -787
rect -183 787 -137 798
rect -183 -798 -137 -787
rect -23 787 23 798
rect -23 -798 23 -787
rect 137 787 183 798
rect 137 -798 183 -787
rect 297 787 343 798
rect 297 -798 343 -787
<< properties >>
string gencell pfet_03v3
string library gf180mcu
string parameters w 8 l 0.280 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {pfet_03v3 pfet_06v0}
<< end >>
