magic
tech gf180mcuD
magscale 1 10
timestamp 1757414845
<< nwell >>
rect -212 -416 212 416
<< pwell >>
rect -374 416 374 536
rect -374 -416 -212 416
rect 212 -416 374 416
rect -374 -536 374 -416
<< psubdiff >>
rect -350 440 350 512
rect -350 396 -278 440
rect -350 -396 -337 396
rect -291 -396 -278 396
rect 278 396 350 440
rect -350 -440 -278 -396
rect 278 -396 291 396
rect 337 -396 350 396
rect 278 -440 350 -396
rect -350 -512 350 -440
<< nsubdiff >>
rect -188 287 -100 300
rect -188 -287 -175 287
rect -129 -287 -100 287
rect -188 -300 -100 -287
rect 100 287 188 300
rect 100 -287 129 287
rect 175 -287 188 287
rect 100 -300 188 -287
<< psubdiffcont >>
rect -337 -396 -291 396
rect 291 -396 337 396
<< nsubdiffcont >>
rect -175 -287 -129 287
rect 129 -287 175 287
<< nvaractor >>
rect -100 -300 100 300
<< polysilicon >>
rect -100 379 100 392
rect -100 333 -87 379
rect 87 333 100 379
rect -100 300 100 333
rect -100 -333 100 -300
rect -100 -379 -87 -333
rect 87 -379 100 -333
rect -100 -392 100 -379
<< polycontact >>
rect -87 333 87 379
rect -87 -379 87 -333
<< metal1 >>
rect -337 453 337 499
rect -337 396 -291 453
rect 291 396 337 453
rect -98 333 -87 379
rect 87 333 98 379
rect -175 287 -129 298
rect -175 -298 -129 -287
rect 129 287 175 298
rect 129 -298 175 -287
rect -98 -379 -87 -333
rect 87 -379 98 -333
rect -337 -453 -291 -396
rect 291 -453 337 -396
rect -337 -499 337 -453
<< properties >>
string FIXED_BBOX -314 -476 314 476
string gencell nmoscap_3p3
string library gf180mcu
string parameters w 3.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {nmoscap_3p3 nmoscap_6p0}
<< end >>
