magic
tech gf180mcuD
magscale 1 10
timestamp 1757859342
<< nwell >>
rect -394 412 3954 823
rect -2258 -98 3954 412
rect -2080 -115 3954 -98
rect -2081 -119 3954 -115
rect -2081 -141 4292 -119
rect -2081 -240 193 -141
rect 3721 -185 4292 -141
rect 4813 -182 5384 -116
rect -1715 -484 -1642 -463
rect -97 -591 25 -323
<< pwell >>
rect -2740 510 -514 909
rect 831 -608 2646 -290
rect 831 -621 2854 -608
rect 803 -906 2854 -621
rect -2079 -964 233 -909
rect 723 -964 2854 -906
rect 3431 -964 3617 -874
rect 3778 -964 4423 -903
rect -2079 -973 4423 -964
rect 4747 -966 5392 -896
rect -2079 -1029 4004 -973
rect -242 -1213 4004 -1029
rect -242 -2286 4011 -1213
rect -235 -2535 4011 -2286
<< nmos >>
rect 1150 -760 1206 -360
rect 2241 -759 2297 -359
rect 262 -1590 318 -1190
rect 613 -1590 669 -1190
rect 1239 -1590 1295 -1190
rect 2139 -1591 2195 -1191
rect 3010 -1990 3066 -1190
rect 3360 -1990 3416 -1190
<< pmos >>
rect 0 0 56 400
rect 205 0 261 400
rect 816 92 872 492
rect 1021 92 1077 492
rect 1199 92 1255 492
rect 1404 92 1460 492
rect 2055 92 2111 492
rect 2260 92 2316 492
rect 2438 92 2494 492
rect 2643 92 2699 492
rect 3316 0 3372 400
rect 3521 0 3577 400
<< ndiff >>
rect 1059 -390 1150 -360
rect 1059 -730 1075 -390
rect 1121 -730 1150 -390
rect 1059 -760 1150 -730
rect 1206 -390 1297 -360
rect 1206 -730 1237 -390
rect 1283 -730 1297 -390
rect 1206 -760 1297 -730
rect 2150 -392 2241 -359
rect 2150 -729 2166 -392
rect 2212 -729 2241 -392
rect 2150 -759 2241 -729
rect 2297 -389 2388 -359
rect 2297 -729 2328 -389
rect 2374 -729 2388 -389
rect 2297 -759 2388 -729
rect 153 -1221 262 -1190
rect 153 -1559 184 -1221
rect 233 -1559 262 -1221
rect 153 -1590 262 -1559
rect 318 -1221 427 -1190
rect 318 -1559 349 -1221
rect 398 -1559 427 -1221
rect 318 -1590 427 -1559
rect 504 -1221 613 -1190
rect 504 -1559 535 -1221
rect 584 -1559 613 -1221
rect 504 -1590 613 -1559
rect 669 -1221 778 -1190
rect 669 -1559 700 -1221
rect 749 -1559 778 -1221
rect 669 -1590 778 -1559
rect 1129 -1222 1239 -1190
rect 1129 -1560 1160 -1222
rect 1209 -1560 1239 -1222
rect 1129 -1590 1239 -1560
rect 1295 -1221 1390 -1190
rect 1295 -1560 1329 -1221
rect 1375 -1560 1390 -1221
rect 1295 -1590 1390 -1560
rect 1129 -1591 1210 -1590
rect 2029 -1223 2139 -1191
rect 2029 -1561 2060 -1223
rect 2109 -1561 2139 -1223
rect 2029 -1591 2139 -1561
rect 2195 -1222 2290 -1191
rect 2195 -1561 2229 -1222
rect 2275 -1561 2290 -1222
rect 2195 -1591 2290 -1561
rect 2029 -1592 2110 -1591
rect 2917 -1219 3010 -1190
rect 2917 -1969 2932 -1219
rect 2980 -1969 3010 -1219
rect 2917 -1990 3010 -1969
rect 3066 -1216 3160 -1190
rect 3066 -1970 3096 -1216
rect 3144 -1970 3160 -1216
rect 3066 -1990 3160 -1970
rect 3267 -1219 3360 -1190
rect 3267 -1969 3282 -1219
rect 3330 -1969 3360 -1219
rect 3267 -1990 3360 -1969
rect 3416 -1216 3510 -1190
rect 3416 -1970 3446 -1216
rect 3494 -1970 3510 -1216
rect 3416 -1990 3510 -1970
<< pdiff >>
rect -110 370 0 400
rect -110 30 -83 370
rect -37 30 0 370
rect -110 0 0 30
rect 56 370 205 400
rect 56 30 106 370
rect 155 30 205 370
rect 56 0 205 30
rect 261 370 360 400
rect 261 31 292 370
rect 339 31 360 370
rect 261 0 360 31
rect 717 461 816 492
rect 717 122 738 461
rect 785 122 816 461
rect 717 92 816 122
rect 872 462 1021 492
rect 872 122 922 462
rect 971 122 1021 462
rect 872 92 1021 122
rect 1077 462 1199 492
rect 1077 122 1114 462
rect 1160 122 1199 462
rect 1077 92 1199 122
rect 1255 462 1404 492
rect 1255 122 1305 462
rect 1354 122 1404 462
rect 1255 92 1404 122
rect 1460 462 1582 492
rect 1460 122 1497 462
rect 1543 122 1582 462
rect 1460 92 1582 122
rect 1956 461 2055 492
rect 1956 122 1977 461
rect 2024 122 2055 461
rect 1956 92 2055 122
rect 2111 462 2260 492
rect 2111 122 2161 462
rect 2210 122 2260 462
rect 2111 92 2260 122
rect 2316 462 2438 492
rect 2316 122 2353 462
rect 2399 122 2438 462
rect 2316 92 2438 122
rect 2494 462 2643 492
rect 2494 122 2544 462
rect 2593 122 2643 462
rect 2494 92 2643 122
rect 2699 462 2821 492
rect 2699 122 2736 462
rect 2782 122 2821 462
rect 2699 92 2821 122
rect 3206 370 3316 400
rect 3206 30 3233 370
rect 3279 30 3316 370
rect 3206 0 3316 30
rect 3372 370 3521 400
rect 3372 30 3422 370
rect 3471 30 3521 370
rect 3372 0 3521 30
rect 3577 370 3676 400
rect 3577 31 3608 370
rect 3655 31 3676 370
rect 3577 0 3676 31
<< mvpdiff >>
rect -1715 -484 -1642 -463
<< ndiffc >>
rect 1075 -730 1121 -390
rect 1237 -730 1283 -390
rect 2166 -729 2212 -392
rect 2328 -729 2374 -389
rect 184 -1559 233 -1221
rect 349 -1559 398 -1221
rect 535 -1559 584 -1221
rect 700 -1559 749 -1221
rect 1160 -1560 1209 -1222
rect 1329 -1560 1375 -1221
rect 2060 -1561 2109 -1223
rect 2229 -1561 2275 -1222
rect 2932 -1969 2980 -1219
rect 3096 -1970 3144 -1216
rect 3282 -1969 3330 -1219
rect 3446 -1970 3494 -1216
<< pdiffc >>
rect -83 30 -37 370
rect 106 30 155 370
rect 292 31 339 370
rect 738 122 785 461
rect 922 122 971 462
rect 1114 122 1160 462
rect 1305 122 1354 462
rect 1497 122 1543 462
rect 1977 122 2024 461
rect 2161 122 2210 462
rect 2353 122 2399 462
rect 2544 122 2593 462
rect 2736 122 2782 462
rect 3233 30 3279 370
rect 3422 30 3471 370
rect 3608 31 3655 370
<< psubdiff >>
rect -2599 806 -2166 833
rect -2599 730 -2569 806
rect -2280 730 -2166 806
rect -2599 712 -2166 730
rect 882 -394 983 -343
rect 1458 -326 1564 -324
rect 882 -819 899 -394
rect 967 -819 983 -394
rect 1458 -378 1582 -326
rect 882 -876 983 -819
rect 1458 -811 1473 -378
rect 1564 -811 1582 -378
rect 1458 -876 1582 -811
rect 1907 -361 2040 -329
rect 1907 -794 1932 -361
rect 2023 -794 2040 -361
rect 2481 -376 2586 -328
rect 1907 -876 2040 -794
rect 2481 -793 2497 -376
rect 2573 -793 2586 -376
rect 2481 -874 2586 -793
rect 2481 -876 2771 -874
rect 882 -892 2771 -876
rect 882 -893 2099 -892
rect 882 -906 1016 -893
rect 723 -981 1016 -906
rect 1373 -980 2099 -893
rect 2456 -980 2771 -892
rect 1373 -981 2771 -980
rect 723 -994 2771 -981
rect -109 -1192 77 -998
rect 723 -1024 1043 -994
rect 893 -1044 1043 -1024
rect -109 -1708 -68 -1192
rect 38 -1708 77 -1192
rect 893 -1514 921 -1044
rect 1028 -1514 1043 -1044
rect 1678 -1061 1828 -994
rect 893 -1581 1043 -1514
rect 1678 -1531 1706 -1061
rect 1813 -1531 1828 -1061
rect 2469 -997 2771 -994
rect 2469 -1061 2624 -997
rect -109 -1900 77 -1708
rect 1678 -1594 1828 -1531
rect 2469 -1531 2497 -1061
rect 2604 -1531 2624 -1061
rect 2469 -1600 2624 -1531
rect 2469 -1635 2623 -1600
rect -109 -1901 102 -1900
rect 2468 -1901 2623 -1635
rect -109 -1925 2623 -1901
rect -109 -1931 1468 -1925
rect -109 -2063 299 -1931
rect 928 -2057 1468 -1931
rect 2097 -2057 2623 -1925
rect 3671 -1316 3824 -986
rect 3671 -1904 3702 -1316
rect 3786 -1904 3824 -1316
rect 928 -2063 2623 -2057
rect -109 -2091 2623 -2063
rect -109 -2094 2348 -2091
rect 2468 -2236 2623 -2091
rect 3671 -2236 3824 -1904
rect 2468 -2271 3825 -2236
rect 2468 -2365 2805 -2271
rect 3466 -2365 3825 -2271
rect 2468 -2391 3825 -2365
<< nsubdiff >>
rect -258 770 -174 771
rect 524 770 2218 771
rect -364 748 3922 770
rect -364 742 846 748
rect -364 675 -212 742
rect 406 675 846 742
rect -364 668 846 675
rect 1434 744 3922 748
rect 1434 676 2082 744
rect 2632 742 3922 744
rect 2632 676 3312 742
rect 1434 668 3312 676
rect -364 660 3312 668
rect 3827 660 3922 742
rect -364 640 3922 660
rect -364 530 -246 640
rect -364 17 -338 530
rect -279 17 -246 530
rect 470 534 588 640
rect 1042 639 3922 640
rect -364 -71 -246 17
rect 470 21 495 534
rect 554 21 588 534
rect 1704 533 1822 639
rect 2208 638 2832 639
rect 2956 544 3074 639
rect 3599 637 3922 639
rect 470 -71 588 21
rect 1704 20 1729 533
rect 1788 20 1822 533
rect 1704 -72 1822 20
rect 2956 31 2981 544
rect 3040 31 3074 544
rect 3805 547 3922 637
rect 2956 -61 3074 31
rect 3805 34 3830 547
rect 3889 34 3922 547
rect 3805 -58 3922 34
<< psubdiffcont >>
rect -2569 730 -2280 806
rect 899 -819 967 -394
rect 1473 -811 1564 -378
rect 1932 -794 2023 -361
rect 2497 -793 2573 -376
rect 1016 -981 1373 -893
rect 2099 -980 2456 -892
rect -68 -1708 38 -1192
rect 921 -1514 1028 -1044
rect 1706 -1531 1813 -1061
rect 2497 -1531 2604 -1061
rect 299 -2063 928 -1931
rect 1468 -2057 2097 -1925
rect 3702 -1904 3786 -1316
rect 2805 -2365 3466 -2271
<< nsubdiffcont >>
rect -212 675 406 742
rect 846 668 1434 748
rect 2082 676 2632 744
rect 3312 660 3827 742
rect -338 17 -279 530
rect 495 21 554 534
rect 1729 20 1788 533
rect 2981 31 3040 544
rect 3830 34 3889 547
<< polysilicon >>
rect -60 520 56 542
rect -60 460 -43 520
rect 40 460 56 520
rect -60 443 56 460
rect 204 524 320 544
rect 204 464 222 524
rect 305 464 320 524
rect 204 445 320 464
rect 0 400 56 443
rect 205 400 261 445
rect 816 492 872 542
rect 1021 492 1077 542
rect 1199 492 1255 542
rect 1404 492 1460 542
rect 0 -50 56 0
rect 205 -50 261 0
rect 816 42 872 92
rect 1021 42 1077 92
rect 816 39 1077 42
rect 1199 42 1255 92
rect 1404 42 1460 92
rect 1199 39 1460 42
rect 816 25 1460 39
rect 816 -29 1139 25
rect 1230 -29 1460 25
rect 816 -49 1460 -29
rect 2055 492 2111 542
rect 2260 492 2316 542
rect 2438 492 2494 542
rect 2643 492 2699 542
rect 1055 -50 1238 -49
rect 2055 42 2111 92
rect 2260 42 2316 92
rect 2055 39 2316 42
rect 2438 42 2494 92
rect 2643 42 2699 92
rect 2438 39 2699 42
rect 2055 26 2699 39
rect 2055 -44 2218 26
rect 2341 -44 2699 26
rect 2055 -49 2699 -44
rect 2056 -60 2699 -49
rect 3257 517 3372 542
rect 3257 461 3272 517
rect 3353 461 3372 517
rect 3257 443 3372 461
rect 3316 400 3372 443
rect 3520 521 3635 541
rect 3520 465 3534 521
rect 3615 465 3635 521
rect 3520 442 3635 465
rect 3521 400 3577 442
rect 3316 -50 3372 0
rect 3521 -50 3577 0
rect 1117 -251 1244 -236
rect 1117 -302 1147 -251
rect 1211 -302 1244 -251
rect 1117 -316 1244 -302
rect 2208 -250 2335 -235
rect 2208 -301 2238 -250
rect 2302 -301 2335 -250
rect 2208 -315 2335 -301
rect 2214 -316 2328 -315
rect 1123 -317 1237 -316
rect 1150 -360 1206 -317
rect 1150 -810 1206 -760
rect 2241 -359 2297 -316
rect 2241 -809 2297 -759
rect 262 -1190 318 -1140
rect 613 -1190 669 -1140
rect 1214 -1089 1330 -1073
rect 1214 -1138 1242 -1089
rect 1300 -1138 1330 -1089
rect 1214 -1151 1330 -1138
rect 1239 -1190 1295 -1151
rect 2114 -1090 2230 -1074
rect 2114 -1139 2142 -1090
rect 2200 -1139 2230 -1090
rect 2114 -1152 2230 -1139
rect 2139 -1191 2195 -1152
rect 262 -1638 318 -1590
rect 613 -1635 669 -1590
rect 259 -1651 360 -1638
rect 259 -1707 277 -1651
rect 339 -1707 360 -1651
rect 259 -1720 360 -1707
rect 568 -1649 670 -1635
rect 1239 -1640 1295 -1590
rect 3010 -1190 3066 -1140
rect 3360 -1190 3416 -1140
rect 2139 -1641 2195 -1591
rect 568 -1705 589 -1649
rect 655 -1705 670 -1649
rect 568 -1720 670 -1705
rect 273 -1721 360 -1720
rect 3010 -2038 3066 -1990
rect 3009 -2050 3066 -2038
rect 3360 -2049 3416 -1990
rect 3009 -2068 3130 -2050
rect 3009 -2125 3039 -2068
rect 3101 -2125 3130 -2068
rect 3009 -2144 3130 -2125
rect 3259 -2067 3416 -2049
rect 3259 -2124 3310 -2067
rect 3372 -2124 3416 -2067
rect 3259 -2142 3416 -2124
rect 3259 -2143 3380 -2142
<< polycontact >>
rect -43 460 40 520
rect 222 464 305 524
rect 1139 -29 1230 25
rect 2218 -44 2341 26
rect 3272 461 3353 517
rect 3534 465 3615 521
rect 1147 -302 1211 -251
rect 2238 -301 2302 -250
rect 1242 -1138 1300 -1089
rect 2142 -1139 2200 -1090
rect 277 -1707 339 -1651
rect 589 -1705 655 -1649
rect 3039 -2125 3101 -2068
rect 3310 -2124 3372 -2067
<< metal1 >>
rect -2600 808 -2166 833
rect -2600 729 -2570 808
rect -2280 729 -2166 808
rect 524 770 2218 771
rect -364 748 3922 770
rect -364 742 846 748
rect -2600 712 -2166 729
rect -364 674 -212 742
rect 406 733 846 742
rect 1434 744 3922 748
rect 1434 733 2082 744
rect 406 674 845 733
rect -364 667 845 674
rect 1463 676 2082 733
rect 2632 742 3922 744
rect 2632 676 3312 742
rect 1463 667 3312 676
rect -364 660 3312 667
rect 3827 660 3922 742
rect -364 640 3922 660
rect -364 531 -246 640
rect -364 17 -340 531
rect -277 17 -246 531
rect -60 520 56 542
rect -60 460 -43 520
rect 40 460 56 520
rect -60 443 56 460
rect 204 524 320 544
rect 204 464 222 524
rect 305 464 320 524
rect 204 445 320 464
rect 470 534 588 640
rect 1042 639 3922 640
rect -92 370 -24 381
rect -92 368 -83 370
rect -37 368 -24 370
rect -92 31 -84 368
rect -32 31 -24 368
rect -92 30 -83 31
rect -37 30 -24 31
rect -92 20 -24 30
rect 90 370 170 381
rect 90 33 103 370
rect 90 30 106 33
rect 155 30 170 370
rect 90 20 170 30
rect 277 370 344 381
rect 277 369 292 370
rect 277 32 287 369
rect 277 31 292 32
rect 339 31 344 370
rect 277 20 344 31
rect 470 20 495 534
rect 558 20 588 534
rect 1704 533 1822 639
rect 2208 638 2832 639
rect 733 461 800 472
rect 733 122 738 461
rect 785 460 800 461
rect 790 123 800 460
rect 785 122 800 123
rect 733 111 800 122
rect 907 462 987 472
rect 907 122 922 462
rect 971 459 987 462
rect 974 122 987 459
rect 907 111 987 122
rect 1101 462 1169 472
rect 1101 461 1114 462
rect 1160 461 1169 462
rect 1101 124 1109 461
rect 1161 124 1169 461
rect 1101 122 1114 124
rect 1160 122 1169 124
rect 1101 111 1169 122
rect 1290 462 1370 472
rect 1290 122 1305 462
rect 1354 459 1370 462
rect 1357 122 1370 459
rect 1290 111 1370 122
rect 1484 462 1552 472
rect 1484 461 1497 462
rect 1543 461 1552 462
rect 1484 124 1492 461
rect 1544 124 1552 461
rect 1484 122 1497 124
rect 1543 122 1552 124
rect 1484 111 1552 122
rect -364 -71 -246 17
rect 470 -70 588 20
rect 1114 25 1252 38
rect 1114 -29 1139 25
rect 1230 -29 1252 25
rect 1114 -47 1252 -29
rect 1704 19 1729 533
rect 1792 19 1822 533
rect 2956 544 3074 639
rect 3599 637 3922 639
rect 1972 461 2039 472
rect 1972 122 1977 461
rect 2024 460 2039 461
rect 2029 123 2039 460
rect 2024 122 2039 123
rect 1972 111 2039 122
rect 2146 462 2226 472
rect 2146 122 2161 462
rect 2210 459 2226 462
rect 2213 122 2226 459
rect 2146 111 2226 122
rect 2340 462 2408 472
rect 2340 461 2353 462
rect 2399 461 2408 462
rect 2340 124 2348 461
rect 2400 124 2408 461
rect 2340 122 2353 124
rect 2399 122 2408 124
rect 2340 111 2408 122
rect 2529 462 2609 472
rect 2529 122 2544 462
rect 2593 459 2609 462
rect 2596 122 2609 459
rect 2529 111 2609 122
rect 2723 462 2791 472
rect 2723 461 2736 462
rect 2782 461 2791 462
rect 2723 124 2731 461
rect 2783 124 2791 461
rect 2723 122 2736 124
rect 2782 122 2791 124
rect 2723 111 2791 122
rect 1704 -71 1822 19
rect 2203 26 2360 37
rect 2203 -44 2218 26
rect 2341 -44 2360 26
rect 2203 -52 2360 -44
rect 2956 30 2981 544
rect 3044 30 3074 544
rect 3805 547 3922 637
rect 3257 517 3372 542
rect 3257 461 3272 517
rect 3353 461 3372 517
rect 3257 443 3372 461
rect 3520 521 3635 541
rect 3520 465 3534 521
rect 3615 465 3635 521
rect 3520 442 3635 465
rect 2956 -90 3074 30
rect 3224 370 3292 381
rect 3224 368 3233 370
rect 3279 368 3292 370
rect 3224 31 3232 368
rect 3284 31 3292 368
rect 3224 30 3233 31
rect 3279 30 3292 31
rect 3224 20 3292 30
rect 3406 370 3486 381
rect 3406 33 3419 370
rect 3406 30 3422 33
rect 3471 30 3486 370
rect 3406 20 3486 30
rect 3593 370 3660 381
rect 3593 369 3608 370
rect 3593 32 3603 369
rect 3593 31 3608 32
rect 3655 31 3660 370
rect 3593 20 3660 31
rect 3805 33 3830 547
rect 3893 33 3922 547
rect 3805 -90 3922 33
rect 2958 -95 3073 -90
rect 3805 -91 3921 -90
rect 3807 -96 3921 -91
rect 1117 -249 1244 -236
rect 1117 -302 1147 -249
rect 1211 -302 1244 -249
rect 1117 -316 1244 -302
rect 2208 -248 2335 -235
rect 2208 -301 2238 -248
rect 2302 -301 2335 -248
rect 2208 -315 2335 -301
rect 2214 -316 2328 -315
rect 1123 -317 1237 -316
rect 1458 -326 1564 -324
rect 882 -394 983 -343
rect 1458 -378 1582 -326
rect 882 -819 899 -394
rect 967 -819 983 -394
rect 1068 -390 1129 -378
rect 1068 -730 1075 -390
rect 1121 -393 1129 -390
rect 1127 -728 1129 -393
rect 1121 -730 1129 -728
rect 1068 -740 1129 -730
rect 1229 -390 1290 -378
rect 1229 -392 1237 -390
rect 1283 -392 1290 -390
rect 1229 -727 1234 -392
rect 1286 -727 1290 -392
rect 1229 -730 1237 -727
rect 1283 -730 1290 -727
rect 1229 -740 1290 -730
rect 882 -876 983 -819
rect 1458 -811 1473 -378
rect 1564 -811 1582 -378
rect 1458 -876 1582 -811
rect 1907 -361 2040 -329
rect 1907 -794 1932 -361
rect 2023 -794 2040 -361
rect 2158 -392 2229 -374
rect 2481 -376 2586 -328
rect 2158 -729 2166 -392
rect 2212 -393 2229 -392
rect 2218 -515 2229 -393
rect 2320 -389 2381 -377
rect 2320 -391 2328 -389
rect 2374 -391 2381 -389
rect 2218 -727 2230 -515
rect 2212 -729 2230 -727
rect 2158 -740 2230 -729
rect 2320 -726 2325 -391
rect 2377 -726 2381 -391
rect 2320 -729 2328 -726
rect 2374 -729 2381 -726
rect 2320 -739 2381 -729
rect 1907 -876 2040 -794
rect 2481 -793 2497 -376
rect 2573 -793 2586 -376
rect 2481 -874 2586 -793
rect 2481 -876 2771 -874
rect 882 -888 2771 -876
rect 882 -906 1016 -888
rect -2079 -928 233 -909
rect -2079 -935 161 -928
rect -2079 -1003 -1627 -935
rect -1089 -939 161 -935
rect -1089 -1003 -739 -939
rect -2079 -1007 -739 -1003
rect -201 -995 161 -939
rect 723 -981 1016 -906
rect 1376 -980 2088 -888
rect 2448 -892 2771 -888
rect 2456 -980 2771 -892
rect 1373 -981 2771 -980
rect 723 -994 2771 -981
rect 3431 -994 3617 -874
rect -201 -1007 233 -995
rect -2079 -1029 233 -1007
rect 723 -1024 1043 -994
rect -109 -1192 77 -1029
rect -109 -1708 -68 -1192
rect 38 -1708 77 -1192
rect 893 -1044 1043 -1024
rect 175 -1221 242 -1208
rect 175 -1229 184 -1221
rect 233 -1229 242 -1221
rect 175 -1552 181 -1229
rect 234 -1552 242 -1229
rect 175 -1559 184 -1552
rect 233 -1559 242 -1552
rect 175 -1570 242 -1559
rect 340 -1221 407 -1208
rect 340 -1229 349 -1221
rect 398 -1229 407 -1221
rect 340 -1552 346 -1229
rect 399 -1552 407 -1229
rect 340 -1559 349 -1552
rect 398 -1559 407 -1552
rect 340 -1570 407 -1559
rect 526 -1221 593 -1208
rect 526 -1229 535 -1221
rect 584 -1229 593 -1221
rect 526 -1552 532 -1229
rect 585 -1552 593 -1229
rect 526 -1559 535 -1552
rect 584 -1559 593 -1552
rect 526 -1570 593 -1559
rect 691 -1221 758 -1208
rect 691 -1229 700 -1221
rect 749 -1229 758 -1221
rect 691 -1552 697 -1229
rect 750 -1552 758 -1229
rect 691 -1559 700 -1552
rect 749 -1559 758 -1552
rect 691 -1570 758 -1559
rect 893 -1514 921 -1044
rect 1028 -1514 1043 -1044
rect 1678 -1061 1828 -994
rect 1214 -1087 1330 -1073
rect 1214 -1139 1241 -1087
rect 1306 -1139 1330 -1087
rect 1214 -1151 1330 -1139
rect 893 -1581 1043 -1514
rect 1151 -1222 1218 -1209
rect 1151 -1230 1160 -1222
rect 1209 -1230 1218 -1222
rect 1151 -1553 1157 -1230
rect 1210 -1553 1218 -1230
rect 1151 -1560 1160 -1553
rect 1209 -1560 1218 -1553
rect 1151 -1571 1218 -1560
rect 1313 -1221 1380 -1209
rect 1313 -1229 1329 -1221
rect 1313 -1552 1322 -1229
rect 1313 -1560 1329 -1552
rect 1375 -1560 1380 -1221
rect 1313 -1571 1380 -1560
rect 1678 -1531 1706 -1061
rect 1813 -1531 1828 -1061
rect 2469 -997 2771 -994
rect 2469 -1061 2624 -997
rect 2114 -1086 2230 -1074
rect 2114 -1139 2142 -1086
rect 2201 -1139 2230 -1086
rect 2114 -1152 2230 -1139
rect 1678 -1594 1828 -1531
rect 2051 -1223 2118 -1210
rect 2213 -1220 2280 -1210
rect 2051 -1231 2060 -1223
rect 2109 -1231 2118 -1223
rect 2051 -1554 2057 -1231
rect 2110 -1554 2118 -1231
rect 2211 -1222 2280 -1220
rect 2211 -1226 2229 -1222
rect 2211 -1349 2222 -1226
rect 2051 -1561 2060 -1554
rect 2109 -1561 2118 -1554
rect 2051 -1572 2118 -1561
rect 2213 -1553 2222 -1349
rect 2213 -1561 2229 -1553
rect 2275 -1561 2280 -1222
rect 2213 -1572 2280 -1561
rect 2469 -1531 2497 -1061
rect 2604 -1531 2624 -1061
rect 2469 -1600 2624 -1531
rect 2927 -1219 2991 -1206
rect 2469 -1635 2623 -1600
rect -109 -1900 77 -1708
rect 259 -1651 360 -1640
rect 259 -1707 277 -1651
rect 339 -1707 360 -1651
rect 259 -1720 360 -1707
rect 568 -1649 670 -1640
rect 568 -1705 589 -1649
rect 655 -1705 670 -1649
rect 568 -1720 670 -1705
rect -109 -1901 102 -1900
rect 2468 -1901 2623 -1635
rect -109 -1925 2623 -1901
rect -109 -1931 1468 -1925
rect -109 -2063 299 -1931
rect 928 -2057 1468 -1931
rect 2097 -2057 2623 -1925
rect 2927 -1969 2932 -1219
rect 2980 -1233 2991 -1219
rect 2985 -1953 2991 -1233
rect 2980 -1969 2991 -1953
rect 2927 -1980 2991 -1969
rect 3088 -1216 3152 -1206
rect 3088 -1238 3096 -1216
rect 3144 -1238 3152 -1216
rect 3088 -1958 3095 -1238
rect 3147 -1958 3152 -1238
rect 3088 -1970 3096 -1958
rect 3144 -1970 3152 -1958
rect 3088 -1980 3152 -1970
rect 3277 -1219 3341 -1206
rect 3277 -1969 3282 -1219
rect 3330 -1233 3341 -1219
rect 3335 -1953 3341 -1233
rect 3330 -1969 3341 -1953
rect 3277 -1980 3341 -1969
rect 3438 -1216 3502 -1206
rect 3438 -1238 3446 -1216
rect 3494 -1238 3502 -1216
rect 3438 -1958 3445 -1238
rect 3497 -1958 3502 -1238
rect 3438 -1970 3446 -1958
rect 3494 -1970 3502 -1958
rect 3438 -1980 3502 -1970
rect 3671 -1316 3824 -986
rect 3671 -1904 3702 -1316
rect 3786 -1904 3824 -1316
rect 928 -2063 2623 -2057
rect -109 -2091 2623 -2063
rect -109 -2094 2348 -2091
rect 2468 -2236 2623 -2091
rect 3009 -2067 3416 -2050
rect 3009 -2068 3310 -2067
rect 3009 -2125 3039 -2068
rect 3101 -2124 3310 -2068
rect 3372 -2124 3416 -2067
rect 3101 -2125 3416 -2124
rect 3009 -2145 3416 -2125
rect 3671 -2236 3824 -1904
rect 2468 -2271 3825 -2236
rect 2468 -2365 2805 -2271
rect 3466 -2365 3825 -2271
rect 2468 -2391 3825 -2365
<< via1 >>
rect -2570 806 -2280 808
rect -2570 730 -2569 806
rect -2569 730 -2280 806
rect -2570 729 -2280 730
rect -1891 730 -1560 812
rect -1134 734 -803 816
rect -212 675 406 740
rect -212 674 406 675
rect 845 668 846 733
rect 846 668 1434 733
rect 1434 668 1463 733
rect 2082 676 2632 744
rect 845 667 1463 668
rect 3312 660 3827 742
rect -2004 358 -1792 424
rect -1054 243 -994 296
rect -1973 -52 -1544 23
rect -1130 -52 -701 23
rect -340 530 -277 531
rect -340 17 -338 530
rect -338 17 -279 530
rect -279 17 -277 530
rect -43 460 40 520
rect 222 464 305 524
rect -84 31 -83 368
rect -83 31 -37 368
rect -37 31 -32 368
rect 103 33 106 370
rect 106 33 155 370
rect 287 32 292 369
rect 292 32 339 369
rect 495 21 554 534
rect 554 21 558 534
rect 495 20 558 21
rect 738 123 785 460
rect 785 123 790 460
rect 922 122 971 459
rect 971 122 974 459
rect 1109 124 1114 461
rect 1114 124 1160 461
rect 1160 124 1161 461
rect 1305 122 1354 459
rect 1354 122 1357 459
rect 1492 124 1497 461
rect 1497 124 1543 461
rect 1543 124 1544 461
rect 1139 -29 1230 25
rect 1729 20 1788 533
rect 1788 20 1792 533
rect 1729 19 1792 20
rect 1977 123 2024 460
rect 2024 123 2029 460
rect 2161 122 2210 459
rect 2210 122 2213 459
rect 2348 124 2353 461
rect 2353 124 2399 461
rect 2399 124 2400 461
rect 2544 122 2593 459
rect 2593 122 2596 459
rect 2731 124 2736 461
rect 2736 124 2782 461
rect 2782 124 2783 461
rect 2218 -44 2341 26
rect 2981 31 3040 544
rect 3040 31 3044 544
rect 2981 30 3044 31
rect 3272 461 3353 517
rect 3534 465 3615 521
rect 3232 31 3233 368
rect 3233 31 3279 368
rect 3279 31 3284 368
rect 3419 33 3422 370
rect 3422 33 3471 370
rect 3603 32 3608 369
rect 3608 32 3655 369
rect 3830 34 3889 547
rect 3889 34 3893 547
rect 3830 33 3893 34
rect -1809 -222 -1404 -148
rect -740 -214 -335 -140
rect 104 -213 638 -143
rect 2834 -181 3374 -111
rect 3721 -185 4292 -119
rect 4813 -182 5384 -116
rect 1147 -251 1211 -249
rect 1147 -302 1211 -251
rect 2238 -250 2302 -248
rect 2238 -301 2302 -250
rect 310 -427 372 -341
rect -1715 -484 -1642 -431
rect -507 -607 -325 -553
rect 249 -618 373 -565
rect 899 -819 967 -394
rect 1075 -728 1121 -393
rect 1121 -728 1127 -393
rect 1234 -727 1237 -392
rect 1237 -727 1283 -392
rect 1283 -727 1286 -392
rect 1473 -811 1564 -378
rect 1932 -794 2023 -361
rect 2166 -727 2212 -393
rect 2212 -727 2218 -393
rect 2325 -726 2328 -391
rect 2328 -726 2374 -391
rect 2374 -726 2377 -391
rect 2497 -793 2573 -376
rect 3022 -396 3082 -303
rect 5154 -457 5249 -402
rect 2976 -584 3138 -527
rect 3908 -572 4309 -520
rect 1016 -893 1376 -888
rect -1627 -1003 -1089 -935
rect -739 -1007 -201 -939
rect 161 -995 638 -928
rect 1016 -980 1373 -893
rect 1373 -980 1376 -893
rect 2088 -892 2448 -888
rect 2088 -980 2099 -892
rect 2099 -980 2448 -892
rect 2910 -982 3280 -901
rect 3778 -973 4423 -903
rect 4747 -966 5392 -896
rect -68 -1708 38 -1192
rect 181 -1552 184 -1229
rect 184 -1552 233 -1229
rect 233 -1552 234 -1229
rect 346 -1552 349 -1229
rect 349 -1552 398 -1229
rect 398 -1552 399 -1229
rect 532 -1552 535 -1229
rect 535 -1552 584 -1229
rect 584 -1552 585 -1229
rect 697 -1552 700 -1229
rect 700 -1552 749 -1229
rect 749 -1552 750 -1229
rect 921 -1514 1028 -1044
rect 1241 -1089 1306 -1087
rect 1241 -1138 1242 -1089
rect 1242 -1138 1300 -1089
rect 1300 -1138 1306 -1089
rect 1241 -1139 1306 -1138
rect 1157 -1553 1160 -1230
rect 1160 -1553 1209 -1230
rect 1209 -1553 1210 -1230
rect 1322 -1552 1329 -1229
rect 1329 -1552 1375 -1229
rect 1706 -1531 1813 -1061
rect 2142 -1090 2201 -1086
rect 2142 -1139 2200 -1090
rect 2200 -1139 2201 -1090
rect 2057 -1554 2060 -1231
rect 2060 -1554 2109 -1231
rect 2109 -1554 2110 -1231
rect 2222 -1553 2229 -1226
rect 2229 -1553 2275 -1226
rect 2497 -1531 2604 -1061
rect 277 -1707 339 -1651
rect 589 -1705 655 -1649
rect 299 -2063 928 -1931
rect 1468 -2057 2097 -1925
rect 2933 -1953 2980 -1233
rect 2980 -1953 2985 -1233
rect 3095 -1958 3096 -1238
rect 3096 -1958 3144 -1238
rect 3144 -1958 3147 -1238
rect 3283 -1953 3330 -1233
rect 3330 -1953 3335 -1233
rect 3445 -1958 3446 -1238
rect 3446 -1958 3494 -1238
rect 3494 -1958 3497 -1238
rect 3702 -1904 3786 -1316
rect 3039 -2125 3101 -2068
rect 3310 -2124 3372 -2067
rect 2805 -2365 3466 -2271
<< metal2 >>
rect -2599 832 -2166 833
rect -2599 831 -2145 832
rect -2599 830 -602 831
rect -2717 816 -602 830
rect -2717 812 -1134 816
rect -2717 808 -1891 812
rect -2717 729 -2570 808
rect -2280 730 -1891 808
rect -1560 734 -1134 812
rect -803 734 -602 816
rect -1560 730 -602 734
rect -2280 729 -602 730
rect -2717 712 -602 729
rect -2716 -904 -2600 712
rect -2171 710 -602 712
rect -363 744 3922 770
rect -363 740 2082 744
rect -363 674 -212 740
rect 406 733 2082 740
rect 406 674 845 733
rect -363 667 845 674
rect 1463 676 2082 733
rect 2632 742 3922 744
rect 2632 676 3312 742
rect 1463 667 3312 676
rect -363 660 3312 667
rect 3827 660 3922 742
rect -363 639 3922 660
rect -363 531 -245 639
rect 204 543 320 544
rect 35 542 320 543
rect -2482 424 -1752 430
rect -2482 358 -2004 424
rect -1792 358 -1752 424
rect -2482 348 -1752 358
rect -1069 297 -977 300
rect -1069 239 -1054 297
rect -993 239 -977 297
rect -1069 236 -977 239
rect -363 50 -340 531
rect -2175 23 -340 50
rect -2175 -52 -1973 23
rect -1544 -52 -1130 23
rect -701 17 -340 23
rect -277 17 -245 531
rect -60 524 320 542
rect -60 520 222 524
rect -60 460 -43 520
rect 40 464 222 520
rect 305 464 320 524
rect 40 460 320 464
rect -60 445 320 460
rect 469 534 588 639
rect -60 443 238 445
rect -93 368 -24 379
rect -93 173 -84 368
rect -32 173 -24 368
rect -93 105 -85 173
rect -29 105 -24 173
rect -93 31 -84 105
rect -32 31 -24 105
rect 92 370 161 382
rect 92 78 103 370
rect -93 20 -24 31
rect 89 33 103 78
rect 155 78 161 370
rect 278 369 347 378
rect 278 344 287 369
rect 339 344 347 369
rect 278 277 282 344
rect 344 277 347 344
rect 155 33 162 78
rect -701 -42 -245 17
rect 89 -42 162 33
rect 278 32 287 277
rect 339 32 347 277
rect 278 19 347 32
rect 469 20 495 534
rect 558 20 588 534
rect 731 473 798 639
rect 730 460 799 473
rect 730 123 738 460
rect 790 123 799 460
rect 916 459 985 473
rect 916 362 922 459
rect 903 349 922 362
rect 974 349 985 459
rect 903 270 912 349
rect 979 270 985 349
rect 903 261 922 270
rect 730 114 799 123
rect 916 122 922 261
rect 974 122 985 270
rect 916 110 985 122
rect 1101 472 1168 639
rect 1101 461 1170 472
rect 1101 124 1109 461
rect 1161 124 1170 461
rect 1299 459 1368 473
rect 1485 472 1552 639
rect 1704 533 1822 639
rect 1969 582 2039 639
rect 2208 638 2832 639
rect 2340 586 2410 638
rect 2724 587 2794 638
rect 1299 360 1305 459
rect 1287 349 1305 360
rect 1357 349 1368 459
rect 1287 270 1297 349
rect 1364 270 1368 349
rect 1287 259 1305 270
rect 1101 113 1170 124
rect 1299 122 1305 259
rect 1357 122 1368 270
rect 1299 110 1368 122
rect 1484 461 1553 472
rect 1484 124 1492 461
rect 1544 124 1553 461
rect 1484 113 1553 124
rect 469 -42 588 20
rect 1114 25 1252 38
rect 1114 -29 1139 25
rect 1230 -29 1252 25
rect -701 -52 590 -42
rect 1114 -47 1252 -29
rect 1704 19 1729 533
rect 1792 19 1822 533
rect 1970 473 2037 582
rect 1969 460 2038 473
rect 1969 123 1977 460
rect 2029 123 2038 460
rect 1969 114 2038 123
rect 2155 459 2224 473
rect 2155 122 2161 459
rect 2213 348 2224 459
rect 2218 280 2224 348
rect 2213 122 2224 280
rect 2155 110 2224 122
rect 2340 472 2407 586
rect 2340 461 2409 472
rect 2340 124 2348 461
rect 2400 124 2409 461
rect 2340 113 2409 124
rect 2538 459 2607 473
rect 2724 472 2791 587
rect 2956 544 3074 639
rect 3599 637 3922 639
rect 2538 347 2544 459
rect 2596 347 2607 459
rect 2538 280 2542 347
rect 2598 280 2607 347
rect 2538 122 2544 280
rect 2596 122 2607 280
rect 2538 110 2607 122
rect 2723 461 2792 472
rect 2723 124 2731 461
rect 2783 124 2792 461
rect 2723 113 2792 124
rect -2175 -79 590 -52
rect -2169 -120 590 -79
rect 1116 -93 1244 -47
rect 1704 -73 1822 19
rect 2203 26 2360 37
rect 2203 -44 2218 26
rect 2341 -44 2360 26
rect 2203 -52 2360 -44
rect 2956 30 2981 544
rect 3044 30 3074 544
rect 3805 547 3922 637
rect 3257 540 3372 542
rect 3520 540 3635 541
rect 3257 521 3635 540
rect 3257 517 3534 521
rect 3257 461 3272 517
rect 3353 465 3534 517
rect 3615 465 3635 521
rect 3353 461 3635 465
rect 3257 443 3635 461
rect 3520 442 3635 443
rect 2956 -47 3074 30
rect 3223 368 3292 379
rect 3223 350 3232 368
rect 3284 350 3292 368
rect 3223 280 3230 350
rect 3286 280 3292 350
rect 3223 31 3232 280
rect 3284 31 3292 280
rect 3408 370 3477 382
rect 3408 48 3419 370
rect 3223 20 3292 31
rect 3406 33 3419 48
rect 3471 48 3477 370
rect 3594 369 3663 378
rect 3594 195 3603 369
rect 3655 195 3663 369
rect 3594 108 3600 195
rect 3656 108 3663 195
rect 3471 33 3486 48
rect 3406 -47 3486 33
rect 3594 32 3603 108
rect 3655 32 3663 108
rect 3594 19 3663 32
rect 3805 33 3830 547
rect 3893 33 3922 547
rect 3805 -47 3922 33
rect -2169 -137 728 -120
rect -2081 -140 728 -137
rect -2081 -148 -740 -140
rect -2081 -222 -1809 -148
rect -1404 -214 -740 -148
rect -335 -143 728 -140
rect -335 -213 104 -143
rect 638 -213 728 -143
rect -335 -214 728 -213
rect -1404 -222 728 -214
rect -2081 -239 728 -222
rect 1116 -176 1139 -93
rect 1220 -176 1244 -93
rect 1116 -239 1244 -176
rect -2081 -240 193 -239
rect 1117 -249 1244 -239
rect 2207 -102 2335 -52
rect 2953 -77 3926 -47
rect 2207 -180 2227 -102
rect 2307 -180 2335 -102
rect 2207 -240 2335 -180
rect 2761 -90 3926 -77
rect 5615 -90 5894 -89
rect 2761 -111 5894 -90
rect 2761 -181 2834 -111
rect 3374 -116 5894 -111
rect 3374 -119 4813 -116
rect 3374 -140 3721 -119
rect 3374 -181 3433 -140
rect 2761 -211 3433 -181
rect 3600 -185 3721 -140
rect 4292 -182 4813 -119
rect 5384 -182 5894 -116
rect 4292 -185 5894 -182
rect 3600 -208 5894 -185
rect 5615 -211 5894 -208
rect 1117 -302 1147 -249
rect 1211 -302 1244 -249
rect 1117 -317 1244 -302
rect 2208 -248 2335 -240
rect 2208 -301 2238 -248
rect 2302 -301 2335 -248
rect 2208 -316 2335 -301
rect 3003 -296 3093 -290
rect 3003 -303 3546 -296
rect 299 -318 390 -317
rect -96 -323 390 -318
rect -97 -341 390 -323
rect -2467 -424 -2279 -422
rect -2467 -431 -1627 -424
rect -2467 -484 -1715 -431
rect -1642 -484 -1627 -431
rect -2467 -489 -1627 -484
rect -97 -427 310 -341
rect 372 -427 390 -341
rect 1458 -326 1564 -324
rect -97 -443 390 -427
rect 882 -394 983 -343
rect 1458 -378 1582 -326
rect -2467 -490 -2279 -489
rect -97 -540 25 -443
rect -522 -553 25 -540
rect -522 -607 -507 -553
rect -325 -607 25 -553
rect -522 -614 25 -607
rect 183 -561 482 -546
rect 183 -618 249 -561
rect 373 -618 482 -561
rect 183 -624 482 -618
rect 882 -819 899 -394
rect 967 -819 983 -394
rect 1068 -393 1139 -381
rect 1068 -408 1075 -393
rect 1127 -408 1139 -393
rect 1068 -484 1072 -408
rect 1132 -484 1139 -408
rect 1068 -728 1075 -484
rect 1127 -728 1139 -484
rect 1068 -740 1139 -728
rect 1223 -392 1294 -381
rect 1223 -650 1234 -392
rect 1286 -650 1294 -392
rect 1223 -718 1231 -650
rect 1287 -718 1294 -650
rect 1223 -727 1234 -718
rect 1286 -727 1294 -718
rect 1223 -740 1294 -727
rect 882 -877 983 -819
rect 1458 -811 1473 -378
rect 1564 -811 1582 -378
rect 1458 -877 1582 -811
rect 1907 -361 2040 -329
rect 1907 -794 1932 -361
rect 2023 -794 2040 -361
rect 2158 -393 2229 -374
rect 2481 -376 2586 -328
rect 2158 -727 2166 -393
rect 2218 -515 2229 -393
rect 2314 -391 2385 -380
rect 2314 -409 2325 -391
rect 2377 -409 2385 -391
rect 2314 -482 2322 -409
rect 2379 -482 2385 -409
rect 2218 -650 2230 -515
rect 2226 -723 2230 -650
rect 2218 -727 2230 -723
rect 2158 -740 2230 -727
rect 2314 -726 2325 -482
rect 2377 -726 2385 -482
rect 2314 -739 2385 -726
rect 1907 -877 2040 -794
rect 2481 -793 2497 -376
rect 2573 -793 2586 -376
rect 3003 -396 3022 -303
rect 3082 -396 3546 -303
rect 3003 -410 3546 -396
rect 5141 -402 5880 -386
rect 2910 -527 3180 -509
rect 2910 -584 2976 -527
rect 3138 -584 3180 -527
rect 3458 -513 3545 -410
rect 5141 -457 5154 -402
rect 5249 -457 5880 -402
rect 5141 -469 5880 -457
rect 3848 -513 4358 -511
rect 3458 -520 4358 -513
rect 3458 -572 3908 -520
rect 4309 -572 4358 -520
rect 3458 -581 4358 -572
rect 3458 -583 3522 -581
rect 2910 -595 3180 -584
rect 2481 -874 2586 -793
rect 5612 -874 5891 -873
rect 2481 -877 5891 -874
rect 882 -888 5891 -877
rect 882 -901 1016 -888
rect -2716 -909 -2045 -904
rect 53 -909 1016 -901
rect -2716 -928 1016 -909
rect -2716 -935 161 -928
rect -2716 -1003 -1627 -935
rect -1089 -939 161 -935
rect -1089 -1003 -739 -939
rect -2716 -1007 -739 -1003
rect -201 -995 161 -939
rect 638 -980 1016 -928
rect 1376 -980 2088 -888
rect 2448 -896 5891 -888
rect 2448 -901 4747 -896
rect 2448 -980 2910 -901
rect 638 -982 2910 -980
rect 3280 -903 4747 -901
rect 3280 -973 3778 -903
rect 4423 -966 4747 -903
rect 5392 -966 5891 -896
rect 4423 -973 5891 -966
rect 3280 -982 5891 -973
rect 638 -994 5891 -982
rect 638 -995 3433 -994
rect -201 -998 3292 -995
rect -201 -1000 2624 -998
rect -201 -1007 1071 -1000
rect -2716 -1024 1071 -1007
rect -2716 -1029 233 -1024
rect -2716 -1033 -2045 -1029
rect -109 -1192 77 -1029
rect -109 -1708 -68 -1192
rect 38 -1708 77 -1192
rect 893 -1044 1043 -1024
rect 173 -1229 244 -1214
rect 173 -1552 181 -1229
rect 234 -1552 244 -1229
rect 173 -1569 244 -1552
rect 338 -1219 409 -1214
rect 524 -1219 595 -1214
rect 338 -1229 595 -1219
rect 338 -1552 346 -1229
rect 399 -1552 532 -1229
rect 585 -1552 595 -1229
rect 338 -1569 595 -1552
rect 689 -1229 760 -1214
rect 689 -1552 697 -1229
rect 750 -1552 760 -1229
rect 689 -1569 760 -1552
rect 893 -1514 921 -1044
rect 1028 -1514 1043 -1044
rect 1678 -1061 1828 -1000
rect 1214 -1083 1330 -1073
rect 1214 -1139 1241 -1083
rect 1306 -1139 1330 -1083
rect 1214 -1150 1330 -1139
rect -109 -1900 77 -1708
rect 178 -1640 241 -1569
rect 340 -1571 592 -1569
rect 420 -1628 509 -1571
rect 420 -1640 510 -1628
rect 690 -1640 759 -1569
rect 893 -1581 1043 -1514
rect 1149 -1230 1220 -1215
rect 1149 -1553 1157 -1230
rect 1210 -1553 1220 -1230
rect 1149 -1570 1220 -1553
rect 1312 -1229 1383 -1215
rect 1312 -1250 1322 -1229
rect 1312 -1327 1319 -1250
rect 1312 -1552 1322 -1327
rect 1375 -1552 1383 -1229
rect 1312 -1570 1383 -1552
rect 1678 -1531 1706 -1061
rect 1813 -1531 1828 -1061
rect 2469 -1061 2624 -1000
rect 2115 -1082 2230 -1073
rect 2115 -1139 2142 -1082
rect 2201 -1139 2230 -1082
rect 2115 -1153 2230 -1139
rect 178 -1649 759 -1640
rect 1151 -1649 1218 -1570
rect 1678 -1594 1828 -1531
rect 2049 -1231 2120 -1216
rect 2049 -1554 2057 -1231
rect 2110 -1254 2120 -1231
rect 2113 -1316 2120 -1254
rect 2110 -1554 2120 -1316
rect 2211 -1226 2281 -1214
rect 2211 -1349 2222 -1226
rect 2049 -1571 2120 -1554
rect 2212 -1553 2222 -1349
rect 2275 -1346 2281 -1226
rect 2275 -1553 2283 -1346
rect 2212 -1565 2283 -1553
rect 2210 -1571 2283 -1565
rect 2469 -1531 2497 -1061
rect 2604 -1531 2624 -1061
rect 3143 -1206 3292 -998
rect 178 -1651 589 -1649
rect 178 -1707 277 -1651
rect 339 -1705 589 -1651
rect 655 -1650 1218 -1649
rect 2210 -1650 2282 -1571
rect 2469 -1600 2624 -1531
rect 2927 -1233 2991 -1206
rect 2469 -1635 2623 -1600
rect 655 -1705 2283 -1650
rect 339 -1707 2283 -1705
rect 178 -1712 2283 -1707
rect 259 -1714 2283 -1712
rect 259 -1720 670 -1714
rect -109 -1901 102 -1900
rect 2468 -1901 2623 -1635
rect -109 -1925 2623 -1901
rect -109 -1931 1468 -1925
rect -109 -2063 299 -1931
rect 928 -2057 1468 -1931
rect 2097 -2057 2623 -1925
rect 2927 -1953 2933 -1233
rect 2985 -1772 2991 -1233
rect 2989 -1860 2991 -1772
rect 2985 -1953 2991 -1860
rect 2927 -1980 2991 -1953
rect 3088 -1233 3341 -1206
rect 3088 -1238 3283 -1233
rect 3088 -1958 3095 -1238
rect 3147 -1953 3283 -1238
rect 3335 -1953 3341 -1233
rect 3147 -1958 3341 -1953
rect 3088 -1964 3341 -1958
rect 3088 -1980 3152 -1964
rect 3277 -1980 3341 -1964
rect 3438 -1238 3502 -1206
rect 3438 -1767 3445 -1238
rect 3497 -1767 3502 -1238
rect 3438 -1849 3443 -1767
rect 3499 -1849 3502 -1767
rect 3438 -1958 3445 -1849
rect 3497 -1958 3502 -1849
rect 3438 -1980 3502 -1958
rect 3671 -1316 3824 -994
rect 5612 -995 5891 -994
rect 3671 -1904 3702 -1316
rect 3786 -1904 3824 -1316
rect 928 -2063 2623 -2057
rect -109 -2091 2623 -2063
rect -109 -2094 2348 -2091
rect 2468 -2236 2623 -2091
rect 3009 -2067 3416 -2050
rect 3009 -2068 3310 -2067
rect 3009 -2125 3039 -2068
rect 3101 -2124 3310 -2068
rect 3372 -2124 3416 -2067
rect 3101 -2125 3416 -2124
rect 3009 -2145 3416 -2125
rect 3671 -2236 3824 -1904
rect 2468 -2271 3825 -2236
rect 2468 -2365 2805 -2271
rect 3466 -2365 3825 -2271
rect 2468 -2391 3825 -2365
<< via2 >>
rect -1054 296 -993 297
rect -1054 243 -994 296
rect -994 243 -993 296
rect -1054 239 -993 243
rect -43 460 40 520
rect 222 464 305 524
rect -85 105 -84 173
rect -84 105 -32 173
rect -32 105 -29 173
rect 282 277 287 344
rect 287 277 339 344
rect 339 277 344 344
rect 912 270 922 349
rect 922 270 974 349
rect 974 270 979 349
rect 1297 270 1305 349
rect 1305 270 1357 349
rect 1357 270 1364 349
rect 2162 280 2213 348
rect 2213 280 2218 348
rect 2542 280 2544 347
rect 2544 280 2596 347
rect 2596 280 2598 347
rect 3272 461 3353 517
rect 3534 465 3615 521
rect 3230 280 3232 350
rect 3232 280 3284 350
rect 3284 280 3286 350
rect 3600 108 3603 195
rect 3603 108 3655 195
rect 3655 108 3656 195
rect 1139 -176 1220 -93
rect 2227 -180 2307 -102
rect 249 -565 373 -561
rect 249 -618 373 -565
rect 1072 -484 1075 -408
rect 1075 -484 1127 -408
rect 1127 -484 1132 -408
rect 1231 -718 1234 -650
rect 1234 -718 1286 -650
rect 1286 -718 1287 -650
rect 2322 -482 2325 -409
rect 2325 -482 2377 -409
rect 2377 -482 2379 -409
rect 2167 -723 2218 -650
rect 2218 -723 2226 -650
rect 2976 -584 3138 -527
rect 1241 -1087 1306 -1083
rect 1241 -1139 1306 -1087
rect 1319 -1327 1322 -1250
rect 1322 -1327 1375 -1250
rect 2142 -1086 2201 -1082
rect 2142 -1139 2201 -1086
rect 2057 -1316 2110 -1254
rect 2110 -1316 2113 -1254
rect 277 -1707 339 -1651
rect 589 -1705 655 -1649
rect 2933 -1860 2985 -1772
rect 2985 -1860 2989 -1772
rect 3443 -1849 3445 -1767
rect 3445 -1849 3497 -1767
rect 3497 -1849 3499 -1767
rect 3039 -2125 3101 -2068
rect 3310 -2124 3372 -2067
<< metal3 >>
rect 204 543 320 544
rect 35 542 3372 543
rect -60 540 3372 542
rect 3520 540 3635 541
rect -404 539 3635 540
rect -511 524 3635 539
rect -511 520 222 524
rect -511 460 -43 520
rect 40 464 222 520
rect 305 517 3407 524
rect 305 464 3272 517
rect 40 461 3272 464
rect 3353 461 3407 517
rect 40 460 3407 461
rect 3480 521 3635 524
rect 3480 465 3534 521
rect 3615 465 3635 521
rect 3480 460 3635 465
rect -511 446 3635 460
rect -511 303 -420 446
rect -60 445 320 446
rect -60 443 238 445
rect 3257 443 3635 446
rect 3520 442 3635 443
rect 278 358 1374 359
rect 278 354 1918 358
rect -1070 297 -420 303
rect -1070 239 -1054 297
rect -993 239 -420 297
rect 277 349 1918 354
rect 277 344 912 349
rect 277 277 282 344
rect 344 277 912 344
rect 277 270 912 277
rect 979 270 1297 349
rect 1364 270 1918 349
rect 2134 350 3298 362
rect 2134 348 3230 350
rect 2134 280 2162 348
rect 2218 347 3230 348
rect 2218 280 2542 347
rect 2598 280 3230 347
rect 3286 280 3298 350
rect 2134 270 3298 280
rect 277 268 1918 270
rect 278 267 1918 268
rect 907 262 1918 267
rect -1070 235 -420 239
rect 728 187 826 189
rect -87 173 826 187
rect -87 105 -85 173
rect -29 105 826 173
rect -87 92 826 105
rect 183 -561 482 -546
rect 183 -618 249 -561
rect 373 -618 482 -561
rect 183 -624 482 -618
rect 728 -638 826 92
rect 911 -393 991 262
rect 1311 259 1918 262
rect 1234 -77 1492 -71
rect 1115 -93 1517 -77
rect 1115 -176 1139 -93
rect 1220 -176 1517 -93
rect 1115 -187 1517 -176
rect 1234 -191 1517 -187
rect 911 -408 1140 -393
rect 911 -422 1072 -408
rect 911 -483 980 -422
rect 1044 -483 1072 -422
rect 911 -484 1072 -483
rect 1132 -484 1140 -408
rect 911 -499 1140 -484
rect 1433 -398 1517 -191
rect 1822 -90 1918 259
rect 1822 -91 2285 -90
rect 1822 -102 2330 -91
rect 1822 -180 2227 -102
rect 2307 -180 2330 -102
rect 1822 -201 2330 -180
rect 1822 -202 2285 -201
rect 2562 -398 2646 270
rect 3222 269 3298 270
rect 2720 195 3659 205
rect 2720 108 3600 195
rect 3656 108 3659 195
rect 2720 95 3659 108
rect 1433 -409 2648 -398
rect 1433 -482 2322 -409
rect 2379 -415 2648 -409
rect 2379 -482 2402 -415
rect 1433 -483 2402 -482
rect 2460 -483 2648 -415
rect 1433 -489 2648 -483
rect 1433 -493 2499 -489
rect 911 -500 1056 -499
rect 728 -650 1589 -638
rect 2720 -639 2831 95
rect 2910 -527 3180 -509
rect 2910 -584 2976 -527
rect 3138 -584 3180 -527
rect 2910 -595 3180 -584
rect 1989 -640 2832 -639
rect 728 -718 1231 -650
rect 1287 -718 1589 -650
rect 728 -729 1589 -718
rect 728 -732 826 -729
rect 1266 -732 1589 -729
rect 1912 -650 2832 -640
rect 1912 -723 2167 -650
rect 2226 -723 2832 -650
rect 1912 -730 2832 -723
rect 1912 -732 2253 -730
rect 1214 -1074 1330 -1073
rect -363 -1075 1331 -1074
rect -605 -1083 1331 -1075
rect -605 -1139 1241 -1083
rect 1306 -1139 1331 -1083
rect -605 -1157 1331 -1139
rect -605 -1158 1089 -1157
rect 1497 -1237 1588 -732
rect 1315 -1238 1588 -1237
rect 1313 -1250 1588 -1238
rect 1313 -1327 1319 -1250
rect 1375 -1327 1588 -1250
rect 1912 -1244 1998 -732
rect 2115 -1082 4464 -1070
rect 2115 -1139 2142 -1082
rect 2201 -1139 4464 -1082
rect 2115 -1153 4464 -1139
rect 1912 -1254 2120 -1244
rect 1912 -1316 2057 -1254
rect 2113 -1316 2120 -1254
rect 1912 -1325 2120 -1316
rect 2049 -1327 2120 -1325
rect 1313 -1340 1588 -1327
rect 1315 -1341 1581 -1340
rect 259 -1649 670 -1640
rect 259 -1651 589 -1649
rect 259 -1707 277 -1651
rect 339 -1705 589 -1651
rect 655 -1705 670 -1649
rect 339 -1707 670 -1705
rect 259 -1720 670 -1707
rect 399 -1756 670 -1720
rect 399 -1758 1780 -1756
rect 399 -1760 1861 -1758
rect 399 -1762 2312 -1760
rect 399 -1767 3515 -1762
rect 399 -1772 3443 -1767
rect 399 -1860 2933 -1772
rect 2989 -1849 3443 -1772
rect 3499 -1849 3515 -1767
rect 2989 -1860 3515 -1849
rect 399 -1863 3515 -1860
rect 480 -1865 3515 -1863
rect 931 -1867 3515 -1865
rect 2149 -1868 3515 -1867
rect 2149 -1874 2887 -1868
rect 3009 -2063 3416 -2050
rect 3009 -2068 3171 -2063
rect 3009 -2125 3039 -2068
rect 3101 -2120 3171 -2068
rect 3239 -2067 3416 -2063
rect 3239 -2120 3310 -2067
rect 3101 -2124 3310 -2120
rect 3372 -2124 3416 -2067
rect 3101 -2125 3416 -2124
rect 3009 -2145 3416 -2125
<< via3 >>
rect 3407 460 3480 524
rect 249 -618 373 -561
rect 980 -483 1044 -422
rect 2402 -483 2460 -415
rect 2976 -584 3138 -527
rect 3171 -2120 3239 -2063
<< metal4 >>
rect 3368 524 3513 548
rect 3368 460 3407 524
rect 3480 460 3513 524
rect 3368 441 3513 460
rect 969 -422 1059 -396
rect 969 -483 980 -422
rect 1044 -483 1059 -422
rect 969 -545 1059 -483
rect 2394 -415 2472 -398
rect 2394 -483 2402 -415
rect 2460 -483 2472 -415
rect 2394 -507 2472 -483
rect 2394 -527 3188 -507
rect 183 -561 1060 -545
rect 183 -618 249 -561
rect 373 -618 1060 -561
rect 2394 -584 2976 -527
rect 3138 -584 3188 -527
rect 2394 -593 3188 -584
rect 2394 -595 3180 -593
rect 183 -624 1060 -618
rect 3368 -2044 3512 441
rect 3360 -2046 3512 -2044
rect 3130 -2063 3512 -2046
rect 3130 -2120 3171 -2063
rect 3239 -2120 3512 -2063
rect 3130 -2146 3512 -2120
use gf180mcu_fd_sc_mcu7t5v0__buf_4  gf180mcu_fd_sc_mcu7t5v0__buf_4_0 ~/conda-gf180mcu-env/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform 1 0 -2172 0 -1 772
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  gf180mcu_fd_sc_mcu7t5v0__inv_2_0 ~/conda-gf180mcu-env/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1757859342
transform 1 0 53 0 1 -965
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  gf180mcu_fd_sc_mcu7t5v0__inv_2_1
timestamp 1757859342
transform 1 0 2760 0 1 -934
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  gf180mcu_fd_sc_mcu7t5v0__inv_8_0 ~/conda-gf180mcu-env/envs/gf180mcu-env/share/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1753044640
transform -1 0 -68 0 1 -965
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  gf180mcu_fd_sc_mcu7t5v0__inv_8_1
timestamp 1753044640
transform 1 0 3601 0 1 -934
box -86 -86 2102 870
<< labels >>
flabel metal3 594 267 694 354 0 FreeSans 320 0 0 0 OUT_NI
flabel metal3 2809 285 2927 346 0 FreeSans 320 0 0 0 OUT_PI
flabel metal3 -570 244 -447 290 0 FreeSans 320 0 0 0 ENi
flabel metal2 -2480 348 -2386 430 0 FreeSans 320 0 0 0 EN
port 5 nsew
flabel metal2 -2466 -490 -2368 -423 0 FreeSans 320 0 0 0 OUT_N
port 6 nsew
flabel metal2 5771 -466 5873 -393 0 FreeSans 320 0 0 0 OUT_P
port 7 nsew
flabel metal3 -603 -1158 -494 -1076 0 FreeSans 320 0 0 0 VIN_P
port 1 nsew
flabel metal3 4351 -1152 4460 -1070 0 FreeSans 320 0 0 0 VIN_N
port 2 nsew
flabel metal2 5615 -211 5894 -89 0 FreeSans 320 0 0 0 VDD
port 3 nsew
flabel metal2 5620 -995 5889 -874 0 FreeSans 320 0 0 0 VSS
port 4 nsew
<< end >>
