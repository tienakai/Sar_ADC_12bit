magic
tech gf180mcuD
magscale 1 10
timestamp 1757235861
<< nwell >>
rect 27 7430 1587 7722
rect 27 7370 1588 7430
rect 28 5491 1588 7370
rect 29 5379 1588 5491
<< pwell >>
rect 1589 7718 3183 7722
rect 1589 7364 3480 7718
rect 1589 7359 3455 7364
rect 1589 5592 3476 7359
rect 1589 5380 3477 5592
<< nmos >>
rect 1764 5692 1820 7292
rect 1924 5692 1980 7292
rect 2084 5692 2140 7292
rect 2244 5692 2300 7292
rect 2532 5692 2588 7292
rect 2692 5692 2748 7292
rect 2852 5692 2908 7292
rect 3012 5692 3068 7292
rect 3308 5691 3364 7291
<< pmos >>
rect 202 5690 258 7290
rect 362 5690 418 7290
rect 522 5690 578 7290
rect 682 5690 738 7290
rect 842 5690 898 7290
rect 1002 5690 1058 7290
rect 1162 5690 1218 7290
rect 1322 5690 1378 7290
<< ndiff >>
rect 1676 7279 1764 7292
rect 1676 5705 1689 7279
rect 1735 5705 1764 7279
rect 1676 5692 1764 5705
rect 1820 7279 1924 7292
rect 1820 5705 1849 7279
rect 1895 5705 1924 7279
rect 1820 5692 1924 5705
rect 1980 7279 2084 7292
rect 1980 5705 2009 7279
rect 2055 5705 2084 7279
rect 1980 5692 2084 5705
rect 2140 7279 2244 7292
rect 2140 5705 2169 7279
rect 2215 5705 2244 7279
rect 2140 5692 2244 5705
rect 2300 7279 2388 7292
rect 2300 5705 2329 7279
rect 2375 5705 2388 7279
rect 2300 5692 2388 5705
rect 2444 7279 2532 7292
rect 2444 5705 2457 7279
rect 2503 5705 2532 7279
rect 2444 5692 2532 5705
rect 2588 7279 2692 7292
rect 2588 5705 2617 7279
rect 2663 5705 2692 7279
rect 2588 5692 2692 5705
rect 2748 7279 2852 7292
rect 2748 5705 2777 7279
rect 2823 5705 2852 7279
rect 2748 5692 2852 5705
rect 2908 7279 3012 7292
rect 2908 5705 2937 7279
rect 2983 5705 3012 7279
rect 2908 5692 3012 5705
rect 3068 7279 3156 7292
rect 3068 5705 3097 7279
rect 3143 5705 3156 7279
rect 3068 5692 3156 5705
rect 3220 7278 3308 7291
rect 3220 5704 3233 7278
rect 3279 5704 3308 7278
rect 3220 5691 3308 5704
rect 3364 7278 3452 7291
rect 3364 5704 3393 7278
rect 3439 5704 3452 7278
rect 3364 5691 3452 5704
<< pdiff >>
rect 114 7277 202 7290
rect 114 5703 127 7277
rect 173 5703 202 7277
rect 114 5690 202 5703
rect 258 7277 362 7290
rect 258 5703 287 7277
rect 333 5703 362 7277
rect 258 5690 362 5703
rect 418 7277 522 7290
rect 418 5703 447 7277
rect 493 5703 522 7277
rect 418 5690 522 5703
rect 578 7277 682 7290
rect 578 5703 607 7277
rect 653 5703 682 7277
rect 578 5690 682 5703
rect 738 7277 842 7290
rect 738 5703 767 7277
rect 813 5703 842 7277
rect 738 5690 842 5703
rect 898 7277 1002 7290
rect 898 5703 927 7277
rect 973 5703 1002 7277
rect 898 5690 1002 5703
rect 1058 7277 1162 7290
rect 1058 5703 1087 7277
rect 1133 5703 1162 7277
rect 1058 5690 1162 5703
rect 1218 7277 1322 7290
rect 1218 5703 1247 7277
rect 1293 5703 1322 7277
rect 1218 5690 1322 5703
rect 1378 7277 1466 7290
rect 1378 5703 1407 7277
rect 1453 5703 1466 7277
rect 1378 5690 1466 5703
<< ndiffc >>
rect 1689 5705 1735 7279
rect 1849 5705 1895 7279
rect 2009 5705 2055 7279
rect 2169 5705 2215 7279
rect 2329 5705 2375 7279
rect 2457 5705 2503 7279
rect 2617 5705 2663 7279
rect 2777 5705 2823 7279
rect 2937 5705 2983 7279
rect 3097 5705 3143 7279
rect 3233 5704 3279 7278
rect 3393 5704 3439 7278
<< pdiffc >>
rect 127 5703 173 7277
rect 287 5703 333 7277
rect 447 5703 493 7277
rect 607 5703 653 7277
rect 767 5703 813 7277
rect 927 5703 973 7277
rect 1087 5703 1133 7277
rect 1247 5703 1293 7277
rect 1407 5703 1453 7277
<< psubdiff >>
rect 1677 5524 3469 5579
rect 1677 5523 2774 5524
rect 1677 5452 1759 5523
rect 2296 5453 2774 5523
rect 3311 5453 3469 5524
rect 2296 5452 3469 5453
rect 1677 5411 3469 5452
<< nsubdiff >>
rect 108 7641 1548 7678
rect 108 7528 148 7641
rect 734 7640 1548 7641
rect 734 7528 923 7640
rect 108 7527 923 7528
rect 1509 7527 1548 7640
rect 108 7510 1548 7527
<< psubdiffcont >>
rect 1759 5452 2296 5523
rect 2774 5453 3311 5524
<< nsubdiffcont >>
rect 148 7528 734 7641
rect 923 7527 1509 7640
<< polysilicon >>
rect 202 7334 1378 7390
rect 202 7290 258 7334
rect 362 7290 418 7334
rect 522 7290 578 7334
rect 682 7290 738 7334
rect 842 7290 898 7334
rect 1002 7290 1058 7334
rect 1162 7290 1218 7334
rect 1322 7290 1378 7334
rect 1764 7331 2301 7392
rect 1764 7292 1820 7331
rect 1924 7292 1980 7331
rect 2084 7292 2140 7331
rect 2244 7292 2300 7331
rect 2532 7330 3069 7391
rect 3263 7330 3401 7391
rect 2532 7292 2588 7330
rect 2692 7292 2748 7330
rect 2852 7292 2908 7330
rect 3012 7292 3068 7330
rect 3308 7291 3364 7330
rect 202 5646 258 5690
rect 362 5646 418 5690
rect 522 5646 578 5690
rect 682 5646 738 5690
rect 842 5646 898 5690
rect 1002 5646 1058 5690
rect 1162 5646 1218 5690
rect 1322 5646 1378 5690
rect 1764 5648 1820 5692
rect 1924 5648 1980 5692
rect 2084 5648 2140 5692
rect 2244 5648 2300 5692
rect 2532 5648 2588 5692
rect 2692 5648 2748 5692
rect 2852 5648 2908 5692
rect 3012 5648 3068 5692
rect 3308 5647 3364 5691
<< metal1 >>
rect 108 7641 1548 7678
rect 108 7528 148 7641
rect 734 7640 1548 7641
rect 734 7528 923 7640
rect 108 7527 923 7528
rect 1509 7527 1548 7640
rect 108 7510 1548 7527
rect 127 7277 173 7288
rect 287 7277 333 7288
rect 173 7240 183 7255
rect 181 7179 183 7240
rect 173 7165 183 7179
rect 127 5692 173 5703
rect 447 7277 493 7288
rect 607 7277 653 7288
rect 493 7241 505 7255
rect 502 7180 505 7241
rect 333 5801 343 5817
rect 339 5731 343 5801
rect 333 5719 343 5731
rect 287 5692 333 5703
rect 493 7165 505 7180
rect 447 5692 493 5703
rect 767 7277 813 7288
rect 927 7277 973 7288
rect 813 7241 826 7255
rect 822 7180 826 7241
rect 653 5800 663 5815
rect 659 5730 663 5800
rect 653 5717 663 5730
rect 607 5692 653 5703
rect 813 7165 826 7180
rect 767 5692 813 5703
rect 1087 7277 1133 7288
rect 1247 7277 1293 7288
rect 1133 7240 1146 7255
rect 1142 7179 1146 7240
rect 973 5801 983 5815
rect 980 5731 983 5801
rect 973 5717 983 5731
rect 927 5692 973 5703
rect 1133 7165 1146 7179
rect 1087 5692 1133 5703
rect 1407 7277 1453 7288
rect 1689 7279 1735 7290
rect 1453 7241 1467 7256
rect 1461 7180 1467 7241
rect 1293 5800 1302 5815
rect 1300 5730 1302 5800
rect 1293 5717 1302 5730
rect 1247 5692 1293 5703
rect 1453 7166 1467 7180
rect 1687 6997 1689 7102
rect 1849 7279 1895 7290
rect 1735 7087 1746 7102
rect 1744 7011 1746 7087
rect 1407 5692 1453 5703
rect 1735 6997 1746 7011
rect 1689 5694 1735 5705
rect 2009 7279 2055 7290
rect 2169 7279 2215 7290
rect 2055 7086 2069 7102
rect 2065 7010 2069 7086
rect 1895 5801 1905 5815
rect 1901 5731 1905 5801
rect 1895 5717 1905 5731
rect 1849 5694 1895 5705
rect 2055 6997 2069 7010
rect 2168 5715 2169 5813
rect 2329 7279 2375 7290
rect 2328 6994 2329 7099
rect 2457 7279 2503 7290
rect 2375 7086 2387 7099
rect 2386 7010 2387 7086
rect 2215 5800 2223 5813
rect 2222 5730 2223 5800
rect 2009 5694 2055 5705
rect 2215 5715 2223 5730
rect 2169 5694 2215 5705
rect 2375 6994 2387 7010
rect 2329 5694 2375 5705
rect 2617 7279 2663 7290
rect 2503 6918 2514 6931
rect 2513 6841 2514 6918
rect 2503 6829 2514 6841
rect 2616 5717 2617 5815
rect 2777 7279 2823 7290
rect 2937 7279 2983 7290
rect 2823 6917 2835 6929
rect 2834 6840 2835 6917
rect 2663 5800 2671 5815
rect 2669 5730 2671 5800
rect 2457 5694 2503 5705
rect 2663 5717 2671 5730
rect 2617 5694 2663 5705
rect 2823 6827 2835 6840
rect 2777 5694 2823 5705
rect 3097 7279 3143 7290
rect 3233 7278 3279 7289
rect 3143 6918 3155 6931
rect 3154 6841 3155 6918
rect 2983 5801 2990 5813
rect 2983 5716 2990 5731
rect 2937 5694 2983 5705
rect 3143 6829 3155 6841
rect 3097 5694 3143 5705
rect 3393 7278 3439 7289
rect 3279 6741 3290 6755
rect 3289 6670 3290 6741
rect 3279 6657 3290 6670
rect 3233 5693 3279 5704
rect 3439 5801 3446 5813
rect 3439 5716 3446 5731
rect 3393 5693 3439 5704
rect 1677 5524 3469 5579
rect 1677 5523 2774 5524
rect 1677 5452 1759 5523
rect 2296 5453 2774 5523
rect 3311 5453 3469 5524
rect 2296 5452 3469 5453
rect 1677 5411 3469 5452
<< via1 >>
rect 127 7179 173 7240
rect 173 7179 181 7240
rect 448 7180 493 7241
rect 493 7180 502 7241
rect 287 5731 333 5801
rect 333 5731 339 5801
rect 768 7180 813 7241
rect 813 7180 822 7241
rect 607 5730 653 5800
rect 653 5730 659 5800
rect 1088 7179 1133 7240
rect 1133 7179 1142 7240
rect 928 5731 973 5801
rect 973 5731 980 5801
rect 1407 7180 1453 7241
rect 1453 7180 1461 7241
rect 1248 5730 1293 5800
rect 1293 5730 1300 5800
rect 1689 7011 1735 7087
rect 1735 7011 1744 7087
rect 2010 7010 2055 7086
rect 2055 7010 2065 7086
rect 1849 5731 1895 5801
rect 1895 5731 1901 5801
rect 2331 7010 2375 7086
rect 2375 7010 2386 7086
rect 2170 5730 2215 5800
rect 2215 5730 2222 5800
rect 2458 6841 2503 6918
rect 2503 6841 2513 6918
rect 2779 6840 2823 6917
rect 2823 6840 2834 6917
rect 2617 5730 2663 5800
rect 2663 5730 2669 5800
rect 3099 6841 3143 6918
rect 3143 6841 3154 6918
rect 2938 5731 2983 5801
rect 2983 5731 2990 5801
rect 3234 6670 3279 6741
rect 3279 6670 3289 6741
rect 3394 5731 3439 5801
rect 3439 5731 3446 5801
<< metal2 >>
rect 116 7241 1474 7258
rect 116 7240 448 7241
rect 116 7179 127 7240
rect 181 7180 448 7240
rect 502 7180 768 7241
rect 822 7240 1407 7241
rect 822 7180 1088 7240
rect 181 7179 1088 7180
rect 1142 7180 1407 7240
rect 1461 7180 1474 7241
rect 1142 7179 1474 7180
rect 116 7171 1474 7179
rect 1679 7087 2403 7100
rect 1679 7011 1689 7087
rect 1744 7086 2403 7087
rect 1744 7011 2010 7086
rect 1679 7010 2010 7011
rect 2065 7010 2331 7086
rect 2386 7010 2403 7086
rect 1679 7003 2403 7010
rect 2445 6918 3163 6931
rect 2445 6841 2458 6918
rect 2513 6917 3099 6918
rect 2513 6841 2779 6917
rect 2445 6840 2779 6841
rect 2834 6841 3099 6917
rect 3154 6841 3163 6918
rect 2834 6840 3163 6841
rect 2445 6828 3163 6840
rect 3231 6741 3293 6754
rect 3231 6670 3234 6741
rect 3289 6670 3293 6741
rect 3231 6657 3293 6670
rect 3392 5810 3448 5814
rect 279 5801 3451 5810
rect 279 5731 287 5801
rect 339 5800 928 5801
rect 339 5731 607 5800
rect 279 5730 607 5731
rect 659 5731 928 5800
rect 980 5800 1849 5801
rect 980 5731 1248 5800
rect 659 5730 1248 5731
rect 1300 5731 1849 5800
rect 1901 5800 2938 5801
rect 1901 5731 2170 5800
rect 1300 5730 2170 5731
rect 2222 5730 2617 5800
rect 2669 5731 2938 5800
rect 2990 5731 3394 5801
rect 3446 5731 3451 5801
rect 2669 5730 3451 5731
rect 279 5722 3451 5730
rect 3392 5716 3448 5722
<< labels >>
flabel metal2 1773 7008 2295 7086 0 FreeSans 320 0 0 0 VCM
port 1 nsew
flabel metal2 2572 6842 3094 6920 0 FreeSans 320 0 0 0 VREF_GND
port 2 nsew
flabel metal2 3235 6661 3290 6750 0 FreeSans 320 0 0 0 VIN
port 3 nsew
flabel metal2 384 7179 1187 7243 0 FreeSans 320 0 0 0 VREF
port 4 nsew
flabel polysilicon 1800 7338 2288 7383 0 FreeSans 320 0 0 0 EN_VCM
port 5 nsew
flabel polysilicon 292 7341 1290 7380 0 FreeSans 320 0 0 0 EN_VREF_Z
port 6 nsew
flabel metal2 1019 5734 2434 5788 0 FreeSans 320 0 0 0 Cbtm
port 7 nsew
flabel metal1 337 7541 1454 7654 0 FreeSans 320 0 0 0 VDD
port 8 nsew
flabel polysilicon 2609 7334 3020 7377 0 FreeSans 320 0 0 0 EN_VSS
port 9 nsew
flabel polysilicon 3270 7336 3398 7386 0 FreeSans 320 0 0 0 EN_VIN
port 10 nsew
flabel metal1 1840 5436 3254 5543 0 FreeSans 320 0 0 0 VSS
port 11 nsew
<< end >>
