magic
tech gf180mcuD
magscale 1 10
timestamp 1757729720
<< pwell >>
rect -220 -268 220 268
<< nmos >>
rect -108 -200 -52 200
rect 52 -200 108 200
<< ndiff >>
rect -196 187 -108 200
rect -196 -187 -183 187
rect -137 -187 -108 187
rect -196 -200 -108 -187
rect -52 187 52 200
rect -52 -187 -23 187
rect 23 -187 52 187
rect -52 -200 52 -187
rect 108 187 196 200
rect 108 -187 137 187
rect 183 -187 196 187
rect 108 -200 196 -187
<< ndiffc >>
rect -183 -187 -137 187
rect -23 -187 23 187
rect 137 -187 183 187
<< polysilicon >>
rect -108 200 -52 244
rect 52 200 108 244
rect -108 -244 -52 -200
rect 52 -244 108 -200
<< metal1 >>
rect -183 187 -137 198
rect -183 -198 -137 -187
rect -23 187 23 198
rect -23 -198 23 -187
rect 137 187 183 198
rect 137 -198 183 -187
<< properties >>
string gencell nfet_03v3
string library gf180mcu
string parameters w 2 l 0.280 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 0 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt}
<< end >>
